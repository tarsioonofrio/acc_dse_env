library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package inmem_package is
  type mem is array(0 to 4000000) of integer;

  constant input_mem : mem := (
    -- bias
    4603, 4862, -1029, -1549, -1741, 104, 1133, -2119, -2893, -2933, -4656, 3088, -1008, 350, -916, -2930, 6183, -2148, -4094, 3410, 7695, 12126, 3075, -3592, -2059, -4520, 7420, -4440, 1656, 550, -2306, 9666, -9757, -3830, -6395, 688, 6821, 11147, -2186, 2130, 10877, -3468, 944, 459, 6164, 5549, 2778, 7982, 1669, -2435, 2656, 2752, -1842, -2322, -2315, -1632, -2046, 48, 1973, 432, 253, 1502, 1413, -1822, 3539, 1569, -4710, 4002, 5073, -1002, 4573, 7031, 3062, -3286, -2061, -1082, 8944, 1909, -738, -4543, -636, -1032, 74, 198, -5642, -1173, -4970, -2191, 9720, -2956, 11478, 678, 1359, 1440, -1223, -829, -494, 2675, -13158, -1782, -3650, 67, -2439, 5762, 3579, 6231, 4887, 7078, -2464, -12046, -1602, 1518, 1069, 640, -5579, -1301, -7060, 3981, 2789, -3005, -5571, -1621, 18799, 119, 971, -943, -5689, 258,

    -- weights
    -- filter=0 channel=0
    -10, -10, 1, 7, 5, -5, -5, -5, -16,
    -- filter=0 channel=1
    28, 38, 10, 36, 51, 29, 19, 27, 32,
    -- filter=0 channel=2
    19, 29, 36, 32, 46, 41, 20, 28, 26,
    -- filter=0 channel=3
    16, 17, 7, 13, 21, -2, -4, 12, -2,
    -- filter=0 channel=4
    -8, -11, -3, -13, -10, -18, -20, -16, -15,
    -- filter=0 channel=5
    -10, -10, -2, -5, -5, -8, 4, -2, 2,
    -- filter=0 channel=6
    7, 9, 11, -3, 12, -1, 7, 1, 3,
    -- filter=0 channel=7
    2, -2, 6, 2, -3, 0, -4, -2, 9,
    -- filter=0 channel=8
    -20, -14, -15, -24, -14, -24, -15, -19, -21,
    -- filter=0 channel=9
    -15, -5, 15, -1, 0, 5, 3, 1, 9,
    -- filter=0 channel=10
    9, 18, 7, 16, 11, 13, 3, 14, 4,
    -- filter=0 channel=11
    6, 12, 7, 7, 1, 8, -2, 0, 6,
    -- filter=0 channel=12
    -2, -10, -6, -8, -4, -4, -7, 1, 4,
    -- filter=0 channel=13
    -6, -15, -7, -9, -22, -4, 0, -16, -1,
    -- filter=0 channel=14
    -9, 6, -4, -14, -5, 7, 6, -10, 6,
    -- filter=0 channel=15
    -18, 0, -15, -14, -6, -11, -5, -22, -17,
    -- filter=0 channel=16
    5, 1, 12, -2, 13, 15, 3, -6, -6,
    -- filter=0 channel=17
    0, -18, -8, -10, -2, -16, -15, -8, -15,
    -- filter=0 channel=18
    -4, -27, -2, -17, -36, -26, -22, -34, -14,
    -- filter=0 channel=19
    17, 15, 6, 15, 22, 10, 19, 26, 18,
    -- filter=0 channel=20
    3, 5, 0, -1, -5, 2, -4, -7, 2,
    -- filter=0 channel=21
    9, -2, 12, -3, -3, -8, -6, 1, 3,
    -- filter=0 channel=22
    -9, -10, 8, 6, 5, -10, -7, -10, -1,
    -- filter=0 channel=23
    24, 17, 3, 23, 23, 0, 2, 21, 8,
    -- filter=0 channel=24
    -15, -21, -15, -18, -12, 3, -14, -13, 0,
    -- filter=0 channel=25
    40, 56, 34, 45, 63, 30, 46, 60, 33,
    -- filter=0 channel=26
    6, 14, -2, 3, 23, 12, 17, 23, -2,
    -- filter=0 channel=27
    9, 32, 16, 15, 23, 12, 25, 29, 19,
    -- filter=0 channel=28
    -11, -6, -7, -23, -11, 5, -8, -15, -12,
    -- filter=0 channel=29
    -3, 4, 8, -20, -15, -11, -19, -7, -15,
    -- filter=0 channel=30
    12, 10, 4, 18, 17, 18, 19, 9, 12,
    -- filter=0 channel=31
    10, 0, 3, 11, 5, -7, 1, 1, 0,
    -- filter=0 channel=32
    20, 29, 24, 31, 35, 38, 19, 25, 18,
    -- filter=0 channel=33
    7, 0, 7, -5, -8, 3, 6, -1, 0,
    -- filter=0 channel=34
    -9, 5, 7, -1, -10, 0, 4, -3, 6,
    -- filter=0 channel=35
    39, 53, 12, 39, 46, 32, 27, 33, 22,
    -- filter=0 channel=36
    0, 1, 10, -5, 14, -4, 12, 5, 12,
    -- filter=0 channel=37
    -9, -4, 0, -2, 2, 4, 3, 12, 12,
    -- filter=0 channel=38
    12, 6, 4, 11, 30, 3, -3, 10, 7,
    -- filter=0 channel=39
    10, 0, 4, -1, 4, -6, -9, 9, 6,
    -- filter=0 channel=40
    8, 14, 13, 2, 0, 3, 14, 12, 12,
    -- filter=0 channel=41
    8, 6, -6, -16, 7, -3, 0, 8, -1,
    -- filter=0 channel=42
    -2, -1, 4, -4, -10, -3, 3, -2, -6,
    -- filter=0 channel=43
    1, 25, 17, 17, 22, 24, 12, 26, 15,
    -- filter=0 channel=44
    16, 16, 14, 20, 25, 16, 28, 21, 23,
    -- filter=0 channel=45
    0, 0, -10, -9, -8, -8, 9, -4, -3,
    -- filter=0 channel=46
    -6, -8, 3, 1, 8, 6, -2, 1, -5,
    -- filter=0 channel=47
    -1, 8, -2, -5, 0, -8, 10, 9, 6,
    -- filter=0 channel=48
    -1, -7, -6, 0, -9, 7, 9, -4, -4,
    -- filter=0 channel=49
    7, 16, 9, 3, -4, -6, 5, -7, 5,
    -- filter=0 channel=50
    9, 11, 3, 3, 19, 7, 11, 5, 0,
    -- filter=0 channel=51
    -11, -4, 0, -4, -10, -12, 1, -9, -11,
    -- filter=0 channel=52
    11, -1, 8, 7, -2, 9, 11, 8, 4,
    -- filter=0 channel=53
    14, 23, 8, 7, 33, 21, 3, 29, 14,
    -- filter=0 channel=54
    5, -4, -5, -8, -6, 8, -12, 2, 2,
    -- filter=0 channel=55
    10, -6, 3, 0, 1, -6, -4, 10, -1,
    -- filter=0 channel=56
    0, 0, -1, -9, -7, -7, 1, 8, -7,
    -- filter=0 channel=57
    -2, -8, -4, 3, 9, 9, -2, -6, -8,
    -- filter=0 channel=58
    13, 14, 0, 11, 14, 5, 2, 10, 0,
    -- filter=0 channel=59
    5, 11, 12, 5, 10, 12, 8, 8, 12,
    -- filter=0 channel=60
    -24, -19, -17, -20, -29, -15, -22, -25, -32,
    -- filter=0 channel=61
    -8, -5, -5, -19, -19, -20, -14, -21, -7,
    -- filter=0 channel=62
    3, 13, 2, 5, 16, 1, -5, -5, 11,
    -- filter=0 channel=63
    8, -3, -4, 3, 0, -3, -4, 4, 3,
    -- filter=1 channel=0
    -5, 6, -8, -5, 9, -10, 8, 8, -3,
    -- filter=1 channel=1
    19, 13, 10, 21, 35, 25, 19, 33, 10,
    -- filter=1 channel=2
    13, 20, 23, 28, 39, 16, 22, 22, 28,
    -- filter=1 channel=3
    0, 13, 7, 1, 18, 3, 10, 19, 4,
    -- filter=1 channel=4
    4, -10, -5, -4, -16, -14, 2, -4, -11,
    -- filter=1 channel=5
    -9, 3, 0, 7, -5, -5, -4, -3, -4,
    -- filter=1 channel=6
    6, -1, 6, 12, 8, 5, 13, 4, 7,
    -- filter=1 channel=7
    -6, 2, 0, -8, 5, -3, 4, 2, 12,
    -- filter=1 channel=8
    -14, -10, -6, 0, 0, -3, -4, -8, -5,
    -- filter=1 channel=9
    -14, -24, -13, -17, -36, -18, -22, -30, -20,
    -- filter=1 channel=10
    0, 5, 8, -1, 13, 5, 12, 23, 20,
    -- filter=1 channel=11
    -6, 3, -10, 9, 16, -9, 2, 4, -3,
    -- filter=1 channel=12
    6, 4, -1, -1, 0, 0, 1, 9, -5,
    -- filter=1 channel=13
    -12, -21, -17, -10, -17, -16, 0, -3, -6,
    -- filter=1 channel=14
    -8, 10, 7, 6, -6, -1, -3, 4, 7,
    -- filter=1 channel=15
    -2, -13, 0, -10, -11, 3, -3, -2, -8,
    -- filter=1 channel=16
    0, -5, -6, 4, 0, -2, -8, 11, 16,
    -- filter=1 channel=17
    -6, -3, -5, -6, -6, -15, -4, 7, 0,
    -- filter=1 channel=18
    -4, -23, -7, -23, -14, -14, -19, -13, -7,
    -- filter=1 channel=19
    10, 23, 13, 15, 17, 5, 9, 3, 8,
    -- filter=1 channel=20
    9, 4, -4, 10, 4, 0, 11, -1, 13,
    -- filter=1 channel=21
    1, -9, 10, 8, 8, 2, 9, 0, -7,
    -- filter=1 channel=22
    0, 5, 10, -7, 6, 7, 3, -2, -10,
    -- filter=1 channel=23
    13, 21, -3, 5, 27, 17, 8, 12, -3,
    -- filter=1 channel=24
    -20, -9, -1, -2, -4, -13, -10, -15, -12,
    -- filter=1 channel=25
    26, 28, 12, 34, 55, 32, 27, 40, 33,
    -- filter=1 channel=26
    5, 6, 17, 12, 7, 16, 22, 4, 4,
    -- filter=1 channel=27
    -2, 12, 11, 15, 29, 20, 10, 15, 17,
    -- filter=1 channel=28
    3, -10, -11, 5, -1, -9, -6, 3, 8,
    -- filter=1 channel=29
    -1, -10, -13, 0, 1, -3, -8, 4, -1,
    -- filter=1 channel=30
    17, 24, 15, 19, 30, 23, 13, 19, 20,
    -- filter=1 channel=31
    -5, 2, 3, -6, 10, 0, -3, 4, 4,
    -- filter=1 channel=32
    19, 13, 17, 23, 39, 14, 10, 33, 10,
    -- filter=1 channel=33
    -7, -5, -9, -3, 5, -2, -8, -9, -1,
    -- filter=1 channel=34
    -1, -4, 8, -1, 4, -6, 6, -4, 5,
    -- filter=1 channel=35
    8, 35, 15, 24, 35, 27, 26, 27, 23,
    -- filter=1 channel=36
    -1, 4, 0, 10, -4, 14, 10, 8, 10,
    -- filter=1 channel=37
    5, 0, -7, 0, -5, 0, -4, 5, 5,
    -- filter=1 channel=38
    -8, 6, 2, 18, 18, -3, 5, 21, 2,
    -- filter=1 channel=39
    -5, 7, 9, -9, 8, 10, 5, 10, 7,
    -- filter=1 channel=40
    4, 16, 13, 0, 0, 4, -5, 10, 2,
    -- filter=1 channel=41
    -1, -8, -4, -6, 15, 12, -8, 0, 6,
    -- filter=1 channel=42
    -6, -6, 4, -9, 9, -2, -4, 0, -9,
    -- filter=1 channel=43
    11, 17, 25, 23, 27, 22, 25, 37, 29,
    -- filter=1 channel=44
    16, 13, 14, 23, 25, 23, 18, 27, 17,
    -- filter=1 channel=45
    -6, -4, -4, 10, 2, 3, 1, 0, -5,
    -- filter=1 channel=46
    9, -1, 12, 5, 3, 0, -4, 0, 13,
    -- filter=1 channel=47
    8, 0, 6, -9, 2, -3, 0, -5, 10,
    -- filter=1 channel=48
    3, -10, -7, -3, 8, 7, 1, 6, 1,
    -- filter=1 channel=49
    4, 6, 0, 4, 19, 4, 3, 8, 9,
    -- filter=1 channel=50
    2, 24, 19, 14, 26, 25, 15, 4, 20,
    -- filter=1 channel=51
    -5, -14, 0, -6, -9, 0, -12, 2, 0,
    -- filter=1 channel=52
    3, -3, -1, 8, -1, -7, -1, -9, -3,
    -- filter=1 channel=53
    15, 27, 13, 20, 30, 33, 14, 20, 22,
    -- filter=1 channel=54
    0, -14, -6, -22, -23, -17, -18, -25, -12,
    -- filter=1 channel=55
    4, -8, -4, -9, -3, 8, -9, 8, 5,
    -- filter=1 channel=56
    0, 0, 5, 13, -6, 0, 3, 6, -5,
    -- filter=1 channel=57
    4, 10, 2, 6, -6, -10, -4, -1, 6,
    -- filter=1 channel=58
    0, 2, 16, 16, 5, 12, -1, 2, 14,
    -- filter=1 channel=59
    1, 6, 2, 7, 26, 5, 0, 19, 20,
    -- filter=1 channel=60
    -16, -12, -26, -7, -15, -20, -8, -18, -18,
    -- filter=1 channel=61
    -11, -17, -9, -8, 4, -15, -5, -6, -14,
    -- filter=1 channel=62
    9, 9, 4, 14, 16, -6, 11, 14, -4,
    -- filter=1 channel=63
    -9, 4, -2, 0, 0, -1, -5, -2, 9,
    -- filter=2 channel=0
    -5, -8, 2, 6, 0, -4, -3, 1, -3,
    -- filter=2 channel=1
    0, -5, 3, 1, 1, -1, -8, 5, -4,
    -- filter=2 channel=2
    -15, -9, -4, 6, -4, -5, 8, 3, 10,
    -- filter=2 channel=3
    0, 7, -8, -6, -3, 11, 2, -5, 4,
    -- filter=2 channel=4
    -2, 0, -10, 7, 3, 0, 11, 10, 7,
    -- filter=2 channel=5
    0, -1, 9, 1, 0, 7, 1, 8, 8,
    -- filter=2 channel=6
    -10, -6, -1, 5, 9, 4, 1, -8, 11,
    -- filter=2 channel=7
    -4, 5, -10, 2, 0, 6, 9, 7, 6,
    -- filter=2 channel=8
    -11, -1, -12, -2, 5, 6, 16, 1, 1,
    -- filter=2 channel=9
    4, -5, 3, 6, -5, 2, -1, 7, 0,
    -- filter=2 channel=10
    8, 0, 1, 6, 0, -5, 9, -4, 5,
    -- filter=2 channel=11
    -6, -10, -13, -9, 8, 7, -2, 10, 13,
    -- filter=2 channel=12
    -1, 4, 0, 7, -7, 7, -2, 5, -2,
    -- filter=2 channel=13
    5, 0, 4, -11, -1, -11, 8, 2, 3,
    -- filter=2 channel=14
    4, 1, 8, 6, -8, -4, -3, -2, 9,
    -- filter=2 channel=15
    0, -8, -3, 12, 11, -5, 3, 1, 0,
    -- filter=2 channel=16
    -7, -18, -15, -3, 3, -5, 6, 2, 0,
    -- filter=2 channel=17
    -10, -10, 5, -4, 0, -9, 7, 15, 12,
    -- filter=2 channel=18
    -1, -1, -6, 9, -2, -5, -2, 9, -2,
    -- filter=2 channel=19
    6, 3, -4, 1, -6, 8, 3, -8, 2,
    -- filter=2 channel=20
    -5, 5, 7, -2, -6, 12, 1, 5, 1,
    -- filter=2 channel=21
    -9, -4, -9, 0, 10, 0, -3, 6, -3,
    -- filter=2 channel=22
    10, 0, 0, 9, 5, 1, 0, 7, -8,
    -- filter=2 channel=23
    -5, -1, 1, 4, -7, -11, 6, 6, 5,
    -- filter=2 channel=24
    5, -1, 3, -10, -7, -6, -7, 12, -1,
    -- filter=2 channel=25
    2, -11, -2, -8, -13, -8, -6, 6, 7,
    -- filter=2 channel=26
    -2, 3, 0, -7, -5, 5, 11, 3, 2,
    -- filter=2 channel=27
    -11, -11, -8, -4, 5, -1, -5, 16, 9,
    -- filter=2 channel=28
    -6, 0, -1, -3, 7, -7, 0, 11, 9,
    -- filter=2 channel=29
    -7, -14, -3, -9, -8, -3, 15, 18, 15,
    -- filter=2 channel=30
    -5, -4, -7, 1, -2, -6, 7, -8, 0,
    -- filter=2 channel=31
    9, 11, 0, 3, 0, -7, 1, 9, 6,
    -- filter=2 channel=32
    -9, -5, -8, -12, -7, -11, -9, 0, 7,
    -- filter=2 channel=33
    -3, 3, 7, 10, 2, -1, 5, -1, -9,
    -- filter=2 channel=34
    -2, -2, -9, 4, -1, 3, 10, 0, 6,
    -- filter=2 channel=35
    -13, -1, 4, 2, -2, 0, -7, -3, 0,
    -- filter=2 channel=36
    3, -5, -9, -4, 0, -5, 9, 0, 0,
    -- filter=2 channel=37
    4, 1, 8, -7, 2, -4, 0, -4, 8,
    -- filter=2 channel=38
    -15, -13, -7, 0, 4, 5, -1, 14, 3,
    -- filter=2 channel=39
    -9, -4, 1, 9, 5, 3, 5, 8, 3,
    -- filter=2 channel=40
    4, -5, 5, -8, -6, -6, 8, 8, 10,
    -- filter=2 channel=41
    -10, -14, -8, 2, -1, 7, 18, 11, 18,
    -- filter=2 channel=42
    3, 4, -7, 9, 2, 0, 9, 6, -3,
    -- filter=2 channel=43
    -3, 11, 3, -1, -4, -4, -2, -6, -4,
    -- filter=2 channel=44
    -6, -1, -9, 9, 11, 7, 3, 4, 7,
    -- filter=2 channel=45
    -8, -2, -2, 2, 9, -2, 4, -8, -7,
    -- filter=2 channel=46
    -1, -1, 7, 0, 0, 9, -1, -1, -6,
    -- filter=2 channel=47
    4, -6, 8, -3, -6, -5, 2, -9, -2,
    -- filter=2 channel=48
    -11, -8, -4, 0, 0, 0, 1, -1, -1,
    -- filter=2 channel=49
    -9, -2, -8, 1, 2, 12, -2, 4, -2,
    -- filter=2 channel=50
    2, 0, 7, 5, 10, 6, -1, 0, 8,
    -- filter=2 channel=51
    -8, 5, -2, 8, -8, 4, 11, 3, 4,
    -- filter=2 channel=52
    6, -2, 0, 6, -10, -7, -3, -7, -6,
    -- filter=2 channel=53
    7, -7, -9, -6, 8, 6, 2, 2, -1,
    -- filter=2 channel=54
    0, 9, 3, 8, 2, 2, 6, -4, 5,
    -- filter=2 channel=55
    -8, -8, -8, 1, -2, -9, 5, 9, -10,
    -- filter=2 channel=56
    -9, -4, 4, 4, -2, -6, 5, 1, -8,
    -- filter=2 channel=57
    5, 0, 7, -5, -3, 0, 9, -8, -1,
    -- filter=2 channel=58
    6, 0, -3, 5, 6, -5, 1, -8, -8,
    -- filter=2 channel=59
    -7, 1, 1, 7, -12, -1, -2, 15, 16,
    -- filter=2 channel=60
    -7, -12, -9, 0, -7, 3, 22, 8, 22,
    -- filter=2 channel=61
    -2, -16, -4, 7, 0, -4, 10, 15, 19,
    -- filter=2 channel=62
    -8, 2, 4, -6, -9, -5, 1, 11, 11,
    -- filter=2 channel=63
    7, 0, 9, 6, -4, -5, 10, -3, 9,
    -- filter=3 channel=0
    5, 11, -3, 14, 8, 15, -3, -16, -3,
    -- filter=3 channel=1
    0, 5, 4, 9, 4, 14, -1, 0, -2,
    -- filter=3 channel=2
    18, 23, 10, -10, -4, -3, -20, -28, -26,
    -- filter=3 channel=3
    9, 14, 1, 7, 0, 1, 3, -8, 3,
    -- filter=3 channel=4
    6, 12, 5, -6, 0, 1, -14, -14, -14,
    -- filter=3 channel=5
    -1, 3, 11, 2, -12, -6, 5, -5, -7,
    -- filter=3 channel=6
    10, 16, 13, 6, -8, -6, -9, -3, -17,
    -- filter=3 channel=7
    1, 1, -3, -2, 0, 3, 0, -7, -5,
    -- filter=3 channel=8
    23, 23, 24, 10, -2, -8, -32, -40, -26,
    -- filter=3 channel=9
    10, 0, 2, -2, 17, 7, -10, 7, -3,
    -- filter=3 channel=10
    -3, -4, -13, 5, 15, 11, 9, 12, 9,
    -- filter=3 channel=11
    -5, 0, 15, 7, 6, 18, -13, -25, -26,
    -- filter=3 channel=12
    -2, -5, -7, -8, 6, 3, -3, -6, -3,
    -- filter=3 channel=13
    5, 5, 5, 11, 21, 11, -14, -12, -8,
    -- filter=3 channel=14
    -8, -8, -2, -6, 7, -5, 2, -8, -3,
    -- filter=3 channel=15
    32, 31, 11, 5, 1, -12, -12, -39, -18,
    -- filter=3 channel=16
    23, 35, 18, 10, 13, 2, -20, -41, -32,
    -- filter=3 channel=17
    8, 22, 27, 4, 0, -5, -15, -31, -30,
    -- filter=3 channel=18
    5, 13, 12, 4, 0, -10, -9, 4, -9,
    -- filter=3 channel=19
    0, -5, 9, 10, 0, -6, -3, -1, -12,
    -- filter=3 channel=20
    -4, 2, -9, -10, -7, 3, -9, 2, 8,
    -- filter=3 channel=21
    -9, -5, 6, 2, -7, 7, 4, 7, 5,
    -- filter=3 channel=22
    9, 10, -1, 8, 5, 6, 10, 0, 6,
    -- filter=3 channel=23
    -1, 1, 0, 16, 14, 7, 0, 7, -5,
    -- filter=3 channel=24
    -5, 15, 12, 0, 14, 11, -6, -9, -9,
    -- filter=3 channel=25
    26, 29, 3, 2, 2, -1, -12, -26, -14,
    -- filter=3 channel=26
    -4, -8, -1, 0, -6, 3, -12, -4, 12,
    -- filter=3 channel=27
    6, 30, 21, 9, -2, 4, -10, -21, -27,
    -- filter=3 channel=28
    20, 22, 19, -12, 1, -8, -14, -23, -12,
    -- filter=3 channel=29
    25, 30, 35, 14, 8, -5, -41, -50, -23,
    -- filter=3 channel=30
    -5, -12, -7, -12, 3, -7, 5, 1, -5,
    -- filter=3 channel=31
    -5, -10, 0, 9, 4, -5, 11, 1, 7,
    -- filter=3 channel=32
    7, 6, -3, -2, 0, -4, 11, -5, -3,
    -- filter=3 channel=33
    8, -4, -7, 4, -2, -4, 1, 10, -4,
    -- filter=3 channel=34
    -1, -11, 5, 2, 0, 1, 2, -11, -7,
    -- filter=3 channel=35
    2, 4, 10, 0, -7, 0, -6, -6, -2,
    -- filter=3 channel=36
    -10, -7, 1, -7, 8, 3, 11, 11, 12,
    -- filter=3 channel=37
    -2, 7, 17, -1, 18, 16, 2, -2, -8,
    -- filter=3 channel=38
    18, 18, 19, 11, 11, 3, -24, -32, -33,
    -- filter=3 channel=39
    10, 0, 2, -8, -9, -5, -4, -4, -3,
    -- filter=3 channel=40
    5, 15, 8, -1, -1, 8, 8, -11, 4,
    -- filter=3 channel=41
    30, 41, 34, -2, -6, 4, -38, -44, -34,
    -- filter=3 channel=42
    5, 8, 9, 5, -1, -8, -10, 3, 2,
    -- filter=3 channel=43
    18, 22, 25, 56, 67, 59, 13, 35, 23,
    -- filter=3 channel=44
    -6, -1, -3, -6, -4, -5, 1, 5, -8,
    -- filter=3 channel=45
    2, -4, 9, -9, 3, 7, 7, -7, 3,
    -- filter=3 channel=46
    -8, -8, -3, 2, 0, 4, -7, 5, 0,
    -- filter=3 channel=47
    10, -1, 3, -9, -1, 6, -1, -6, -6,
    -- filter=3 channel=48
    12, 9, 8, 0, -3, -9, -6, -5, -9,
    -- filter=3 channel=49
    23, 22, 7, -5, -15, -12, -11, -7, -17,
    -- filter=3 channel=50
    -1, -13, 9, -1, 17, 15, 10, -1, 0,
    -- filter=3 channel=51
    4, -1, 1, 6, 3, 8, 10, 8, -5,
    -- filter=3 channel=52
    2, 0, 2, -1, 7, -7, -5, 1, 9,
    -- filter=3 channel=53
    0, -12, -6, 1, -1, -1, 12, 12, 4,
    -- filter=3 channel=54
    0, 22, 15, -2, -1, 13, -5, -7, 4,
    -- filter=3 channel=55
    0, 7, 7, 3, 0, 9, 5, 0, -7,
    -- filter=3 channel=56
    -10, -3, 3, 11, -8, 9, 9, 3, 1,
    -- filter=3 channel=57
    5, -7, 1, -9, 0, 5, 0, -2, 4,
    -- filter=3 channel=58
    8, -9, 0, -3, 9, -10, -3, 5, 0,
    -- filter=3 channel=59
    11, 30, 23, 3, 10, 2, -22, -14, -9,
    -- filter=3 channel=60
    21, 22, 21, 19, 8, 2, -42, -46, -25,
    -- filter=3 channel=61
    13, 12, 21, 6, 16, 13, -25, -32, -31,
    -- filter=3 channel=62
    17, 21, 8, -1, 6, -1, -6, -6, -12,
    -- filter=3 channel=63
    -3, -1, -8, 7, 0, -6, 2, 9, 6,
    -- filter=4 channel=0
    -16, -16, -16, 4, -8, -7, 8, 20, 19,
    -- filter=4 channel=1
    6, 8, -13, -1, -12, -14, 4, 13, 3,
    -- filter=4 channel=2
    -6, -19, -26, -2, 2, 9, 7, 21, 8,
    -- filter=4 channel=3
    3, -14, 4, 10, -2, 14, 13, 12, 14,
    -- filter=4 channel=4
    -6, -15, -19, -4, 1, 0, 6, 21, 20,
    -- filter=4 channel=5
    5, -4, -11, 0, -4, 7, 0, 11, 11,
    -- filter=4 channel=6
    -12, -19, -1, -7, -3, 13, 15, 4, 6,
    -- filter=4 channel=7
    2, -5, -3, -10, -4, 6, -1, -1, -2,
    -- filter=4 channel=8
    -30, -40, -27, 8, -6, -2, 22, 29, 38,
    -- filter=4 channel=9
    2, -4, 8, -11, -1, 2, -8, 3, 13,
    -- filter=4 channel=10
    -7, 12, 3, -12, -10, -11, -5, 11, -3,
    -- filter=4 channel=11
    -13, -21, -16, 0, -7, 0, 0, 12, 26,
    -- filter=4 channel=12
    6, 11, -5, 0, 6, -6, -7, 9, -6,
    -- filter=4 channel=13
    -19, -16, -3, -14, -4, -17, 19, 13, 10,
    -- filter=4 channel=14
    9, -7, -12, -7, -6, -1, -11, 6, 1,
    -- filter=4 channel=15
    -14, -29, -33, 10, 7, 11, 30, 42, 19,
    -- filter=4 channel=16
    -18, -52, -48, -2, -12, 3, 16, 43, 46,
    -- filter=4 channel=17
    -6, -16, -36, 0, 7, 4, 21, 30, 38,
    -- filter=4 channel=18
    -12, -11, 7, -7, -3, 3, 2, 2, 10,
    -- filter=4 channel=19
    3, -6, -6, 0, 5, -8, 1, -3, 0,
    -- filter=4 channel=20
    -1, 6, 3, 5, -2, -1, 0, 2, -4,
    -- filter=4 channel=21
    -1, -4, 10, 10, 2, -1, 4, 1, -6,
    -- filter=4 channel=22
    3, -4, -5, 4, 4, 4, 5, 11, -6,
    -- filter=4 channel=23
    2, -1, -10, 9, -10, 0, -2, 8, 15,
    -- filter=4 channel=24
    8, -14, -5, -9, -5, -4, -3, 9, 26,
    -- filter=4 channel=25
    -18, -23, -27, 3, 12, 10, 6, 11, 11,
    -- filter=4 channel=26
    2, -3, 13, -2, -9, 3, 0, -5, -2,
    -- filter=4 channel=27
    -15, -29, -33, 7, 0, 6, 17, 36, 33,
    -- filter=4 channel=28
    -6, -14, -33, 3, 17, -1, 16, 9, 35,
    -- filter=4 channel=29
    -37, -58, -29, 2, 0, 2, 21, 45, 49,
    -- filter=4 channel=30
    2, 8, -5, 7, 1, 0, -2, -4, 13,
    -- filter=4 channel=31
    -9, 7, 0, 9, 3, -9, -6, 5, 1,
    -- filter=4 channel=32
    14, -2, 7, 10, 8, -8, -9, 9, 1,
    -- filter=4 channel=33
    0, 9, -2, 3, -3, -8, 9, -6, -9,
    -- filter=4 channel=34
    -8, 3, -9, -1, -6, -9, -7, -2, 5,
    -- filter=4 channel=35
    -10, -26, -19, 4, 14, -1, 4, 2, 10,
    -- filter=4 channel=36
    9, 2, 0, 8, 7, 4, 7, -8, -2,
    -- filter=4 channel=37
    0, -14, -14, -10, -6, -9, 17, 21, 22,
    -- filter=4 channel=38
    -8, -38, -30, -17, -10, -2, 17, 38, 31,
    -- filter=4 channel=39
    -3, 0, 10, 1, 7, 0, -8, 0, -2,
    -- filter=4 channel=40
    1, 8, -6, 10, 12, 15, -1, 16, 0,
    -- filter=4 channel=41
    -37, -53, -49, 4, 3, 20, 32, 42, 48,
    -- filter=4 channel=42
    2, -3, -6, 5, 6, 8, 9, -3, 7,
    -- filter=4 channel=43
    29, 39, 37, 21, 9, 9, 31, 26, 34,
    -- filter=4 channel=44
    0, -8, -12, 2, 4, 0, -1, -7, -3,
    -- filter=4 channel=45
    -9, -3, 2, -7, 0, -6, 1, -4, 0,
    -- filter=4 channel=46
    -13, 0, 8, 0, 10, 0, 1, -1, 0,
    -- filter=4 channel=47
    0, 3, 2, 10, 8, 0, -6, -1, -3,
    -- filter=4 channel=48
    -16, -21, -1, 2, 2, -1, 2, 7, 16,
    -- filter=4 channel=49
    -8, -12, -12, 12, 16, 31, 17, 17, 14,
    -- filter=4 channel=50
    16, 22, 9, -12, 0, 0, -10, 7, 8,
    -- filter=4 channel=51
    9, 6, -5, 1, -8, 5, 2, -8, -6,
    -- filter=4 channel=52
    7, -6, -4, 5, -4, 2, -8, 3, 6,
    -- filter=4 channel=53
    0, 14, -1, 0, 8, -2, 0, 2, 14,
    -- filter=4 channel=54
    -12, 0, -5, 0, 14, 7, 10, 12, 23,
    -- filter=4 channel=55
    -7, -2, -9, 5, 1, 9, 3, 6, -10,
    -- filter=4 channel=56
    10, 9, 2, -3, -9, -10, 4, 9, -2,
    -- filter=4 channel=57
    -8, 9, -8, -1, 8, 2, -1, -3, -9,
    -- filter=4 channel=58
    1, 10, 14, -1, 11, -2, -9, -8, -2,
    -- filter=4 channel=59
    -29, -38, -31, 10, -10, -3, 18, 34, 30,
    -- filter=4 channel=60
    -39, -53, -42, -6, -10, -3, 29, 54, 39,
    -- filter=4 channel=61
    -9, -24, -37, -13, -7, -1, 14, 26, 28,
    -- filter=4 channel=62
    -12, -22, -23, -7, 8, -7, 10, 26, 11,
    -- filter=4 channel=63
    2, 1, -3, -8, -10, -2, 3, 8, 2,
    -- filter=5 channel=0
    14, 7, 12, 5, 19, 21, -5, 7, -1,
    -- filter=5 channel=1
    12, 14, 16, 3, 27, 16, 9, 14, 9,
    -- filter=5 channel=2
    9, 10, 22, 1, 4, 5, 4, 10, 5,
    -- filter=5 channel=3
    0, 5, 16, 8, 3, 10, 9, 4, 12,
    -- filter=5 channel=4
    4, -5, -11, 3, -15, -7, 0, 1, -1,
    -- filter=5 channel=5
    -15, 0, -11, -5, -10, 1, 2, -6, -2,
    -- filter=5 channel=6
    -3, 14, 12, -5, 6, 14, 5, 11, 9,
    -- filter=5 channel=7
    -11, 3, 6, -3, -7, -9, -8, 0, -4,
    -- filter=5 channel=8
    -15, -9, -3, -9, -5, -13, -17, -14, -19,
    -- filter=5 channel=9
    -7, -28, -19, -14, -19, -19, -3, -20, -19,
    -- filter=5 channel=10
    2, 20, 21, 11, 30, 18, 0, 27, 20,
    -- filter=5 channel=11
    -5, 2, 11, -5, -4, 6, 4, 0, -3,
    -- filter=5 channel=12
    4, 3, -5, 10, -6, 1, 4, 6, -1,
    -- filter=5 channel=13
    -7, -9, -2, 2, -10, -15, -7, -4, -15,
    -- filter=5 channel=14
    -14, 0, -3, -4, -6, 4, -8, 4, 1,
    -- filter=5 channel=15
    3, -4, -7, -21, -17, -7, -9, -19, -14,
    -- filter=5 channel=16
    -11, -3, 8, -8, -21, 0, -13, -20, -6,
    -- filter=5 channel=17
    -5, -2, 10, -2, -12, -5, -4, 0, -2,
    -- filter=5 channel=18
    6, -6, -8, 1, -12, -9, -6, -20, -15,
    -- filter=5 channel=19
    -13, -5, -5, -11, -5, 1, -2, 4, 0,
    -- filter=5 channel=20
    5, -13, 4, 4, -13, -12, -1, 4, -10,
    -- filter=5 channel=21
    -1, -7, -4, 3, -8, -8, 10, 3, -7,
    -- filter=5 channel=22
    -10, 3, 6, -7, 10, 7, 0, -7, -2,
    -- filter=5 channel=23
    15, 33, 30, 26, 31, 34, 18, 20, 21,
    -- filter=5 channel=24
    -15, -9, 4, -1, -4, 0, -16, -5, -8,
    -- filter=5 channel=25
    15, 33, 24, 4, 23, 31, 9, 29, 22,
    -- filter=5 channel=26
    11, 5, 7, 7, 9, 11, -3, -6, 2,
    -- filter=5 channel=27
    3, 23, 19, 6, 22, 17, 18, 18, 18,
    -- filter=5 channel=28
    -12, -15, -20, -14, -29, -20, -16, -19, -20,
    -- filter=5 channel=29
    -24, -14, 0, -15, -30, -8, -26, -32, -22,
    -- filter=5 channel=30
    -11, 3, -8, -8, -5, -2, 0, -4, 6,
    -- filter=5 channel=31
    11, 6, 4, 12, 5, -2, 0, 0, 9,
    -- filter=5 channel=32
    20, 27, 21, 17, 36, 32, 5, 30, 14,
    -- filter=5 channel=33
    5, 0, 8, -7, 1, -3, 0, 8, -1,
    -- filter=5 channel=34
    5, -10, -3, -8, -10, 1, -9, 3, -11,
    -- filter=5 channel=35
    29, 49, 37, 15, 55, 41, 29, 30, 38,
    -- filter=5 channel=36
    9, 10, 7, 4, 9, 1, 1, 11, 6,
    -- filter=5 channel=37
    -1, 4, 4, -4, 5, 0, -11, -12, 1,
    -- filter=5 channel=38
    6, 24, 20, -3, 25, 15, -5, 7, 9,
    -- filter=5 channel=39
    10, 2, 8, 10, -6, 0, 8, -3, 5,
    -- filter=5 channel=40
    -6, 8, 12, 5, 14, 5, -5, 0, 15,
    -- filter=5 channel=41
    7, -2, 14, -6, 6, 8, 2, -5, -3,
    -- filter=5 channel=42
    6, 6, -5, -8, 3, 0, 3, 3, 1,
    -- filter=5 channel=43
    -2, 9, 7, 12, 21, 10, -1, 5, 11,
    -- filter=5 channel=44
    9, 20, 8, 7, 7, 22, 20, 15, 16,
    -- filter=5 channel=45
    0, 1, -1, -1, -4, -5, 0, 9, -4,
    -- filter=5 channel=46
    1, -2, 1, -7, -4, 0, -11, -13, -7,
    -- filter=5 channel=47
    -7, 10, -3, 6, 3, -4, 3, -9, 6,
    -- filter=5 channel=48
    -14, 1, -8, 2, -6, -11, -3, -1, 0,
    -- filter=5 channel=49
    8, 17, 15, -2, 17, 1, 12, 15, 16,
    -- filter=5 channel=50
    1, 0, -9, -12, -9, -8, 0, -5, -5,
    -- filter=5 channel=51
    6, 2, 9, 1, 7, 15, 14, 17, 11,
    -- filter=5 channel=52
    7, 0, 6, -6, -8, -7, -9, 5, -9,
    -- filter=5 channel=53
    -2, -2, 4, 1, 2, 13, 7, 11, 5,
    -- filter=5 channel=54
    -8, -7, 5, -3, -14, -9, -3, -1, 0,
    -- filter=5 channel=55
    9, 1, 9, 0, 6, -9, -4, 6, 4,
    -- filter=5 channel=56
    6, 8, -11, 8, -1, 2, 3, -7, 8,
    -- filter=5 channel=57
    5, 10, -8, 1, -3, 3, -4, -9, -7,
    -- filter=5 channel=58
    10, 0, -6, -3, 5, 3, -1, -7, 6,
    -- filter=5 channel=59
    3, 6, 12, -4, 6, 4, -4, 5, 2,
    -- filter=5 channel=60
    -1, 4, -6, -11, -9, 6, -13, -12, -11,
    -- filter=5 channel=61
    -7, 4, -2, 0, -7, 6, -11, -4, 2,
    -- filter=5 channel=62
    -7, 5, 7, 0, -3, -8, 1, -2, -1,
    -- filter=5 channel=63
    10, 0, -1, 1, 6, -1, -7, 3, -5,
    -- filter=6 channel=0
    1, 0, -13, -12, -13, -13, -5, -3, -3,
    -- filter=6 channel=1
    5, 13, 6, 5, 15, -2, 5, 1, 14,
    -- filter=6 channel=2
    2, 0, -3, 8, 11, 16, 10, 12, 12,
    -- filter=6 channel=3
    0, -3, 3, 2, 15, 14, 13, 8, 3,
    -- filter=6 channel=4
    -1, -9, 4, 3, -8, -12, 6, 0, 2,
    -- filter=6 channel=5
    11, 5, 8, 3, 0, 12, 13, -4, 1,
    -- filter=6 channel=6
    6, -2, -5, -6, 7, 9, 2, -7, -9,
    -- filter=6 channel=7
    6, 9, 0, 11, 10, 9, 9, 9, 0,
    -- filter=6 channel=8
    -5, -11, -7, -13, -16, 4, -12, -2, -5,
    -- filter=6 channel=9
    3, 14, 22, 8, 36, 32, 18, 15, 12,
    -- filter=6 channel=10
    6, 0, 9, -2, 1, -5, -8, 1, -3,
    -- filter=6 channel=11
    0, -6, -10, -8, -1, 3, -10, 2, -2,
    -- filter=6 channel=12
    -4, 6, -5, 9, 6, -9, 4, 4, -7,
    -- filter=6 channel=13
    -13, -3, 5, 6, 11, 11, -7, 0, 7,
    -- filter=6 channel=14
    2, 9, -8, 4, 7, 7, -2, -2, -6,
    -- filter=6 channel=15
    -13, -6, -6, -13, 7, 1, -6, -8, -10,
    -- filter=6 channel=16
    -8, -7, -2, 7, 4, 12, 7, -7, 0,
    -- filter=6 channel=17
    -7, -8, -7, -4, -7, -9, 9, -5, -9,
    -- filter=6 channel=18
    -4, 1, -2, -5, -7, -9, -10, 0, 7,
    -- filter=6 channel=19
    3, 1, 13, 12, 16, 13, 6, 3, -3,
    -- filter=6 channel=20
    2, 17, 0, 9, 3, 5, 3, 12, 0,
    -- filter=6 channel=21
    10, 10, -2, 10, 9, 10, -3, 12, 10,
    -- filter=6 channel=22
    4, -3, -2, 0, -2, -3, -1, 0, -1,
    -- filter=6 channel=23
    1, -5, -13, 8, -6, 0, 3, -5, 3,
    -- filter=6 channel=24
    -2, -6, 3, -5, -2, -3, 3, -9, 7,
    -- filter=6 channel=25
    3, 2, 10, 11, 0, 3, 12, 9, 4,
    -- filter=6 channel=26
    8, 6, 6, 10, 8, 13, 11, 6, 0,
    -- filter=6 channel=27
    -2, -10, 3, 3, -7, -2, 2, -1, 0,
    -- filter=6 channel=28
    0, 2, 8, -7, -1, 0, -6, 5, 10,
    -- filter=6 channel=29
    2, 6, 13, 5, 1, 5, 6, 3, -10,
    -- filter=6 channel=30
    -1, 12, 12, 8, 7, 13, 7, 4, 1,
    -- filter=6 channel=31
    5, -8, 3, 11, 0, 11, 3, 2, -7,
    -- filter=6 channel=32
    4, 13, 12, 5, 16, 10, 7, 16, 2,
    -- filter=6 channel=33
    -3, -7, -2, -1, 0, 8, 5, -1, 6,
    -- filter=6 channel=34
    3, -3, 7, 6, 11, 3, -7, 2, 6,
    -- filter=6 channel=35
    -8, -10, 1, 0, 5, -3, -1, -7, -9,
    -- filter=6 channel=36
    8, 7, 0, 5, 5, -5, 3, -1, -1,
    -- filter=6 channel=37
    -4, 11, 13, 4, 5, 17, 13, 11, 8,
    -- filter=6 channel=38
    -7, -6, 0, -1, 0, 2, -5, -7, 0,
    -- filter=6 channel=39
    -4, -8, -3, 5, 9, -9, -3, 1, -3,
    -- filter=6 channel=40
    -5, -7, 6, -1, 8, 1, -8, -1, -9,
    -- filter=6 channel=41
    2, 1, 2, 7, 8, -10, -9, -6, -4,
    -- filter=6 channel=42
    5, 8, -2, 4, 6, -9, -6, -10, -10,
    -- filter=6 channel=43
    -9, 5, -2, -4, -9, -3, 7, 5, -3,
    -- filter=6 channel=44
    -4, 12, 10, 17, -3, 6, 9, 8, -4,
    -- filter=6 channel=45
    -3, 1, -5, -3, -5, 7, 10, -10, -8,
    -- filter=6 channel=46
    11, 5, -3, -5, 4, 9, -7, -1, -1,
    -- filter=6 channel=47
    -2, 9, -1, -5, 2, 4, 0, 2, -8,
    -- filter=6 channel=48
    -10, 7, 8, 1, -4, 11, -7, -6, 0,
    -- filter=6 channel=49
    -7, 1, -3, 3, -11, -13, 9, 4, -2,
    -- filter=6 channel=50
    4, -2, -4, 0, 11, 15, -1, 9, 12,
    -- filter=6 channel=51
    -3, -15, -11, 6, 0, -10, -3, 2, -6,
    -- filter=6 channel=52
    0, 3, -1, -8, 1, -7, 3, -8, 5,
    -- filter=6 channel=53
    16, 12, 3, 12, 15, 0, 2, 6, 14,
    -- filter=6 channel=54
    11, 6, 25, 17, 31, 13, 11, 9, 15,
    -- filter=6 channel=55
    0, -4, 7, 6, -5, 8, 0, 5, 1,
    -- filter=6 channel=56
    9, 3, -4, -8, -5, -6, 4, 5, 6,
    -- filter=6 channel=57
    -2, -4, -6, -5, -5, 7, 8, -5, -8,
    -- filter=6 channel=58
    -3, 9, 13, 11, 1, 6, 13, 3, -6,
    -- filter=6 channel=59
    -6, -4, 3, 0, 8, 8, 9, 2, -4,
    -- filter=6 channel=60
    -6, -15, 0, -16, -3, 3, 3, -1, 2,
    -- filter=6 channel=61
    -16, -4, -18, 3, -5, -13, -8, -14, -8,
    -- filter=6 channel=62
    10, -5, 4, 10, 3, -1, 1, -2, 11,
    -- filter=6 channel=63
    -9, 9, -9, 7, -8, 1, -3, -4, -2,
    -- filter=7 channel=0
    -4, -3, 4, -8, -2, 4, -9, -2, -2,
    -- filter=7 channel=1
    4, 8, -10, 2, -10, -7, -3, -5, 8,
    -- filter=7 channel=2
    2, -5, 4, 0, 3, 0, 7, -4, -7,
    -- filter=7 channel=3
    5, -2, -4, -1, 6, -10, 0, -9, -10,
    -- filter=7 channel=4
    -3, -10, 0, -5, 0, -7, 10, -10, -1,
    -- filter=7 channel=5
    -7, 0, -9, -5, 7, 9, -2, -2, -2,
    -- filter=7 channel=6
    2, 10, -2, -8, -1, 2, 8, 9, 6,
    -- filter=7 channel=7
    -10, -4, -8, -8, 6, -7, 5, 2, -2,
    -- filter=7 channel=8
    -1, -3, 9, 2, 2, 8, 1, 7, 1,
    -- filter=7 channel=9
    -8, 8, -2, -7, -8, 0, -3, 1, -6,
    -- filter=7 channel=10
    -7, -6, 0, -1, -3, 0, 10, 4, 0,
    -- filter=7 channel=11
    7, 1, 5, 0, 0, -6, -5, -8, 7,
    -- filter=7 channel=12
    -9, 0, 4, 10, 4, -7, -5, -8, -2,
    -- filter=7 channel=13
    7, -9, -4, -7, -8, -2, 5, -2, 1,
    -- filter=7 channel=14
    9, 4, 7, -2, 7, -2, 1, -2, 6,
    -- filter=7 channel=15
    6, 7, -1, 4, -3, -8, 9, 10, 10,
    -- filter=7 channel=16
    -3, -5, -10, 1, 2, -9, 9, -9, 9,
    -- filter=7 channel=17
    -3, -6, 5, 8, -8, 3, -1, -10, 4,
    -- filter=7 channel=18
    3, 7, 6, 9, -8, 0, 8, 6, -7,
    -- filter=7 channel=19
    -3, 0, 6, -1, 4, -5, 6, 5, 4,
    -- filter=7 channel=20
    -3, 6, -8, -6, -9, 2, 8, 2, 4,
    -- filter=7 channel=21
    7, 2, 1, -6, 9, -2, 10, -5, -3,
    -- filter=7 channel=22
    9, 10, 0, -1, -5, 0, 6, 9, -6,
    -- filter=7 channel=23
    -9, -4, -2, -5, -9, -5, -6, -5, -10,
    -- filter=7 channel=24
    -4, -7, -10, -2, 4, 9, -9, 5, 0,
    -- filter=7 channel=25
    -5, 6, -2, -8, 2, -2, 9, 10, -7,
    -- filter=7 channel=26
    0, 5, -7, -2, 4, -6, -8, -2, 3,
    -- filter=7 channel=27
    9, 5, 5, 9, 0, 8, -3, 7, -4,
    -- filter=7 channel=28
    -3, 1, -1, 8, 5, 8, 4, 9, 0,
    -- filter=7 channel=29
    -6, 5, 0, -10, -1, 8, 3, -2, -10,
    -- filter=7 channel=30
    -3, 0, 6, 0, 8, 1, -1, -8, -7,
    -- filter=7 channel=31
    4, 6, 0, -9, 6, -5, 8, -5, 9,
    -- filter=7 channel=32
    -5, 5, -4, -10, -4, -2, -1, 9, 7,
    -- filter=7 channel=33
    -1, 1, -3, 2, -10, -2, 0, 0, 2,
    -- filter=7 channel=34
    2, 9, 2, 10, -4, -8, -3, 6, 2,
    -- filter=7 channel=35
    -4, 3, 3, -7, 4, -10, 8, -7, -2,
    -- filter=7 channel=36
    -3, -3, -8, -9, 6, 5, 4, -3, 9,
    -- filter=7 channel=37
    -3, 10, 6, -6, 10, 7, -9, 1, 5,
    -- filter=7 channel=38
    -5, 6, -2, 8, -3, 4, -10, -7, 3,
    -- filter=7 channel=39
    1, 9, 1, -8, 10, -10, 7, -5, -5,
    -- filter=7 channel=40
    5, -5, -7, -1, 0, -7, 8, -5, 4,
    -- filter=7 channel=41
    -9, 8, 2, 4, -2, -7, -1, -3, -6,
    -- filter=7 channel=42
    -10, -4, 8, -3, -4, 9, 2, -6, -4,
    -- filter=7 channel=43
    -5, -2, -8, 5, 7, 8, 0, 3, -10,
    -- filter=7 channel=44
    3, -2, -4, 0, 10, 5, 4, 1, 7,
    -- filter=7 channel=45
    -8, -10, 5, -8, 3, 4, 9, 0, -8,
    -- filter=7 channel=46
    -7, 0, -2, -9, -8, 8, 8, -9, 9,
    -- filter=7 channel=47
    0, 9, -5, -2, 6, -1, 8, -9, -1,
    -- filter=7 channel=48
    4, 7, -4, 9, 0, 10, 0, -9, 9,
    -- filter=7 channel=49
    -8, 2, -6, 1, -7, -6, -6, 7, -2,
    -- filter=7 channel=50
    -8, 2, -4, -7, -5, 5, -8, 4, 5,
    -- filter=7 channel=51
    -3, 3, 3, 7, -8, -8, -1, 8, -3,
    -- filter=7 channel=52
    10, -6, -6, -6, -5, 9, -10, 0, 10,
    -- filter=7 channel=53
    -7, -7, 0, 6, 10, 0, -5, -9, -4,
    -- filter=7 channel=54
    -4, -3, 7, 7, -8, 7, -2, -3, 7,
    -- filter=7 channel=55
    0, 0, 3, -1, 0, 3, -4, 0, -8,
    -- filter=7 channel=56
    7, -2, 5, -3, -6, 8, 2, 8, -8,
    -- filter=7 channel=57
    -6, -6, 9, 6, 9, -2, 6, 0, -5,
    -- filter=7 channel=58
    -10, -3, 3, -7, -7, 8, 2, -1, -10,
    -- filter=7 channel=59
    5, 6, 0, -7, 3, 8, 0, 9, 3,
    -- filter=7 channel=60
    0, -9, 1, -10, -8, -10, -1, 1, -8,
    -- filter=7 channel=61
    3, -7, -1, -9, 7, 5, 0, 0, -9,
    -- filter=7 channel=62
    7, 0, 9, -6, 0, -7, -7, 0, 3,
    -- filter=7 channel=63
    -4, 5, -5, -10, -2, -4, 1, 3, -9,
    -- filter=8 channel=0
    -7, -3, -6, -15, 0, 0, -6, 12, 15,
    -- filter=8 channel=1
    0, 5, 9, 0, -15, 4, -14, -10, 5,
    -- filter=8 channel=2
    -11, -4, 6, 2, -10, 0, -1, 9, 3,
    -- filter=8 channel=3
    1, -9, 11, 2, 7, 9, 5, 7, 17,
    -- filter=8 channel=4
    0, 1, -6, -8, 4, 4, 1, 9, 12,
    -- filter=8 channel=5
    -2, 0, -2, -5, 7, -6, 2, 9, 4,
    -- filter=8 channel=6
    2, 0, 7, -3, -1, 9, -7, 5, 12,
    -- filter=8 channel=7
    10, 1, 11, 3, 6, -1, 0, 11, 14,
    -- filter=8 channel=8
    -3, -13, 0, -8, -12, 7, 4, 12, 6,
    -- filter=8 channel=9
    4, -10, 2, -9, -11, 10, -2, 2, 11,
    -- filter=8 channel=10
    -1, -5, -7, 8, -4, -2, 3, 0, 4,
    -- filter=8 channel=11
    -5, -11, 5, -5, -1, 0, -12, -6, 5,
    -- filter=8 channel=12
    -8, 7, 8, 2, -8, 1, 4, -7, -5,
    -- filter=8 channel=13
    0, 4, 7, -2, 4, 7, -8, 6, 10,
    -- filter=8 channel=14
    1, 8, 11, 5, 1, 10, 5, 3, 8,
    -- filter=8 channel=15
    -7, -3, 4, -16, 12, 12, -4, 4, 20,
    -- filter=8 channel=16
    -15, -18, -3, -20, 5, 5, 7, 2, 10,
    -- filter=8 channel=17
    -2, 0, -7, -6, -7, 6, -6, 0, 7,
    -- filter=8 channel=18
    -11, 4, 6, -5, -3, 2, 5, 8, 6,
    -- filter=8 channel=19
    4, -3, -4, 6, -14, 2, -6, 0, -2,
    -- filter=8 channel=20
    -8, 5, 9, 10, 11, 0, 4, 5, 8,
    -- filter=8 channel=21
    4, 2, -6, -9, -10, 2, 10, -5, 1,
    -- filter=8 channel=22
    10, 8, -3, -7, -4, -7, -1, 9, 2,
    -- filter=8 channel=23
    9, -9, -11, 3, -13, -5, -5, 5, 10,
    -- filter=8 channel=24
    6, -12, -8, -7, -8, 6, -1, 6, 12,
    -- filter=8 channel=25
    -9, -17, 0, -16, 5, -2, -8, 6, 1,
    -- filter=8 channel=26
    -1, 8, -1, 5, -2, 7, -5, 13, 9,
    -- filter=8 channel=27
    -11, -6, -9, -3, -4, 14, 5, -7, 8,
    -- filter=8 channel=28
    -12, -8, 1, -14, 0, 0, -5, 11, 16,
    -- filter=8 channel=29
    -6, -6, -3, -6, 9, 26, -11, 17, 9,
    -- filter=8 channel=30
    26, 15, 9, 25, -2, 20, 12, 15, 9,
    -- filter=8 channel=31
    9, 0, -8, 7, -1, 8, -10, 2, 6,
    -- filter=8 channel=32
    -2, -4, 7, -1, 2, -8, 1, -5, -5,
    -- filter=8 channel=33
    7, -2, 8, -10, 0, -2, 8, 5, -3,
    -- filter=8 channel=34
    3, 0, 10, -3, 1, 12, 6, -2, -2,
    -- filter=8 channel=35
    -4, -5, 0, -15, 3, 9, 3, 0, -3,
    -- filter=8 channel=36
    4, 4, -3, 5, -5, -5, 8, 5, -11,
    -- filter=8 channel=37
    8, -11, -7, -7, -12, 3, -8, 5, 2,
    -- filter=8 channel=38
    3, -1, 10, -11, -10, 2, -11, 0, 11,
    -- filter=8 channel=39
    7, 2, -7, 8, -1, 4, 3, 9, 0,
    -- filter=8 channel=40
    2, 7, 9, -5, 5, 2, 6, 10, -6,
    -- filter=8 channel=41
    1, -21, 9, -4, 9, 17, 4, 11, 9,
    -- filter=8 channel=42
    -1, -3, 6, -1, 7, 0, 8, -10, -9,
    -- filter=8 channel=43
    7, 18, 11, 15, 14, 13, 12, 17, 6,
    -- filter=8 channel=44
    -1, 2, -5, 4, 3, -6, 0, 4, -4,
    -- filter=8 channel=45
    9, 7, 3, -8, -5, 1, 8, -10, -10,
    -- filter=8 channel=46
    -4, 7, 6, 13, 11, 13, 8, 0, 5,
    -- filter=8 channel=47
    -6, 0, 5, -8, 0, -3, 5, 0, 2,
    -- filter=8 channel=48
    -14, -10, 0, 5, 7, 15, 2, -5, -6,
    -- filter=8 channel=49
    -13, 3, -7, 6, 10, 4, 13, -2, 4,
    -- filter=8 channel=50
    18, 20, -2, 10, 8, 7, -1, 2, 7,
    -- filter=8 channel=51
    3, -6, -7, 9, -2, 6, -4, -9, -4,
    -- filter=8 channel=52
    3, 2, 0, 0, 7, 2, 4, 8, 3,
    -- filter=8 channel=53
    10, 1, -4, 19, 0, 13, 4, 13, 5,
    -- filter=8 channel=54
    -7, -2, 10, -6, -5, -2, -6, -2, 0,
    -- filter=8 channel=55
    0, 2, 3, 0, 0, -4, -3, 10, -4,
    -- filter=8 channel=56
    1, -1, -2, -3, 5, 6, 8, 10, 5,
    -- filter=8 channel=57
    0, -7, 3, -6, -9, 9, -2, 4, 5,
    -- filter=8 channel=58
    5, -4, -6, 7, 11, 7, -5, -1, 5,
    -- filter=8 channel=59
    0, -8, -4, 0, -9, 1, -1, 3, 5,
    -- filter=8 channel=60
    -6, -6, 0, -16, -4, 6, 0, 21, 21,
    -- filter=8 channel=61
    10, -6, 0, 2, -16, 16, -6, 0, 21,
    -- filter=8 channel=62
    -7, -9, 7, 0, -8, 2, 0, 8, -1,
    -- filter=8 channel=63
    8, -4, -6, 2, 4, -9, 8, 7, -5,
    -- filter=9 channel=0
    -1, 0, -7, 3, 9, 9, 5, 1, 10,
    -- filter=9 channel=1
    -5, 0, 0, -8, 6, -8, 4, -4, 0,
    -- filter=9 channel=2
    7, 5, 5, -3, 10, 6, 1, 3, 5,
    -- filter=9 channel=3
    12, 5, -9, 13, -6, -7, 3, -3, 5,
    -- filter=9 channel=4
    -10, 5, -10, 0, 2, -3, 9, 0, -2,
    -- filter=9 channel=5
    -7, -9, 2, 0, 2, 1, 0, 2, -15,
    -- filter=9 channel=6
    -11, 0, -3, -2, -3, 0, -10, 6, 0,
    -- filter=9 channel=7
    -11, 0, -7, 4, 5, -11, 0, -1, -6,
    -- filter=9 channel=8
    -1, 5, -2, 11, 8, 13, -2, -1, -2,
    -- filter=9 channel=9
    -4, 8, 1, 1, 1, 4, 4, -8, 0,
    -- filter=9 channel=10
    0, -7, 8, 2, 5, -6, 5, -5, 3,
    -- filter=9 channel=11
    5, -10, -2, -2, 9, 6, 1, 2, 1,
    -- filter=9 channel=12
    -8, -2, -10, 11, -2, -2, 5, 10, 9,
    -- filter=9 channel=13
    -1, -8, 5, -4, 6, 0, -6, 8, -8,
    -- filter=9 channel=14
    0, 0, -5, -6, -7, 2, 5, 0, -10,
    -- filter=9 channel=15
    6, -6, 0, 6, -5, 12, -11, -11, 4,
    -- filter=9 channel=16
    -4, -13, -13, 0, -8, -2, -1, 1, -9,
    -- filter=9 channel=17
    8, 0, 0, 8, 0, 14, -10, -2, 0,
    -- filter=9 channel=18
    1, 7, 4, 10, 8, -8, -8, -5, -8,
    -- filter=9 channel=19
    7, 4, 0, -9, -13, -8, -5, -12, -14,
    -- filter=9 channel=20
    0, -14, -5, -8, -7, -3, 0, -7, -3,
    -- filter=9 channel=21
    2, 4, -3, 4, -3, -7, -8, -5, 4,
    -- filter=9 channel=22
    -2, -6, -6, 6, -2, 10, 4, -1, 4,
    -- filter=9 channel=23
    -10, 6, 10, -3, 4, 6, -4, 3, 12,
    -- filter=9 channel=24
    -5, 7, 0, 9, 8, 10, 9, -3, 7,
    -- filter=9 channel=25
    -7, -4, 1, 7, -6, 0, 4, -3, 9,
    -- filter=9 channel=26
    -6, -14, -15, -5, -13, 2, -9, -14, -12,
    -- filter=9 channel=27
    -8, 8, -4, -1, 7, 17, -5, -6, -1,
    -- filter=9 channel=28
    5, -11, -4, 4, 8, -6, -5, -14, -3,
    -- filter=9 channel=29
    2, -4, 4, 9, 7, -8, -7, 3, -4,
    -- filter=9 channel=30
    -7, -14, -4, -19, -13, -12, -18, -23, -24,
    -- filter=9 channel=31
    3, 4, 8, 5, -5, -7, 7, -5, 3,
    -- filter=9 channel=32
    -8, 0, 11, 5, -8, 8, 7, 2, 8,
    -- filter=9 channel=33
    -6, -1, -7, -6, 1, -3, 0, -9, 9,
    -- filter=9 channel=34
    2, 1, 6, -3, -3, -4, -13, -9, 5,
    -- filter=9 channel=35
    -6, 4, 14, 3, 3, 12, 10, 15, 1,
    -- filter=9 channel=36
    0, -9, -6, 10, 8, -7, -7, 0, -4,
    -- filter=9 channel=37
    2, 1, 2, 4, -5, 5, 8, -6, 1,
    -- filter=9 channel=38
    -7, 6, 9, -5, 10, 5, -2, -1, 14,
    -- filter=9 channel=39
    5, 8, 9, 4, -1, 4, -10, 8, -5,
    -- filter=9 channel=40
    -3, -7, 8, -3, -1, -7, -5, -7, 9,
    -- filter=9 channel=41
    2, 10, -5, -6, 7, 12, -2, -5, 10,
    -- filter=9 channel=42
    -1, -5, 6, 3, 7, 7, 1, 0, 7,
    -- filter=9 channel=43
    -6, -20, -22, -3, -6, -18, 1, -6, 8,
    -- filter=9 channel=44
    -5, 7, -2, -5, -8, 8, -10, -2, 5,
    -- filter=9 channel=45
    4, 0, 8, 9, 0, -4, 4, 0, -7,
    -- filter=9 channel=46
    5, -2, -5, -11, -13, -11, -13, -2, -12,
    -- filter=9 channel=47
    3, 9, 8, -6, 5, -5, 7, -5, 1,
    -- filter=9 channel=48
    -2, -5, 4, -5, 2, -9, 6, -4, -3,
    -- filter=9 channel=49
    3, 3, -1, 7, 11, -1, -3, 5, 8,
    -- filter=9 channel=50
    -11, -3, -18, -16, -18, -8, -9, 2, -12,
    -- filter=9 channel=51
    -12, 0, 13, 9, 8, -4, -4, 6, 10,
    -- filter=9 channel=52
    -6, 8, 0, 6, -6, -6, -8, 7, -2,
    -- filter=9 channel=53
    4, 2, -5, -1, -13, -11, -1, -3, -3,
    -- filter=9 channel=54
    12, 8, 7, 9, 6, -10, -1, -3, -7,
    -- filter=9 channel=55
    8, 4, 7, 3, -10, -9, 10, 8, -8,
    -- filter=9 channel=56
    5, -10, -7, 2, 4, -10, 0, -4, 4,
    -- filter=9 channel=57
    -9, 10, 0, 7, -4, 8, -7, 0, -2,
    -- filter=9 channel=58
    -8, 4, -9, -5, -4, -9, 9, 5, 8,
    -- filter=9 channel=59
    7, -6, -8, 9, 4, 11, -7, -2, 9,
    -- filter=9 channel=60
    -5, -9, 5, 8, 2, 17, 6, 5, 2,
    -- filter=9 channel=61
    -1, 1, 6, 10, 5, 15, 1, 7, 5,
    -- filter=9 channel=62
    -5, 7, -1, 7, 12, 1, 7, -4, -7,
    -- filter=9 channel=63
    -4, 1, -1, 9, 2, 6, 0, 0, 4,
    -- filter=10 channel=0
    8, 11, 0, 4, 19, 8, 3, 8, -7,
    -- filter=10 channel=1
    -22, -11, 0, -12, -15, -2, -5, -13, -20,
    -- filter=10 channel=2
    -18, -6, 0, -19, -25, -8, -21, -23, -8,
    -- filter=10 channel=3
    -4, 0, 14, 5, 12, 11, 4, -3, 0,
    -- filter=10 channel=4
    2, 14, 2, 11, 12, 14, 4, 0, -2,
    -- filter=10 channel=5
    9, 8, 2, 8, 6, -5, -6, -5, -9,
    -- filter=10 channel=6
    2, -4, -3, 0, 0, 0, -11, -15, -11,
    -- filter=10 channel=7
    4, -3, 11, 3, 12, 9, -4, 9, 5,
    -- filter=10 channel=8
    24, 24, 14, 9, 17, 11, 4, -9, 1,
    -- filter=10 channel=9
    0, -3, 0, 3, 11, 3, 4, -9, 3,
    -- filter=10 channel=10
    -6, 0, 7, -3, 3, -7, 6, 9, 8,
    -- filter=10 channel=11
    2, -1, -4, -2, -3, -2, -1, 7, 0,
    -- filter=10 channel=12
    -7, 1, -3, -2, -4, -3, -2, 9, -8,
    -- filter=10 channel=13
    10, 11, -4, 17, 3, 0, 7, 11, -4,
    -- filter=10 channel=14
    9, 1, 3, 3, 12, 4, 7, 9, 2,
    -- filter=10 channel=15
    6, 20, 7, 3, 9, -5, -9, 4, -1,
    -- filter=10 channel=16
    3, 0, 0, 2, -8, -12, 0, -15, -13,
    -- filter=10 channel=17
    14, 13, 10, 9, 20, 2, 9, -2, 4,
    -- filter=10 channel=18
    10, 13, -7, 4, 11, 11, 12, 16, 8,
    -- filter=10 channel=19
    -9, -13, -4, -8, -1, -12, 0, -3, 0,
    -- filter=10 channel=20
    -3, -7, 1, -4, 6, 0, 10, -9, 10,
    -- filter=10 channel=21
    8, -5, -6, 1, -5, -3, 6, 5, -8,
    -- filter=10 channel=22
    9, 1, 8, 0, -6, 0, -1, 0, 0,
    -- filter=10 channel=23
    3, 8, -4, 4, -1, -1, 8, 9, 0,
    -- filter=10 channel=24
    5, 6, 0, 0, 20, 10, 12, 7, 1,
    -- filter=10 channel=25
    -13, -22, -17, -13, -11, -19, -23, -17, -8,
    -- filter=10 channel=26
    -7, 0, 7, 8, -6, -1, 1, -7, -8,
    -- filter=10 channel=27
    7, 0, -6, -5, -9, 3, 0, -3, -9,
    -- filter=10 channel=28
    -2, 13, 3, 3, -3, -2, -12, -3, -6,
    -- filter=10 channel=29
    7, 13, 3, 7, 6, -7, -7, -21, -23,
    -- filter=10 channel=30
    7, 12, -1, -4, 15, 2, 9, -3, 5,
    -- filter=10 channel=31
    5, 10, 8, -1, -2, -9, 7, 5, 1,
    -- filter=10 channel=32
    -11, -8, -8, -2, -10, -13, -16, -12, -4,
    -- filter=10 channel=33
    7, -9, 10, 7, 6, 2, 4, 2, -6,
    -- filter=10 channel=34
    2, 2, -5, -2, 0, 1, -6, -4, 1,
    -- filter=10 channel=35
    0, -2, -3, -7, -17, -1, -11, -11, -11,
    -- filter=10 channel=36
    -4, -2, 9, 0, 1, -6, -6, 4, -1,
    -- filter=10 channel=37
    11, -4, -4, 5, 1, -4, 6, 4, -9,
    -- filter=10 channel=38
    6, 10, 13, -1, 11, 9, -6, -17, -13,
    -- filter=10 channel=39
    7, -9, 2, 0, 7, -3, 7, 6, 3,
    -- filter=10 channel=40
    4, 5, -8, -1, -1, 2, 2, -12, -1,
    -- filter=10 channel=41
    15, 5, 0, 0, 0, -5, -3, -15, -10,
    -- filter=10 channel=42
    -10, -1, -1, 10, 7, -10, 1, 0, 6,
    -- filter=10 channel=43
    -17, -8, -10, -1, -4, -13, -19, -3, -14,
    -- filter=10 channel=44
    -12, -3, 0, -11, -5, -6, -8, 2, -1,
    -- filter=10 channel=45
    -6, 7, -8, 9, -7, 9, -5, 0, 9,
    -- filter=10 channel=46
    10, 12, 8, 6, 4, 11, 0, 8, 0,
    -- filter=10 channel=47
    2, -6, -9, -7, 9, 8, 3, -7, 5,
    -- filter=10 channel=48
    -2, 6, 8, 11, -8, -9, 0, 0, -14,
    -- filter=10 channel=49
    10, 1, -2, -2, -2, -4, 1, 11, -9,
    -- filter=10 channel=50
    7, -3, -3, 8, -5, 11, 4, -6, -3,
    -- filter=10 channel=51
    1, 0, -1, 17, 4, 0, 12, 10, 1,
    -- filter=10 channel=52
    4, -5, 8, -2, -2, -6, -7, -5, 0,
    -- filter=10 channel=53
    -12, -4, 0, 0, -2, 2, -6, 0, -4,
    -- filter=10 channel=54
    -4, -2, -6, 11, 6, -9, 10, 2, -6,
    -- filter=10 channel=55
    -10, 6, -8, -5, 9, 3, 4, -9, 0,
    -- filter=10 channel=56
    -6, 5, 11, -3, -2, -7, -2, 7, 3,
    -- filter=10 channel=57
    8, 10, 0, 1, -4, 4, -3, 6, -9,
    -- filter=10 channel=58
    -7, -9, -5, 6, 2, -4, 7, 4, -2,
    -- filter=10 channel=59
    6, 15, 15, 4, -9, -4, -13, -20, 3,
    -- filter=10 channel=60
    26, 33, 17, 22, 19, 2, 0, 9, 5,
    -- filter=10 channel=61
    19, 14, 21, 17, 24, 7, -5, 12, 6,
    -- filter=10 channel=62
    -5, 15, 13, -5, 4, -8, 3, -8, 3,
    -- filter=10 channel=63
    -10, -2, 0, -1, 3, 6, 1, 0, -6,
    -- filter=11 channel=0
    0, -2, 1, -5, 1, -6, -7, -9, 9,
    -- filter=11 channel=1
    -4, 3, -12, 6, -3, -7, 2, -6, 3,
    -- filter=11 channel=2
    -13, -1, 1, -1, -1, -2, -3, -5, -4,
    -- filter=11 channel=3
    -9, 0, 10, 7, -7, 0, 9, 2, 3,
    -- filter=11 channel=4
    -2, 11, 0, 0, 9, 4, 1, 6, -2,
    -- filter=11 channel=5
    7, -2, 9, -7, -7, -3, -5, 4, -10,
    -- filter=11 channel=6
    6, -3, 4, 4, 10, 0, 1, -5, -3,
    -- filter=11 channel=7
    -4, -4, -2, 4, 3, -4, -1, 6, 0,
    -- filter=11 channel=8
    8, -8, 7, -1, 4, 12, 7, -10, -8,
    -- filter=11 channel=9
    3, 36, 35, 22, 45, 41, 17, 37, 49,
    -- filter=11 channel=10
    -6, -2, 0, 7, -8, -14, 10, -8, 0,
    -- filter=11 channel=11
    3, 4, -10, 4, -8, 5, -4, 0, -9,
    -- filter=11 channel=12
    -6, 0, 3, 6, -4, -6, 3, 5, -7,
    -- filter=11 channel=13
    9, -3, 1, 9, 0, 1, 8, -3, 7,
    -- filter=11 channel=14
    0, 3, -8, 0, -10, -11, -8, -3, 1,
    -- filter=11 channel=15
    1, -7, 2, 5, 13, 13, -8, 4, 10,
    -- filter=11 channel=16
    -10, 4, -9, 4, -2, -5, -6, 7, 5,
    -- filter=11 channel=17
    3, -2, -7, -5, 10, 2, 3, 0, -10,
    -- filter=11 channel=18
    1, 4, 22, 13, 4, 10, 11, 12, 13,
    -- filter=11 channel=19
    0, 9, 7, 1, 10, -4, 1, 9, -2,
    -- filter=11 channel=20
    -1, -3, 16, 11, 13, 9, 13, 17, 7,
    -- filter=11 channel=21
    -7, -1, 12, -1, 11, 4, -7, -7, 14,
    -- filter=11 channel=22
    -7, -10, 1, -9, 5, -2, 0, -1, 10,
    -- filter=11 channel=23
    -5, 3, -3, -8, -11, -13, 8, 0, 2,
    -- filter=11 channel=24
    -8, 2, 3, 2, 7, -4, 0, 5, 3,
    -- filter=11 channel=25
    -1, -18, -6, -10, -16, -9, 5, -3, -15,
    -- filter=11 channel=26
    -14, -14, 5, -1, -13, -13, -6, 3, -11,
    -- filter=11 channel=27
    1, -4, -4, -8, -17, -10, 3, -10, -18,
    -- filter=11 channel=28
    11, 12, 11, 0, 12, 2, -7, 11, 0,
    -- filter=11 channel=29
    4, 5, 2, 6, -1, 18, 5, 7, 4,
    -- filter=11 channel=30
    -5, -21, -16, -22, -19, -4, -9, -9, -6,
    -- filter=11 channel=31
    9, -6, 1, -8, 10, 5, 4, -1, 7,
    -- filter=11 channel=32
    3, -1, -5, -6, -8, -9, -3, -13, -5,
    -- filter=11 channel=33
    1, 7, 3, 4, 8, -9, 0, 8, -10,
    -- filter=11 channel=34
    3, -11, 4, 3, -12, -2, -3, -2, -3,
    -- filter=11 channel=35
    -9, -5, -13, -14, -14, -20, -13, -19, -4,
    -- filter=11 channel=36
    8, 1, -6, 6, -4, -1, -2, -8, 9,
    -- filter=11 channel=37
    -2, 7, 6, 10, 5, 3, 5, -4, 11,
    -- filter=11 channel=38
    -6, -8, -12, -11, -11, 3, -4, -4, 5,
    -- filter=11 channel=39
    -5, -5, 10, 0, 5, 7, -4, 0, -4,
    -- filter=11 channel=40
    -6, 8, -11, -11, -3, -3, -9, -3, 6,
    -- filter=11 channel=41
    -10, 1, 1, 7, 7, -1, -12, -4, -1,
    -- filter=11 channel=42
    5, 8, -8, 5, -4, 7, 2, -7, -9,
    -- filter=11 channel=43
    -6, -5, -10, -19, -16, 0, -10, -3, -8,
    -- filter=11 channel=44
    0, -14, -13, -15, 0, 2, -8, -5, -13,
    -- filter=11 channel=45
    0, 0, -10, 4, 5, 4, -9, 8, -9,
    -- filter=11 channel=46
    -4, -5, -6, -3, -8, 6, -2, 0, -11,
    -- filter=11 channel=47
    2, -5, -2, -7, 0, -7, 4, 0, -5,
    -- filter=11 channel=48
    0, 0, -6, -8, 12, 15, 0, 7, 9,
    -- filter=11 channel=49
    12, -4, -7, 7, -1, -7, -7, -6, 6,
    -- filter=11 channel=50
    -6, -14, -2, -4, -10, 4, -4, -1, 7,
    -- filter=11 channel=51
    9, 10, 5, 4, -6, -7, 1, 9, -2,
    -- filter=11 channel=52
    10, 10, 2, 9, 3, -5, -2, -3, 1,
    -- filter=11 channel=53
    -7, -12, -17, -1, -8, -7, -2, -20, -7,
    -- filter=11 channel=54
    16, 13, 18, 7, 20, 26, 20, 15, 24,
    -- filter=11 channel=55
    4, 5, 3, -10, 8, 9, 6, 6, -10,
    -- filter=11 channel=56
    4, -8, 0, 2, -6, -6, 1, 3, -7,
    -- filter=11 channel=57
    -7, -1, 0, -1, -9, -9, -5, -4, -7,
    -- filter=11 channel=58
    -2, 0, 5, 9, -1, 7, 17, 12, 14,
    -- filter=11 channel=59
    -2, -4, -1, 3, -9, 2, 5, -8, -4,
    -- filter=11 channel=60
    9, -13, 0, 3, 4, 9, 6, -9, 7,
    -- filter=11 channel=61
    4, -11, 0, -2, -11, 5, 7, 2, -5,
    -- filter=11 channel=62
    -1, 0, -8, -6, 0, -9, -3, -8, 7,
    -- filter=11 channel=63
    4, 4, 0, 0, -10, 1, 3, -2, -7,
    -- filter=12 channel=0
    1, 3, -17, 13, 2, -10, 1, -2, -16,
    -- filter=12 channel=1
    -13, 7, 8, -7, 4, 0, -15, 2, 3,
    -- filter=12 channel=2
    -8, 3, -5, -13, 20, -4, 1, 11, -11,
    -- filter=12 channel=3
    -7, 9, -13, 8, 17, -12, -6, 6, -11,
    -- filter=12 channel=4
    -2, 1, -1, -6, 6, -7, 0, 5, -6,
    -- filter=12 channel=5
    -11, 0, 4, -3, -5, 6, -10, 3, 16,
    -- filter=12 channel=6
    -2, 11, 0, -2, -2, -3, 5, -6, -9,
    -- filter=12 channel=7
    -3, -6, 16, 9, 2, 6, -5, 2, 7,
    -- filter=12 channel=8
    -10, 16, 0, -3, 13, -5, -4, 10, -16,
    -- filter=12 channel=9
    -11, 0, 5, -3, 2, -7, -3, 9, 0,
    -- filter=12 channel=10
    11, -10, 0, -1, 0, 0, 8, 7, -5,
    -- filter=12 channel=11
    -16, 8, -5, -18, 5, -12, -4, 0, -6,
    -- filter=12 channel=12
    5, -10, -9, 7, -4, 2, 2, -7, 4,
    -- filter=12 channel=13
    -7, 10, -2, 1, 12, -6, -6, 9, -9,
    -- filter=12 channel=14
    0, -3, 7, 3, 2, 18, 12, -2, 8,
    -- filter=12 channel=15
    -11, 22, -4, 6, 22, -19, 1, 21, 0,
    -- filter=12 channel=16
    -18, 9, -6, -14, 23, -9, -9, 12, -17,
    -- filter=12 channel=17
    -3, 0, 9, -9, 23, -2, -11, 2, -5,
    -- filter=12 channel=18
    -3, -2, 3, 5, 8, -2, 3, 7, -13,
    -- filter=12 channel=19
    -6, -6, 13, -19, 4, 13, -10, -6, 8,
    -- filter=12 channel=20
    -1, 8, 10, 13, 7, -4, 10, 0, -4,
    -- filter=12 channel=21
    -10, 7, -10, -10, 3, -4, 7, -10, 8,
    -- filter=12 channel=22
    0, 6, -3, -8, 3, -1, -8, -2, 7,
    -- filter=12 channel=23
    -1, 0, 1, -4, 13, -12, 0, -1, -11,
    -- filter=12 channel=24
    -9, 8, 8, -3, 12, 0, -5, 8, 0,
    -- filter=12 channel=25
    -4, 10, -6, -12, 15, -11, -12, 0, 0,
    -- filter=12 channel=26
    4, 2, -3, 21, 9, -4, 11, 13, 6,
    -- filter=12 channel=27
    -12, 2, -4, 4, 13, -11, 7, 11, 1,
    -- filter=12 channel=28
    -6, 15, 3, -9, 18, -3, -5, 5, -7,
    -- filter=12 channel=29
    -15, 21, -6, -3, 33, -18, 5, 21, -8,
    -- filter=12 channel=30
    11, 22, 28, 4, 12, 23, 5, 12, 21,
    -- filter=12 channel=31
    0, -6, 1, 7, 7, -8, 9, 6, -10,
    -- filter=12 channel=32
    -2, -1, 2, -8, 10, 14, 1, 7, -7,
    -- filter=12 channel=33
    -8, -4, 0, 5, 7, 9, -9, 9, 4,
    -- filter=12 channel=34
    6, 3, 3, 9, 0, 10, 7, 0, 10,
    -- filter=12 channel=35
    -7, 16, -19, 9, 10, -23, 4, 10, -14,
    -- filter=12 channel=36
    0, -6, -9, 5, -1, 9, 0, -3, 4,
    -- filter=12 channel=37
    -4, -2, 3, -15, 14, 3, -5, 15, -4,
    -- filter=12 channel=38
    -12, 19, 2, -8, 13, -16, -10, 12, -18,
    -- filter=12 channel=39
    -8, 1, -6, 8, -7, -7, 7, -6, 9,
    -- filter=12 channel=40
    -1, 10, -4, -7, -7, -7, 2, 4, 6,
    -- filter=12 channel=41
    -2, 15, -3, 4, 23, -27, -8, 15, -6,
    -- filter=12 channel=42
    1, -8, -6, 6, 4, -3, -4, 1, 5,
    -- filter=12 channel=43
    3, -4, 12, -8, 8, 3, -1, 6, 2,
    -- filter=12 channel=44
    6, -4, 0, 4, 0, 11, 0, -7, 4,
    -- filter=12 channel=45
    8, -7, 1, -5, -8, -3, -9, -1, -1,
    -- filter=12 channel=46
    5, 20, 10, 16, 3, 1, 11, 13, 12,
    -- filter=12 channel=47
    -5, 0, -9, 9, 7, 9, -4, -7, -5,
    -- filter=12 channel=48
    -8, 8, 5, 12, 4, 1, -7, 5, -2,
    -- filter=12 channel=49
    -5, 9, -4, -2, 5, -13, 8, -4, 6,
    -- filter=12 channel=50
    4, -2, 25, 1, 1, 31, 13, 4, 18,
    -- filter=12 channel=51
    9, 8, 4, 15, -5, -3, 10, -3, -10,
    -- filter=12 channel=52
    6, -1, -1, -7, -3, -9, 10, -8, 2,
    -- filter=12 channel=53
    15, 0, 14, 8, 12, 18, 7, 8, 25,
    -- filter=12 channel=54
    -9, 2, -4, -1, 8, 2, 1, -1, -8,
    -- filter=12 channel=55
    0, -1, -7, -7, 3, 7, -9, -9, 4,
    -- filter=12 channel=56
    -5, 4, 0, 8, 0, 12, 0, -3, 13,
    -- filter=12 channel=57
    -10, 6, 8, 3, -9, 8, -9, 9, 1,
    -- filter=12 channel=58
    -4, -1, -6, -5, -3, 0, 8, -11, 7,
    -- filter=12 channel=59
    -16, 19, 1, -6, 21, -19, 8, 13, -11,
    -- filter=12 channel=60
    -6, 31, -18, -10, 38, -34, -1, 21, -16,
    -- filter=12 channel=61
    -18, -1, 0, -2, 26, -8, -5, 5, -14,
    -- filter=12 channel=62
    -7, 10, -2, -13, -1, -11, -2, 5, -2,
    -- filter=12 channel=63
    6, 10, -5, 2, 5, 1, 1, 7, -9,
    -- filter=13 channel=0
    1, -5, -14, 10, 0, -14, 2, -7, 1,
    -- filter=13 channel=1
    -10, 7, -11, -11, 13, -2, -8, -1, 6,
    -- filter=13 channel=2
    5, 0, -9, 9, 8, -8, -19, -6, -8,
    -- filter=13 channel=3
    2, 5, -4, 9, 16, 8, -9, 0, -11,
    -- filter=13 channel=4
    0, -3, 0, -2, 4, 7, 7, 1, -7,
    -- filter=13 channel=5
    4, 14, 1, -3, 7, 5, -4, 13, 11,
    -- filter=13 channel=6
    2, 0, 0, 9, 8, 5, 6, -6, -2,
    -- filter=13 channel=7
    -3, 6, 0, -6, 16, 4, 3, 15, 0,
    -- filter=13 channel=8
    2, 12, 2, 20, 17, 9, -10, 10, -8,
    -- filter=13 channel=9
    -6, 0, -4, 9, 18, -2, 3, 1, -2,
    -- filter=13 channel=10
    2, 1, -3, 5, 0, 5, 2, -7, 3,
    -- filter=13 channel=11
    -14, 8, -10, 7, 5, 10, -8, 8, -11,
    -- filter=13 channel=12
    -3, -3, -5, 3, 0, 8, 4, -5, -9,
    -- filter=13 channel=13
    0, 8, -1, 17, 4, 3, 3, 2, -11,
    -- filter=13 channel=14
    0, 1, 9, 9, 10, 1, -1, 16, 6,
    -- filter=13 channel=15
    8, 3, -1, 9, 22, -8, 1, 11, -2,
    -- filter=13 channel=16
    0, 0, -3, 20, 14, -6, 1, -2, -2,
    -- filter=13 channel=17
    -1, 5, -5, 13, 16, 14, -11, -4, -8,
    -- filter=13 channel=18
    2, 3, 6, 16, 0, 2, 13, 0, -11,
    -- filter=13 channel=19
    6, -2, 0, -11, 10, 9, -8, 1, -2,
    -- filter=13 channel=20
    -3, 8, 10, 16, 1, 5, 12, 15, 7,
    -- filter=13 channel=21
    -7, 0, 10, 4, -8, 2, 0, 2, -9,
    -- filter=13 channel=22
    -1, 3, 10, 9, 9, -1, 5, -4, 3,
    -- filter=13 channel=23
    -7, 3, -7, -16, 2, 1, 0, -12, -2,
    -- filter=13 channel=24
    8, 7, 0, 6, 2, 6, -3, 0, 2,
    -- filter=13 channel=25
    -3, 7, -12, -1, 12, -6, -1, -10, -3,
    -- filter=13 channel=26
    -4, 9, 5, 10, 15, -2, -1, 3, 4,
    -- filter=13 channel=27
    6, 0, -10, -9, 12, -2, -18, -3, -9,
    -- filter=13 channel=28
    -7, 3, -13, 14, 27, 8, 0, 9, -1,
    -- filter=13 channel=29
    12, 0, -15, 26, 28, -9, -7, 0, -5,
    -- filter=13 channel=30
    7, 34, 28, 16, 25, 27, 0, 21, 22,
    -- filter=13 channel=31
    -6, 8, 1, 3, -7, -1, -2, -8, -1,
    -- filter=13 channel=32
    -5, -3, -5, -7, -3, -5, -6, -9, 1,
    -- filter=13 channel=33
    -3, -3, -10, -5, 1, -4, 0, -4, 9,
    -- filter=13 channel=34
    1, 10, 7, -4, 2, -3, -3, -1, 5,
    -- filter=13 channel=35
    -7, -6, 4, -4, 3, -13, -1, -1, -14,
    -- filter=13 channel=36
    2, 3, -8, 3, 7, -8, -7, 8, 0,
    -- filter=13 channel=37
    7, -2, -10, 7, 2, 8, -8, 8, -11,
    -- filter=13 channel=38
    6, 4, -15, 0, 3, -15, -5, 3, -13,
    -- filter=13 channel=39
    10, 1, 6, -2, 3, -7, 2, 8, 2,
    -- filter=13 channel=40
    -4, 6, -3, 9, 9, 1, -3, -11, -6,
    -- filter=13 channel=41
    7, 1, -1, 11, 23, -5, -2, -10, -7,
    -- filter=13 channel=42
    -3, -5, -8, 6, -2, 1, -3, 10, 4,
    -- filter=13 channel=43
    -6, 4, -5, 13, 4, 11, 14, 18, 16,
    -- filter=13 channel=44
    -9, 11, 4, 1, 4, 0, -11, 10, 14,
    -- filter=13 channel=45
    -4, 10, 10, 10, -4, -7, 0, 7, 4,
    -- filter=13 channel=46
    5, 19, 10, 4, 12, 7, 15, 8, 13,
    -- filter=13 channel=47
    -3, -7, 3, 2, -2, -8, 3, 7, -1,
    -- filter=13 channel=48
    9, 13, -5, 2, 2, 7, 7, 9, 2,
    -- filter=13 channel=49
    -5, 12, -6, 11, 6, 4, -8, -12, -15,
    -- filter=13 channel=50
    4, 12, 16, -2, 18, 19, 14, 21, 17,
    -- filter=13 channel=51
    -1, 6, -6, 0, -11, -10, 9, -10, -6,
    -- filter=13 channel=52
    -9, -5, -2, 0, 1, 8, 8, -9, -5,
    -- filter=13 channel=53
    0, 17, 9, -1, 16, 21, 6, 23, 7,
    -- filter=13 channel=54
    -5, 14, -6, 5, 12, 3, -11, -1, -3,
    -- filter=13 channel=55
    -2, 0, 8, 5, -2, -4, -5, -8, -3,
    -- filter=13 channel=56
    0, 3, 7, 1, 5, 8, 12, 8, 8,
    -- filter=13 channel=57
    7, -1, 0, -9, -4, -5, -7, -4, 5,
    -- filter=13 channel=58
    0, 3, 4, -2, -8, -10, 0, -6, -8,
    -- filter=13 channel=59
    6, 12, -15, 1, 0, -10, -7, -11, -1,
    -- filter=13 channel=60
    10, 15, -14, 10, 19, 1, 5, 9, -8,
    -- filter=13 channel=61
    1, 0, -8, 8, 22, 0, -3, -5, -9,
    -- filter=13 channel=62
    5, 6, -11, -1, 15, 4, 4, 8, -13,
    -- filter=13 channel=63
    3, 6, 0, 3, 6, 5, -2, 3, -1,
    -- filter=14 channel=0
    7, 5, -3, -6, 0, 8, 3, -1, -10,
    -- filter=14 channel=1
    -8, -7, -7, -7, 2, 5, 1, 2, -4,
    -- filter=14 channel=2
    6, -7, -5, 5, 8, 3, 0, 7, -8,
    -- filter=14 channel=3
    -6, 3, 7, 5, 5, 7, -7, -5, 0,
    -- filter=14 channel=4
    6, -9, -4, 6, -4, 8, 0, 0, -8,
    -- filter=14 channel=5
    -2, 4, -4, -3, -9, 6, -8, 0, -4,
    -- filter=14 channel=6
    6, 5, -5, 6, -6, 0, -4, -6, 8,
    -- filter=14 channel=7
    -9, 6, 0, -2, 5, 9, -8, 2, 5,
    -- filter=14 channel=8
    6, 4, -5, 7, 7, -7, 2, -3, 1,
    -- filter=14 channel=9
    6, -4, 3, 1, -6, -9, 8, 1, -9,
    -- filter=14 channel=10
    -5, 7, 0, 2, 3, -6, -1, -6, 10,
    -- filter=14 channel=11
    -8, 9, 3, 4, -4, -8, -6, 4, -7,
    -- filter=14 channel=12
    0, -2, 0, -8, 2, 3, 1, 4, 4,
    -- filter=14 channel=13
    -8, 2, 3, 1, -3, -7, -2, 8, -9,
    -- filter=14 channel=14
    -2, -1, 10, -6, 7, 1, -1, 7, 1,
    -- filter=14 channel=15
    -7, 8, 10, -6, -8, -2, 5, 3, 0,
    -- filter=14 channel=16
    -5, 6, -1, 0, -7, 5, -3, 4, -9,
    -- filter=14 channel=17
    -2, 2, -9, 0, -9, 1, 5, -10, -8,
    -- filter=14 channel=18
    0, 0, -3, 5, 8, -1, 6, -2, 1,
    -- filter=14 channel=19
    -9, -1, 2, 7, -1, 0, -9, -9, 9,
    -- filter=14 channel=20
    6, 10, -4, 3, 4, -3, 4, 0, 0,
    -- filter=14 channel=21
    5, -3, -1, 0, 9, -8, -2, -9, -5,
    -- filter=14 channel=22
    5, -5, 8, -1, 5, -5, 9, 0, -9,
    -- filter=14 channel=23
    0, -3, 4, -3, 1, 5, -4, -5, -4,
    -- filter=14 channel=24
    3, 8, 1, 8, 4, 6, 1, -3, -9,
    -- filter=14 channel=25
    0, -8, 7, -6, 0, 1, -6, -6, 3,
    -- filter=14 channel=26
    9, -5, -7, -9, 5, 0, -9, -1, 0,
    -- filter=14 channel=27
    -8, -7, 0, -8, 7, 2, 5, -7, 4,
    -- filter=14 channel=28
    -8, -9, 3, -4, 2, 4, 2, 8, -8,
    -- filter=14 channel=29
    9, -10, -1, -10, -6, -6, 1, -4, -2,
    -- filter=14 channel=30
    0, 8, 0, -8, -10, 0, 8, 1, 0,
    -- filter=14 channel=31
    4, 8, 0, -9, -10, 5, -2, 4, 0,
    -- filter=14 channel=32
    0, -1, 5, -5, 10, -3, -2, -6, -7,
    -- filter=14 channel=33
    -1, 2, 2, -3, -1, 5, -5, -8, -6,
    -- filter=14 channel=34
    10, -7, 3, 1, -8, 0, 0, 3, 6,
    -- filter=14 channel=35
    -6, 1, 4, 1, 4, 0, 10, -9, -1,
    -- filter=14 channel=36
    -5, -8, 0, -7, -6, 1, -9, 7, 3,
    -- filter=14 channel=37
    -1, 9, -4, -5, -3, -4, 9, 5, 8,
    -- filter=14 channel=38
    -4, -3, 9, 0, 6, -4, -1, -6, -7,
    -- filter=14 channel=39
    7, -1, -3, 10, -2, 3, 0, 0, -3,
    -- filter=14 channel=40
    10, 6, 3, 4, -3, -10, 6, -5, 7,
    -- filter=14 channel=41
    0, -7, -9, 4, 6, -6, -7, -2, 8,
    -- filter=14 channel=42
    1, -5, -8, 7, 1, 7, -7, -2, -4,
    -- filter=14 channel=43
    -8, 0, 4, 7, -1, 4, -5, 5, -5,
    -- filter=14 channel=44
    -4, 8, -7, 8, 9, 0, 9, 5, -6,
    -- filter=14 channel=45
    0, 7, 0, -5, -7, 7, -7, -5, 3,
    -- filter=14 channel=46
    -5, -8, 0, 0, -10, 0, 2, -6, -6,
    -- filter=14 channel=47
    -7, -6, -4, -1, 0, 8, 6, -5, -8,
    -- filter=14 channel=48
    -4, 0, -6, 8, -4, 8, 0, 9, -9,
    -- filter=14 channel=49
    5, 2, 8, 8, 0, 0, 8, -5, -3,
    -- filter=14 channel=50
    3, -6, -2, 9, -3, -4, -6, -6, -4,
    -- filter=14 channel=51
    4, 0, -3, 6, -6, -5, -10, 9, -8,
    -- filter=14 channel=52
    -4, 9, 10, 9, -4, 10, 9, 5, 7,
    -- filter=14 channel=53
    -2, 6, -4, 0, -2, 6, 0, -4, 0,
    -- filter=14 channel=54
    9, -9, -2, 6, 3, 10, 3, -1, 8,
    -- filter=14 channel=55
    -10, 5, 3, -8, 0, 2, -10, 7, -4,
    -- filter=14 channel=56
    4, -8, 6, -9, -1, -3, -3, -5, -2,
    -- filter=14 channel=57
    -1, 6, 1, 2, -8, 0, -6, -7, 0,
    -- filter=14 channel=58
    1, -5, -3, -6, 9, -6, 3, -4, -9,
    -- filter=14 channel=59
    -8, 4, 3, -2, 8, -2, 0, 4, -1,
    -- filter=14 channel=60
    3, -1, 6, -7, 1, -3, 6, -2, 0,
    -- filter=14 channel=61
    -2, -5, -7, -3, -5, 7, -2, 10, -7,
    -- filter=14 channel=62
    1, 4, -10, -6, 9, -1, 3, -3, -6,
    -- filter=14 channel=63
    4, -7, 0, 2, -9, -1, -9, 3, 10,
    -- filter=15 channel=0
    -10, -6, 1, 0, -1, -13, -14, -13, 0,
    -- filter=15 channel=1
    -7, 11, 12, 13, 10, 16, 10, 13, 2,
    -- filter=15 channel=2
    9, 2, 2, 0, 5, 15, 5, -1, 0,
    -- filter=15 channel=3
    9, 8, 18, 5, 9, 16, 3, 5, 14,
    -- filter=15 channel=4
    -10, -9, 0, 6, -3, 1, 1, -3, -3,
    -- filter=15 channel=5
    3, 12, 1, 16, 17, 5, 10, 4, -5,
    -- filter=15 channel=6
    3, 9, -2, 9, 9, 5, 2, 1, -8,
    -- filter=15 channel=7
    8, -9, 0, 12, 6, 4, 5, -4, -8,
    -- filter=15 channel=8
    4, 8, 0, 0, -5, -8, -1, -21, 2,
    -- filter=15 channel=9
    16, 26, 31, 27, 30, 34, 18, 37, 16,
    -- filter=15 channel=10
    3, -8, -11, 2, 1, 0, -11, -9, 0,
    -- filter=15 channel=11
    -8, 0, 2, -7, 0, 8, -9, 4, 4,
    -- filter=15 channel=12
    -4, 1, 10, 10, -3, -5, -7, 11, -1,
    -- filter=15 channel=13
    -7, 0, -9, 14, 6, -2, 0, 4, -4,
    -- filter=15 channel=14
    6, 10, -5, 3, 1, 9, 3, 3, 7,
    -- filter=15 channel=15
    14, 9, 4, -5, -4, 1, -4, -7, -8,
    -- filter=15 channel=16
    9, 5, 16, 4, 4, 20, -4, -7, 12,
    -- filter=15 channel=17
    -5, -7, 5, -6, -8, 4, 2, 2, 4,
    -- filter=15 channel=18
    8, -7, 0, 5, -6, -5, -10, 4, -2,
    -- filter=15 channel=19
    6, 25, 4, 18, 16, 19, 14, 19, 0,
    -- filter=15 channel=20
    -3, 16, 6, 7, 16, 4, 5, 8, 4,
    -- filter=15 channel=21
    -8, -7, 0, -8, 4, 8, 11, 4, -7,
    -- filter=15 channel=22
    2, -6, -6, -7, 2, 0, 10, -8, -1,
    -- filter=15 channel=23
    -16, -16, -8, -17, -16, 4, 0, -13, -3,
    -- filter=15 channel=24
    4, 3, 3, -10, -11, 0, 3, 1, 2,
    -- filter=15 channel=25
    4, 13, 5, -2, 10, 21, -2, 20, 7,
    -- filter=15 channel=26
    12, 3, -3, 12, 7, 4, 0, 3, 13,
    -- filter=15 channel=27
    -9, -6, 0, -12, -9, 11, -10, -10, 4,
    -- filter=15 channel=28
    7, 16, 2, -1, 8, 5, -6, -5, 12,
    -- filter=15 channel=29
    10, 14, 10, 20, 15, 5, -9, 1, 3,
    -- filter=15 channel=30
    -4, 2, 6, 0, -3, -4, -5, 0, -5,
    -- filter=15 channel=31
    -4, 7, 3, -4, -2, -12, 0, -7, 5,
    -- filter=15 channel=32
    -1, 7, 12, -10, -6, 11, 6, -1, 3,
    -- filter=15 channel=33
    -3, 3, -9, -4, -3, 4, -9, -2, 6,
    -- filter=15 channel=34
    3, 7, 0, -7, -7, 1, -8, -4, -6,
    -- filter=15 channel=35
    -5, -2, 1, -13, 0, -1, -4, 0, -9,
    -- filter=15 channel=36
    9, 8, -8, 0, -10, -8, 2, -10, -3,
    -- filter=15 channel=37
    14, 2, 13, 5, 19, 1, 14, 1, 13,
    -- filter=15 channel=38
    2, -4, -3, 4, -9, -4, -13, -2, 3,
    -- filter=15 channel=39
    -8, 0, -8, 10, 3, 4, -4, 5, 0,
    -- filter=15 channel=40
    0, -9, 3, 4, 2, 9, -9, 5, -4,
    -- filter=15 channel=41
    14, 11, 4, 3, 6, -7, -13, 1, 2,
    -- filter=15 channel=42
    -1, 7, 4, -6, 1, 3, 2, 8, 7,
    -- filter=15 channel=43
    4, -1, -8, 20, 1, -2, 13, 11, 0,
    -- filter=15 channel=44
    1, 16, -1, -6, 5, 9, 9, 15, 15,
    -- filter=15 channel=45
    8, 2, -1, 2, 8, -7, 2, -6, 4,
    -- filter=15 channel=46
    -3, 6, 6, -6, -3, -8, 2, 14, -3,
    -- filter=15 channel=47
    6, -8, 6, 6, 8, 0, -6, -4, 9,
    -- filter=15 channel=48
    0, 0, -4, 9, 20, -3, 8, 7, 11,
    -- filter=15 channel=49
    6, -13, 4, -1, -13, -13, -1, -9, 0,
    -- filter=15 channel=50
    0, -5, 10, 7, 15, -4, 0, 0, 11,
    -- filter=15 channel=51
    -7, -23, 0, -16, -8, -12, -13, -1, -16,
    -- filter=15 channel=52
    3, -10, 0, 9, -6, 0, 4, -1, 2,
    -- filter=15 channel=53
    5, 11, -3, -4, 0, 2, -10, 12, 1,
    -- filter=15 channel=54
    21, 15, 20, 25, 33, 24, 14, 4, 12,
    -- filter=15 channel=55
    -4, 5, 7, 0, 6, -6, 9, -3, -5,
    -- filter=15 channel=56
    -5, -3, 8, 0, -5, 4, -4, -7, -9,
    -- filter=15 channel=57
    0, 4, 2, -8, -5, 7, 8, 0, 2,
    -- filter=15 channel=58
    4, 13, 11, 8, -3, 4, -4, 2, -5,
    -- filter=15 channel=59
    2, -1, 6, 6, 5, 15, 1, 3, 12,
    -- filter=15 channel=60
    13, -5, -10, 7, -8, -10, -9, -17, 0,
    -- filter=15 channel=61
    -6, 2, -1, 5, -5, -8, -6, -9, -14,
    -- filter=15 channel=62
    10, 8, 13, -1, -1, 0, -4, 2, -2,
    -- filter=15 channel=63
    -7, -9, 4, -6, -5, 4, 0, 5, 0,
    -- filter=16 channel=0
    9, 17, 0, 21, 10, 18, 4, 13, 9,
    -- filter=16 channel=1
    -9, -3, 3, -12, -2, -4, -17, 4, -2,
    -- filter=16 channel=2
    -2, -6, 8, -15, -13, -4, -18, -15, -1,
    -- filter=16 channel=3
    -15, 1, -9, 1, 4, 0, -2, 3, -8,
    -- filter=16 channel=4
    13, 11, -7, 13, 3, 11, -5, 4, 4,
    -- filter=16 channel=5
    -10, -5, 9, 3, 7, 4, -4, 4, -2,
    -- filter=16 channel=6
    -5, -4, 8, -7, 8, 7, 8, -1, 7,
    -- filter=16 channel=7
    0, 5, 13, -5, 3, 12, -2, 3, 15,
    -- filter=16 channel=8
    10, 10, -5, 0, 18, 0, 5, 6, 8,
    -- filter=16 channel=9
    -25, -34, -36, -17, -37, -20, -15, -23, -33,
    -- filter=16 channel=10
    3, 13, 9, 9, 20, 20, 9, 19, 20,
    -- filter=16 channel=11
    -8, 1, -2, -2, 7, 3, -9, 2, 5,
    -- filter=16 channel=12
    -9, -1, -9, 8, 9, 2, 6, -8, 7,
    -- filter=16 channel=13
    -2, -9, -7, 9, 13, -4, -3, 8, 6,
    -- filter=16 channel=14
    -5, 0, 4, 3, 0, 12, -6, 3, -1,
    -- filter=16 channel=15
    12, 11, 0, 8, -1, 12, -4, 1, -6,
    -- filter=16 channel=16
    -12, -8, 0, -10, -8, -14, -20, -17, -2,
    -- filter=16 channel=17
    -8, 1, 2, 5, 8, 12, -10, 9, 10,
    -- filter=16 channel=18
    14, 4, -1, 17, 8, 8, 15, 2, -2,
    -- filter=16 channel=19
    0, -9, 7, -5, -16, 1, -8, -4, 4,
    -- filter=16 channel=20
    5, -9, 11, -1, 6, 0, 9, 5, 1,
    -- filter=16 channel=21
    8, 4, 6, 9, -2, 4, 2, -7, -5,
    -- filter=16 channel=22
    6, 5, 0, -4, -3, -3, 3, 5, -3,
    -- filter=16 channel=23
    5, 22, 13, 6, 10, 16, 6, 5, 4,
    -- filter=16 channel=24
    1, 0, -3, -3, 14, -5, 9, 11, 0,
    -- filter=16 channel=25
    -3, 0, -1, -16, -13, -8, -21, -14, -7,
    -- filter=16 channel=26
    9, 8, 13, 12, 6, -1, 0, -3, 6,
    -- filter=16 channel=27
    -13, 3, 7, -12, 6, 15, -9, -6, -3,
    -- filter=16 channel=28
    2, 0, -11, -2, 0, 0, -5, -12, -1,
    -- filter=16 channel=29
    -4, -9, -7, -1, -15, -13, -12, -19, -5,
    -- filter=16 channel=30
    4, 3, 6, -5, 21, 24, 10, 13, 22,
    -- filter=16 channel=31
    -2, -7, -8, 2, -5, 1, -6, 4, 5,
    -- filter=16 channel=32
    -11, 0, 13, -5, -1, 14, 6, 9, 6,
    -- filter=16 channel=33
    -2, -10, 9, 0, 0, 3, -6, -4, 2,
    -- filter=16 channel=34
    -2, 7, 11, -4, -1, 5, -7, 12, 3,
    -- filter=16 channel=35
    2, 22, 11, 8, 23, 18, 5, 0, 4,
    -- filter=16 channel=36
    9, 6, 3, 5, 10, -2, 11, -8, -2,
    -- filter=16 channel=37
    -14, -16, -18, -4, -18, 2, 0, -7, -14,
    -- filter=16 channel=38
    -11, 8, -6, 2, 13, 1, -8, -4, -6,
    -- filter=16 channel=39
    -9, 4, -1, 0, -3, -7, -3, -3, 6,
    -- filter=16 channel=40
    -4, 2, 3, 3, 9, -7, -7, 11, 11,
    -- filter=16 channel=41
    -2, 17, -1, 4, 9, -2, -13, -9, -7,
    -- filter=16 channel=42
    -8, -1, 0, 9, 9, -1, -4, 8, -9,
    -- filter=16 channel=43
    -12, 3, -3, 3, 7, 14, 7, -2, 7,
    -- filter=16 channel=44
    -12, 0, -5, -8, 1, 2, -1, -6, 0,
    -- filter=16 channel=45
    3, 0, 0, -3, -1, -7, 4, -10, 4,
    -- filter=16 channel=46
    -6, -5, -1, 13, 5, 8, -1, -7, 9,
    -- filter=16 channel=47
    -6, 0, -6, 3, 4, -10, 5, 5, 3,
    -- filter=16 channel=48
    7, -12, 0, -4, 0, 2, 1, -10, -10,
    -- filter=16 channel=49
    11, 11, 16, 16, 8, 20, 11, 6, 1,
    -- filter=16 channel=50
    0, 4, 1, -8, 2, 12, 11, 16, 6,
    -- filter=16 channel=51
    12, 20, 14, 12, 23, 5, 15, 24, 12,
    -- filter=16 channel=52
    10, -4, 0, 10, 4, 6, 5, -2, 0,
    -- filter=16 channel=53
    8, 16, 19, 3, 7, 5, 7, 4, 16,
    -- filter=16 channel=54
    -19, -27, -12, -21, -19, -18, -20, -11, -8,
    -- filter=16 channel=55
    -10, 8, -1, 6, -9, 1, -4, -10, 1,
    -- filter=16 channel=56
    0, -6, -4, 11, -5, -3, -3, 12, 12,
    -- filter=16 channel=57
    -5, 7, -8, 0, -2, -8, -8, 4, 7,
    -- filter=16 channel=58
    4, -7, 6, -1, 8, 8, 1, 9, 7,
    -- filter=16 channel=59
    2, -7, -1, -5, -2, 12, -16, -2, 7,
    -- filter=16 channel=60
    4, 18, -5, 5, 17, -2, -10, 4, 6,
    -- filter=16 channel=61
    11, 12, 0, 11, 26, 8, 3, 8, 4,
    -- filter=16 channel=62
    -2, -5, 2, -17, 0, -6, -12, 5, 4,
    -- filter=16 channel=63
    -8, 4, 4, 0, -4, -10, -10, 3, -6,
    -- filter=17 channel=0
    5, -7, 0, 7, -1, -7, 2, 3, 7,
    -- filter=17 channel=1
    0, -5, -8, -6, 7, 1, -5, 0, -8,
    -- filter=17 channel=2
    -5, -8, 2, 4, -9, -3, -3, 0, -8,
    -- filter=17 channel=3
    -3, -3, -4, 10, -2, 10, -2, 3, 0,
    -- filter=17 channel=4
    0, 5, -7, 5, 6, 0, -3, 2, -6,
    -- filter=17 channel=5
    -1, -9, -10, 2, -4, 3, 1, 9, -5,
    -- filter=17 channel=6
    1, -4, 5, 5, 9, -9, -9, -4, -7,
    -- filter=17 channel=7
    -1, -5, -6, 7, 0, -3, 5, 3, 8,
    -- filter=17 channel=8
    1, 8, 10, 6, -1, 3, 5, -1, -7,
    -- filter=17 channel=9
    6, -4, 2, -7, -2, -3, -10, 0, 4,
    -- filter=17 channel=10
    -3, -9, 8, 2, 8, 0, 8, 7, -5,
    -- filter=17 channel=11
    4, 0, -6, 0, 8, -8, 4, -2, -6,
    -- filter=17 channel=12
    6, 3, -8, 7, 6, 0, -1, -4, 7,
    -- filter=17 channel=13
    2, -2, 7, -9, 4, 5, 7, -5, 6,
    -- filter=17 channel=14
    0, 1, -5, -8, -5, -5, -6, 5, 2,
    -- filter=17 channel=15
    3, -3, -6, 1, 4, -9, -9, -10, 0,
    -- filter=17 channel=16
    7, -6, 3, -3, -6, 1, -3, -10, 0,
    -- filter=17 channel=17
    2, -2, -1, 2, 0, 1, 4, 10, 8,
    -- filter=17 channel=18
    2, 8, 6, 0, -9, 10, 1, 3, -7,
    -- filter=17 channel=19
    -8, -8, -8, 1, 8, 4, -9, -5, -5,
    -- filter=17 channel=20
    9, -8, 3, -2, 0, 4, 1, 1, -5,
    -- filter=17 channel=21
    -2, -8, -7, -8, -5, -8, -5, -9, 9,
    -- filter=17 channel=22
    0, 0, -5, -3, -7, 8, -2, 10, -7,
    -- filter=17 channel=23
    4, 3, 1, -7, 2, 7, 6, 4, 3,
    -- filter=17 channel=24
    -7, 0, -5, 0, 7, 9, -10, 0, 6,
    -- filter=17 channel=25
    -4, -6, -5, 1, 3, 8, 4, 7, 3,
    -- filter=17 channel=26
    -2, 3, -2, 2, -7, -1, 4, 8, -1,
    -- filter=17 channel=27
    4, 4, -6, -6, -2, 4, 5, 4, -3,
    -- filter=17 channel=28
    -7, -4, 3, 7, -9, -10, -6, -7, -7,
    -- filter=17 channel=29
    3, 9, -4, 3, -2, 2, 2, -6, -9,
    -- filter=17 channel=30
    -2, 8, 5, 7, 5, 7, -7, -7, 7,
    -- filter=17 channel=31
    -2, -4, 3, 3, 9, -8, 3, -5, 5,
    -- filter=17 channel=32
    -6, 5, 3, 3, -3, -1, -9, 7, -10,
    -- filter=17 channel=33
    -8, 5, 0, -4, 0, -2, -7, 0, 2,
    -- filter=17 channel=34
    5, -6, -4, -2, -9, 0, 10, -7, 0,
    -- filter=17 channel=35
    2, -5, -5, -8, -1, -10, 5, -8, -9,
    -- filter=17 channel=36
    -10, 5, 0, 8, -6, -1, 5, 3, 0,
    -- filter=17 channel=37
    9, 0, 0, 3, -1, -4, -10, -7, 3,
    -- filter=17 channel=38
    -9, 0, 0, -3, -1, -4, -7, 0, 10,
    -- filter=17 channel=39
    9, -6, 5, 1, -7, 5, 0, -10, 0,
    -- filter=17 channel=40
    -6, -8, -4, -3, 0, -3, 0, 9, 6,
    -- filter=17 channel=41
    2, 2, -1, -8, 10, 7, 0, 4, 1,
    -- filter=17 channel=42
    4, 0, 3, 8, 8, -8, 0, -4, -1,
    -- filter=17 channel=43
    7, 3, -6, 8, 8, -1, 6, -2, 0,
    -- filter=17 channel=44
    -4, 8, 1, -2, -6, 8, -9, -1, -1,
    -- filter=17 channel=45
    9, -5, -9, -3, -4, -6, -3, -6, 4,
    -- filter=17 channel=46
    10, 3, -1, 2, 3, 3, -3, 0, -5,
    -- filter=17 channel=47
    0, 6, 4, -7, -7, -7, -10, 5, -4,
    -- filter=17 channel=48
    3, 0, -5, -1, 6, 1, -6, 7, -4,
    -- filter=17 channel=49
    -6, -6, 1, -9, 0, 8, -2, -4, -4,
    -- filter=17 channel=50
    -8, 9, 2, 6, 1, 9, 9, 2, 8,
    -- filter=17 channel=51
    -2, -10, 3, 3, 2, 0, 7, 10, 5,
    -- filter=17 channel=52
    -1, -8, 6, 9, -7, 8, -5, -3, 6,
    -- filter=17 channel=53
    2, 0, 2, -4, -5, -3, -9, -10, 1,
    -- filter=17 channel=54
    1, 0, -4, -9, 1, 10, -7, 4, -4,
    -- filter=17 channel=55
    -2, 10, -4, -5, -3, 0, -3, 8, 6,
    -- filter=17 channel=56
    -7, -8, 9, -2, 0, 5, 5, 8, 4,
    -- filter=17 channel=57
    -7, 2, -5, -5, -4, -10, -8, 10, 6,
    -- filter=17 channel=58
    -3, -8, -1, -10, -2, 10, 3, -9, -9,
    -- filter=17 channel=59
    -7, 4, -2, -6, 9, -5, 6, 5, -2,
    -- filter=17 channel=60
    -7, -3, -5, -5, -10, -10, -9, 5, 4,
    -- filter=17 channel=61
    -4, -6, 0, 7, 5, 0, 0, -2, 4,
    -- filter=17 channel=62
    -1, -10, 9, 6, 3, 8, -10, 3, 1,
    -- filter=17 channel=63
    8, 0, -2, -6, 7, -2, 6, 4, 3,
    -- filter=18 channel=0
    -11, -22, -19, -14, -4, -18, -16, -8, -17,
    -- filter=18 channel=1
    10, 18, 24, 17, 20, 28, 9, 18, 25,
    -- filter=18 channel=2
    5, 28, 12, 19, 30, 14, 6, 23, 1,
    -- filter=18 channel=3
    23, 16, 15, 32, 19, 24, 29, 22, 16,
    -- filter=18 channel=4
    0, -3, -14, 2, 0, -16, 3, -14, -4,
    -- filter=18 channel=5
    10, 3, 13, 14, 18, 12, 4, 14, -7,
    -- filter=18 channel=6
    -8, 10, -2, 4, 0, -9, 5, -2, 1,
    -- filter=18 channel=7
    5, 1, -9, -6, 1, 0, 10, 11, -9,
    -- filter=18 channel=8
    4, 3, -14, -3, 1, -19, 0, -3, -19,
    -- filter=18 channel=9
    23, 33, 27, 17, 31, 34, 15, 31, 21,
    -- filter=18 channel=10
    -12, -8, 6, -5, -18, 0, 4, -4, 5,
    -- filter=18 channel=11
    -5, -6, 2, 5, -1, 5, 0, 4, -11,
    -- filter=18 channel=12
    12, 6, 9, -8, 2, 3, -5, -6, -5,
    -- filter=18 channel=13
    0, -8, -11, 5, -1, -6, 9, 0, -5,
    -- filter=18 channel=14
    2, -4, 7, 3, 1, 0, 8, 0, -8,
    -- filter=18 channel=15
    5, 6, -14, 13, 2, -4, -11, -4, -18,
    -- filter=18 channel=16
    19, 17, 11, 27, 26, 0, 12, 3, -11,
    -- filter=18 channel=17
    3, -12, -12, -5, -3, -11, -4, 4, -19,
    -- filter=18 channel=18
    -9, -8, -10, -6, -17, -5, -10, -12, -19,
    -- filter=18 channel=19
    23, 15, 13, 19, 38, 9, 7, 21, 10,
    -- filter=18 channel=20
    -5, 0, -3, 1, 3, -5, 1, 2, 0,
    -- filter=18 channel=21
    12, -1, 8, 11, -4, 2, -1, 6, -6,
    -- filter=18 channel=22
    9, 10, -5, 1, -5, 3, 7, 0, -10,
    -- filter=18 channel=23
    -9, -11, -10, -17, -5, 2, -12, -2, 1,
    -- filter=18 channel=24
    3, -5, -4, 1, 0, -18, -11, 4, -7,
    -- filter=18 channel=25
    12, 21, 23, 19, 35, 26, 23, 16, 22,
    -- filter=18 channel=26
    8, 14, 4, 12, 7, 4, 13, 5, 0,
    -- filter=18 channel=27
    2, 0, 0, -1, 10, 3, 9, 15, 9,
    -- filter=18 channel=28
    7, 18, -10, 20, 19, 0, 4, 14, -10,
    -- filter=18 channel=29
    6, 15, 6, 18, 14, -7, 14, 9, -2,
    -- filter=18 channel=30
    -1, 17, 4, 1, 27, -4, 14, 7, 5,
    -- filter=18 channel=31
    0, -5, -6, -5, 5, -2, 11, -9, -7,
    -- filter=18 channel=32
    -4, -4, 17, -6, 14, 13, 3, 5, 9,
    -- filter=18 channel=33
    -5, -7, 5, -4, -8, -6, 10, 2, -6,
    -- filter=18 channel=34
    6, 2, 5, 7, 4, -8, -5, 9, 1,
    -- filter=18 channel=35
    -18, 0, 13, -14, -7, 12, -10, 1, -2,
    -- filter=18 channel=36
    0, 3, 5, 0, 0, -6, 3, -9, 3,
    -- filter=18 channel=37
    8, 18, 13, 11, 30, 5, 14, 14, -1,
    -- filter=18 channel=38
    -8, -1, -7, 6, -4, -11, 14, 7, 0,
    -- filter=18 channel=39
    7, 1, 4, -5, -8, 8, 7, -3, -2,
    -- filter=18 channel=40
    -7, 4, -8, 10, -4, -3, 7, 5, -5,
    -- filter=18 channel=41
    14, 11, -3, -4, 4, 0, 9, -13, -4,
    -- filter=18 channel=42
    -4, 6, 0, -6, 2, 2, -3, 3, -6,
    -- filter=18 channel=43
    -13, -14, -13, 7, -4, -1, 0, -1, -8,
    -- filter=18 channel=44
    9, 8, 7, 15, 25, 18, 10, 6, 5,
    -- filter=18 channel=45
    9, 0, -4, -3, 6, -9, 9, 0, 2,
    -- filter=18 channel=46
    -1, 15, 9, 1, 13, 0, -1, 11, 2,
    -- filter=18 channel=47
    7, -5, 8, 7, -3, 4, -1, -5, 3,
    -- filter=18 channel=48
    0, 10, -3, 5, 0, 5, 10, -1, -10,
    -- filter=18 channel=49
    2, -18, -16, -4, -5, -15, -18, -8, -3,
    -- filter=18 channel=50
    -1, 4, -7, 2, 7, 5, 5, 2, 7,
    -- filter=18 channel=51
    -17, -20, -4, -20, -16, -22, -13, -27, 0,
    -- filter=18 channel=52
    11, -7, -10, -4, 3, 7, 11, 9, -8,
    -- filter=18 channel=53
    10, 3, 2, 0, 12, 0, 0, 22, 13,
    -- filter=18 channel=54
    24, 20, 23, 26, 33, 11, 19, 12, 0,
    -- filter=18 channel=55
    -5, 0, -10, 10, 9, -10, -2, 3, 1,
    -- filter=18 channel=56
    -1, 7, -6, 1, 6, -1, -6, -6, 4,
    -- filter=18 channel=57
    -9, 8, 0, -10, -9, -8, 2, -7, -4,
    -- filter=18 channel=58
    7, 2, 0, 15, 12, 1, 3, 13, 10,
    -- filter=18 channel=59
    24, 19, 16, 23, 3, 0, 10, 8, 7,
    -- filter=18 channel=60
    -4, -10, -17, 4, -5, -29, -9, -10, -24,
    -- filter=18 channel=61
    -16, -5, -21, -16, -21, -9, 4, -2, -16,
    -- filter=18 channel=62
    15, 14, 3, 22, 19, 9, 22, 9, 9,
    -- filter=18 channel=63
    9, 9, 8, -9, 2, -2, 6, 1, -3,
    -- filter=19 channel=0
    10, 4, -1, -1, -7, -9, 1, -3, -1,
    -- filter=19 channel=1
    -5, -5, 3, -8, -4, -8, 0, -3, 4,
    -- filter=19 channel=2
    -9, -9, 0, 2, 2, 3, -4, 0, 0,
    -- filter=19 channel=3
    2, -7, 8, -1, 1, 2, -3, 0, 0,
    -- filter=19 channel=4
    -5, 6, -1, -10, -8, 4, 7, -4, -6,
    -- filter=19 channel=5
    10, 5, -1, 2, -3, 0, -6, -5, 2,
    -- filter=19 channel=6
    8, 1, -6, 9, -4, 6, -2, 11, 4,
    -- filter=19 channel=7
    0, -7, 0, -8, 2, 4, 9, 7, 9,
    -- filter=19 channel=8
    6, -5, 1, 1, 0, -6, 0, -5, 9,
    -- filter=19 channel=9
    -6, -1, 8, 3, -4, -6, -1, 4, 10,
    -- filter=19 channel=10
    3, 1, -5, 9, 9, -1, 6, -4, 3,
    -- filter=19 channel=11
    -4, -5, 1, -10, -3, -2, 0, -5, 0,
    -- filter=19 channel=12
    4, 4, -3, 2, -7, 0, 0, -2, 1,
    -- filter=19 channel=13
    10, -3, 3, -1, 0, -3, -8, 0, 4,
    -- filter=19 channel=14
    5, -9, -8, -3, 8, 0, 1, 8, 3,
    -- filter=19 channel=15
    -3, -3, -1, -1, 6, -4, 10, 1, -2,
    -- filter=19 channel=16
    -10, 0, -5, 1, -4, 1, 8, -1, 0,
    -- filter=19 channel=17
    0, -4, -3, 7, -4, -3, -6, 2, -4,
    -- filter=19 channel=18
    11, -8, 10, 6, -5, -5, 11, 9, -4,
    -- filter=19 channel=19
    2, -7, 5, -5, -3, -3, -8, 2, 6,
    -- filter=19 channel=20
    -7, 1, 9, -7, 8, -4, 0, -9, 9,
    -- filter=19 channel=21
    7, 3, 1, 9, 10, 3, 5, 5, 10,
    -- filter=19 channel=22
    -6, -5, -4, -9, 8, -4, -6, 7, 1,
    -- filter=19 channel=23
    -3, -9, -2, -2, -5, -8, 4, 0, 3,
    -- filter=19 channel=24
    3, -3, -3, -9, 8, -6, -3, 2, -4,
    -- filter=19 channel=25
    1, 0, 0, 6, -9, 0, 10, 10, -2,
    -- filter=19 channel=26
    -6, 0, 7, -8, -7, -1, -3, -5, 5,
    -- filter=19 channel=27
    3, -3, 6, 0, -10, -4, -3, -9, -1,
    -- filter=19 channel=28
    5, 3, -8, 2, -8, -5, -9, -1, 0,
    -- filter=19 channel=29
    -11, -7, -8, 10, -4, 9, -5, 8, 6,
    -- filter=19 channel=30
    3, 7, -8, -10, 5, 2, 0, -4, -10,
    -- filter=19 channel=31
    0, 7, 0, 10, 5, -5, -7, 9, -2,
    -- filter=19 channel=32
    -10, 9, -9, -2, -6, -5, 4, 4, -1,
    -- filter=19 channel=33
    7, -6, -9, -9, -1, -7, 1, 7, 2,
    -- filter=19 channel=34
    -2, -5, -4, -6, -4, 4, -1, -2, -4,
    -- filter=19 channel=35
    -5, 0, 1, 4, -2, 4, -1, 8, 6,
    -- filter=19 channel=36
    -6, 10, 4, 11, 5, 9, 3, -7, 4,
    -- filter=19 channel=37
    6, -2, 8, 1, -5, 9, 7, 5, -1,
    -- filter=19 channel=38
    3, -7, -10, 2, -9, 8, -1, -8, -1,
    -- filter=19 channel=39
    -4, 6, -7, -9, -7, 4, 0, -3, 0,
    -- filter=19 channel=40
    9, -2, 10, -9, -7, 5, -8, 9, 5,
    -- filter=19 channel=41
    6, 5, -4, 1, -8, 8, 5, 4, 0,
    -- filter=19 channel=42
    -8, 5, 4, 7, -7, -10, 0, -7, -3,
    -- filter=19 channel=43
    -1, 1, -8, -1, 5, -9, 4, 3, 0,
    -- filter=19 channel=44
    -9, -1, -6, 9, -1, 7, -1, -4, 3,
    -- filter=19 channel=45
    7, -1, -8, -1, -1, -5, 0, -5, -1,
    -- filter=19 channel=46
    -10, -7, 7, 1, 7, 0, 9, 1, 3,
    -- filter=19 channel=47
    1, 10, -7, -4, 2, -2, -1, 9, 2,
    -- filter=19 channel=48
    1, 9, -3, 10, -4, -9, 4, 10, 10,
    -- filter=19 channel=49
    -8, -6, 4, 10, -7, 2, -5, -4, 3,
    -- filter=19 channel=50
    5, 3, -6, -1, -8, 10, -3, -1, -9,
    -- filter=19 channel=51
    4, 8, 5, 0, -1, 10, 0, 8, 8,
    -- filter=19 channel=52
    -6, 1, 0, 5, -2, 8, 4, 9, -9,
    -- filter=19 channel=53
    -9, 2, -1, -4, -9, 3, 4, 9, 5,
    -- filter=19 channel=54
    9, 3, -9, 7, -3, 3, -2, 6, 5,
    -- filter=19 channel=55
    -4, 3, 2, -1, -1, -2, -7, -9, -6,
    -- filter=19 channel=56
    9, -7, -2, -8, 5, -3, -3, 7, 5,
    -- filter=19 channel=57
    -5, -7, 5, -8, -5, -8, 1, 7, 6,
    -- filter=19 channel=58
    12, -3, -6, 1, -7, 9, 6, 4, -2,
    -- filter=19 channel=59
    -5, -2, -9, -3, 9, -7, -5, 7, -3,
    -- filter=19 channel=60
    -4, -7, -4, -4, -10, 8, 7, -7, 9,
    -- filter=19 channel=61
    -5, 5, 8, -2, -8, -1, -2, -3, -6,
    -- filter=19 channel=62
    -3, 0, -7, 1, 3, -7, 4, 8, -3,
    -- filter=19 channel=63
    4, -1, 7, 2, -1, 3, -1, -8, 10,
    -- filter=20 channel=0
    -3, -13, -9, 1, -5, -5, 8, 5, 5,
    -- filter=20 channel=1
    -13, -15, -10, -11, 1, 0, 3, -6, 5,
    -- filter=20 channel=2
    -18, -7, -3, -4, 1, 1, -17, -4, -10,
    -- filter=20 channel=3
    0, 0, 13, -12, 5, 8, 1, 10, 10,
    -- filter=20 channel=4
    11, -6, -6, 5, 2, 10, -2, -4, 9,
    -- filter=20 channel=5
    6, 8, 7, 2, 0, 14, 1, 7, 1,
    -- filter=20 channel=6
    7, 2, 0, -2, 9, 0, -3, -8, 1,
    -- filter=20 channel=7
    4, 7, -1, -4, 1, -1, -5, 0, 4,
    -- filter=20 channel=8
    -9, -5, 11, 0, 7, 5, -5, 2, -11,
    -- filter=20 channel=9
    37, 68, 61, 46, 78, 69, 36, 72, 69,
    -- filter=20 channel=10
    1, -11, 7, -1, 0, 0, 10, -7, 5,
    -- filter=20 channel=11
    -3, -7, -7, 4, 4, -9, -11, 3, 1,
    -- filter=20 channel=12
    3, 8, -4, 4, 9, 0, 7, 6, 6,
    -- filter=20 channel=13
    0, 16, 4, 8, 5, 11, 12, 2, 1,
    -- filter=20 channel=14
    0, -2, 8, 9, 0, -8, 6, -6, 6,
    -- filter=20 channel=15
    -4, 9, -4, -6, 8, 1, -10, 4, 6,
    -- filter=20 channel=16
    0, -5, -14, -3, 13, 0, -20, -5, -10,
    -- filter=20 channel=17
    -1, 8, -4, 2, 0, 3, 5, -10, -12,
    -- filter=20 channel=18
    10, 23, 21, 14, 29, 21, 9, 32, 14,
    -- filter=20 channel=19
    0, 20, 14, 14, 21, 10, 15, 21, 11,
    -- filter=20 channel=20
    10, 17, 16, 24, 23, 20, 21, 20, 19,
    -- filter=20 channel=21
    1, 0, 13, 11, 0, -3, 2, 7, 1,
    -- filter=20 channel=22
    5, -1, -10, 3, -10, -3, -4, 8, -1,
    -- filter=20 channel=23
    -3, -15, -13, -6, -11, -4, 6, -17, -11,
    -- filter=20 channel=24
    0, 0, 0, -3, 2, 3, 2, -9, 10,
    -- filter=20 channel=25
    -14, -7, -5, -8, -16, -20, -18, -25, -23,
    -- filter=20 channel=26
    6, 8, 10, 2, 4, 8, -6, 4, -5,
    -- filter=20 channel=27
    -11, -24, -3, -6, -11, -16, -18, -29, -15,
    -- filter=20 channel=28
    0, 17, 13, 16, 28, 9, 9, 4, 9,
    -- filter=20 channel=29
    5, 11, -11, -2, 22, 16, 1, 0, 3,
    -- filter=20 channel=30
    -9, -3, 0, -7, -12, 1, -4, -16, -9,
    -- filter=20 channel=31
    3, 10, 15, -2, 11, -7, 2, -5, -1,
    -- filter=20 channel=32
    11, -6, -1, -4, -12, -4, 0, 0, -10,
    -- filter=20 channel=33
    2, -1, -3, -7, 6, 10, 10, 0, 4,
    -- filter=20 channel=34
    -4, -5, 0, 8, 2, -8, -8, 1, 5,
    -- filter=20 channel=35
    -15, -17, -14, -23, -21, -30, -27, -21, -10,
    -- filter=20 channel=36
    10, 4, 9, 9, -6, 0, 14, 5, 4,
    -- filter=20 channel=37
    -1, 13, -5, 6, 9, 17, 4, 0, 6,
    -- filter=20 channel=38
    -18, -21, -3, -12, -13, -5, -10, -2, -1,
    -- filter=20 channel=39
    9, 8, 5, -2, 5, -4, -5, -5, 4,
    -- filter=20 channel=40
    4, -1, -8, -11, -13, -6, 1, 4, 3,
    -- filter=20 channel=41
    5, 4, -6, -2, -8, 2, -2, -20, -1,
    -- filter=20 channel=42
    -2, -4, 6, 0, 10, -3, -7, -5, -10,
    -- filter=20 channel=43
    -6, -18, -23, -13, -20, -17, 0, 3, -10,
    -- filter=20 channel=44
    -11, 6, 4, -12, -12, 2, 0, -15, 3,
    -- filter=20 channel=45
    -1, -3, 0, 3, 10, 9, 5, 9, -10,
    -- filter=20 channel=46
    0, 6, 0, 6, -2, -6, 4, 10, -1,
    -- filter=20 channel=47
    -9, -10, -3, -2, 0, -1, 0, -5, -3,
    -- filter=20 channel=48
    -2, 12, 9, -2, 7, 11, -5, 0, 13,
    -- filter=20 channel=49
    0, -10, 15, 4, 2, -7, 9, -16, 8,
    -- filter=20 channel=50
    -6, -9, 7, -6, -6, 0, 3, 0, 0,
    -- filter=20 channel=51
    14, -5, 5, -1, -3, 5, 0, 2, 7,
    -- filter=20 channel=52
    5, -9, 1, -8, -8, 10, 10, 5, -8,
    -- filter=20 channel=53
    -13, -12, -8, 1, -10, 4, -3, -2, 3,
    -- filter=20 channel=54
    20, 43, 28, 38, 42, 51, 19, 48, 45,
    -- filter=20 channel=55
    -7, 3, -7, -7, 8, 7, -4, 0, -9,
    -- filter=20 channel=56
    -4, -3, 8, -2, 7, 0, -6, 7, 10,
    -- filter=20 channel=57
    5, -7, 0, 8, 8, -4, 6, 7, 2,
    -- filter=20 channel=58
    10, 20, 5, 9, 15, 15, 17, 13, 11,
    -- filter=20 channel=59
    -4, -7, 0, -2, 0, -2, -13, -21, 2,
    -- filter=20 channel=60
    1, 0, -8, 11, 0, 1, -9, 4, 0,
    -- filter=20 channel=61
    0, -12, 1, 5, -3, -1, -4, -5, -12,
    -- filter=20 channel=62
    -8, -4, 0, -6, -4, -3, -1, 4, 6,
    -- filter=20 channel=63
    3, -6, -2, 8, 5, 0, -4, -3, 0,
    -- filter=21 channel=0
    11, 4, -2, 20, 23, 18, 9, 26, 17,
    -- filter=21 channel=1
    -1, -18, -17, -6, -22, -12, -9, -11, 0,
    -- filter=21 channel=2
    -10, -10, -10, 3, -22, -6, -13, -7, -12,
    -- filter=21 channel=3
    -1, -20, -16, -15, -6, -13, -15, -17, -10,
    -- filter=21 channel=4
    10, 15, 3, 11, 20, 7, 11, 17, 5,
    -- filter=21 channel=5
    -10, -8, 6, -12, -3, -4, 0, -15, -5,
    -- filter=21 channel=6
    0, 7, 3, 4, 12, 6, 10, 7, 9,
    -- filter=21 channel=7
    4, -6, 1, -11, -3, -9, 0, 2, 6,
    -- filter=21 channel=8
    5, 11, 2, 10, 26, 16, 17, 4, 4,
    -- filter=21 channel=9
    -14, -21, -15, 0, -31, -23, -12, -25, -26,
    -- filter=21 channel=10
    10, 14, 9, 11, 19, 13, 3, 9, 8,
    -- filter=21 channel=11
    9, 5, 6, -5, 4, 6, 14, 7, 5,
    -- filter=21 channel=12
    0, 10, 10, -3, 0, -4, -6, 8, 3,
    -- filter=21 channel=13
    1, 5, 0, 20, 7, 12, 16, 5, 10,
    -- filter=21 channel=14
    -7, 2, -3, 4, -11, 11, 7, 5, 12,
    -- filter=21 channel=15
    5, 6, 13, 1, 16, 6, 8, 0, 6,
    -- filter=21 channel=16
    -2, 2, 0, 0, 3, -8, -8, -12, -18,
    -- filter=21 channel=17
    11, 5, 4, 7, 2, 3, -1, 1, -1,
    -- filter=21 channel=18
    25, 11, 10, 31, 33, 9, 6, 24, 19,
    -- filter=21 channel=19
    -9, -14, -1, -13, -22, -19, -4, -19, -12,
    -- filter=21 channel=20
    -3, -2, 1, -5, 2, 1, 0, -3, -3,
    -- filter=21 channel=21
    -5, -5, 5, 2, -4, -1, 9, 7, -7,
    -- filter=21 channel=22
    -7, 2, -2, 4, 4, 7, -2, 0, -7,
    -- filter=21 channel=23
    11, 16, 4, 17, 21, 28, 15, 19, 27,
    -- filter=21 channel=24
    7, 8, 0, 0, 13, 1, 4, 5, -1,
    -- filter=21 channel=25
    -17, -20, -24, -11, -22, -26, -19, -14, -16,
    -- filter=21 channel=26
    -2, 2, -10, -3, -14, 2, 0, -13, 4,
    -- filter=21 channel=27
    2, 0, 2, 4, 5, 9, 1, 0, 2,
    -- filter=21 channel=28
    10, 5, -7, 2, -9, 0, 12, 0, 2,
    -- filter=21 channel=29
    9, -14, -12, 10, -8, -11, -5, -12, -15,
    -- filter=21 channel=30
    -2, 0, 10, -21, -3, 3, -15, -14, -5,
    -- filter=21 channel=31
    13, 2, 13, 0, 3, 9, -1, 13, 12,
    -- filter=21 channel=32
    -11, -2, 3, -11, -15, -12, -12, 4, 5,
    -- filter=21 channel=33
    4, -6, 0, 6, -4, 0, -2, 2, -9,
    -- filter=21 channel=34
    -9, -1, 0, -9, -7, -8, -2, 3, -10,
    -- filter=21 channel=35
    -7, -2, 14, -5, 14, 10, 8, 18, -3,
    -- filter=21 channel=36
    2, 11, 1, 3, 12, 10, 0, 9, -1,
    -- filter=21 channel=37
    -10, -3, -11, -10, -6, -12, 0, -17, -12,
    -- filter=21 channel=38
    12, 0, -9, 4, -3, 8, -1, 0, -7,
    -- filter=21 channel=39
    -8, 7, 8, -9, -3, -1, -1, -1, 4,
    -- filter=21 channel=40
    0, -9, -6, -1, -4, -11, -7, 7, 6,
    -- filter=21 channel=41
    0, 4, -2, 6, -4, 10, -1, 11, 7,
    -- filter=21 channel=42
    -8, -8, -1, 5, -9, 1, 4, -10, 6,
    -- filter=21 channel=43
    -26, -15, -21, -23, -20, -19, -18, -25, -16,
    -- filter=21 channel=44
    -4, -11, -9, -4, -15, -5, -4, -9, 0,
    -- filter=21 channel=45
    -9, 2, 2, 2, -3, 6, -1, 3, -3,
    -- filter=21 channel=46
    0, 5, -11, -7, 0, 2, -11, -3, -3,
    -- filter=21 channel=47
    6, -3, 1, 4, 10, 1, -1, 5, 8,
    -- filter=21 channel=48
    0, -3, -12, 5, 1, -4, -4, 5, -15,
    -- filter=21 channel=49
    6, 12, 18, 10, 17, 14, 6, 20, 13,
    -- filter=21 channel=50
    -16, -9, 0, -14, -3, -10, -6, -13, 10,
    -- filter=21 channel=51
    21, 25, 11, 28, 29, 16, 25, 31, 21,
    -- filter=21 channel=52
    -7, -7, -7, 7, 0, -9, -3, 10, 1,
    -- filter=21 channel=53
    -18, -18, -10, -11, -15, -6, -12, -8, 3,
    -- filter=21 channel=54
    -14, -15, -14, -16, -15, -16, -11, -17, -14,
    -- filter=21 channel=55
    2, -10, -10, 10, -5, 10, -4, 0, 0,
    -- filter=21 channel=56
    -6, 3, 5, 4, 3, 3, -6, 1, 6,
    -- filter=21 channel=57
    -3, 9, 6, -1, 1, -4, 5, -8, 5,
    -- filter=21 channel=58
    8, 6, 14, 0, 8, 4, 11, 12, 1,
    -- filter=21 channel=59
    -10, -11, -14, -15, -12, -9, -4, -9, -8,
    -- filter=21 channel=60
    19, 20, -2, 12, 27, 14, 17, 13, 5,
    -- filter=21 channel=61
    4, 14, 5, 14, 18, 18, 16, 15, 8,
    -- filter=21 channel=62
    2, -9, -3, -9, -16, -7, 2, -15, -10,
    -- filter=21 channel=63
    -3, -8, -6, 3, 1, 4, 5, -9, 2,
    -- filter=22 channel=0
    4, 5, 0, -4, -1, 8, 0, -6, 5,
    -- filter=22 channel=1
    0, 3, 15, -4, 11, 22, -6, 6, 7,
    -- filter=22 channel=2
    10, 3, 9, -8, 19, 17, -3, 16, 14,
    -- filter=22 channel=3
    15, 2, 16, -4, 4, 15, -5, -3, 9,
    -- filter=22 channel=4
    7, -10, -9, -9, -14, 4, -4, -15, -2,
    -- filter=22 channel=5
    11, 11, 4, -7, -1, 1, 5, 11, -6,
    -- filter=22 channel=6
    -1, 4, 12, -6, -2, -4, 8, 3, 0,
    -- filter=22 channel=7
    4, 7, -2, 3, 5, 5, 8, 2, 0,
    -- filter=22 channel=8
    6, 0, 0, -16, -15, 0, -17, 1, -2,
    -- filter=22 channel=9
    17, 15, 14, 9, 12, -1, 10, 8, -7,
    -- filter=22 channel=10
    -11, 5, 0, -10, -8, 11, 8, 0, -4,
    -- filter=22 channel=11
    7, -9, 0, 1, -6, 1, -6, 1, -3,
    -- filter=22 channel=12
    1, 3, 5, 0, -5, 0, -4, -5, -4,
    -- filter=22 channel=13
    -1, -4, 6, 1, 8, 3, 6, 1, -2,
    -- filter=22 channel=14
    10, 8, 1, 8, 1, 9, 4, 0, 8,
    -- filter=22 channel=15
    -9, 3, -6, 2, -12, -4, -4, -1, 0,
    -- filter=22 channel=16
    -2, 5, 19, -2, 11, 5, -1, 4, 0,
    -- filter=22 channel=17
    -4, 1, -1, -11, -3, 1, -12, -10, -5,
    -- filter=22 channel=18
    0, -12, 4, -7, -17, -11, -3, 3, -13,
    -- filter=22 channel=19
    15, 4, 7, 2, 15, 0, -3, 10, 1,
    -- filter=22 channel=20
    12, -3, 11, 3, 0, 3, 8, 6, -5,
    -- filter=22 channel=21
    4, -5, -10, -6, -10, 0, 8, 9, 2,
    -- filter=22 channel=22
    -9, -7, 0, 1, 4, -3, 5, 4, 2,
    -- filter=22 channel=23
    7, 1, -8, -6, -3, 8, 3, 0, -3,
    -- filter=22 channel=24
    1, -6, -1, 4, 0, -7, 1, -5, -1,
    -- filter=22 channel=25
    2, 11, 23, 5, 17, 29, -6, 11, 17,
    -- filter=22 channel=26
    8, 6, 12, 4, 12, 7, 7, 8, 0,
    -- filter=22 channel=27
    -6, 7, 16, -15, -8, 1, -11, -2, 16,
    -- filter=22 channel=28
    3, -5, -2, 0, -5, 5, 0, -1, -12,
    -- filter=22 channel=29
    14, -2, -3, 1, 6, 1, -8, -4, -1,
    -- filter=22 channel=30
    14, 21, 11, 7, 10, 14, 12, 8, 13,
    -- filter=22 channel=31
    5, 9, -8, 10, 8, 5, 1, -7, -5,
    -- filter=22 channel=32
    0, 8, -2, 5, 0, 16, 5, 3, 14,
    -- filter=22 channel=33
    -6, 4, 1, -10, 6, -4, -3, -2, -3,
    -- filter=22 channel=34
    -6, 4, 2, -6, 12, 10, -5, 1, -6,
    -- filter=22 channel=35
    -5, 0, 14, -3, 10, 19, 1, 0, 4,
    -- filter=22 channel=36
    -10, -5, 10, 5, -4, 0, -9, 10, 4,
    -- filter=22 channel=37
    11, 4, 3, 8, 14, 0, -7, 8, 7,
    -- filter=22 channel=38
    -4, 4, 5, -9, 2, 12, -5, -4, 7,
    -- filter=22 channel=39
    0, -1, -7, 1, -2, -5, 0, -8, 5,
    -- filter=22 channel=40
    0, 0, -4, 2, -7, -4, -4, 0, -6,
    -- filter=22 channel=41
    5, 0, 0, -12, 2, -4, -8, 1, 6,
    -- filter=22 channel=42
    7, 0, 5, 0, -7, -5, 2, 2, 1,
    -- filter=22 channel=43
    -1, 2, -3, 5, 15, 12, 5, 14, 12,
    -- filter=22 channel=44
    11, 19, 2, 4, 10, 6, 2, 11, 16,
    -- filter=22 channel=45
    2, 9, 0, 7, 0, 9, -7, -4, 2,
    -- filter=22 channel=46
    11, -6, 7, 13, 9, 11, -4, 8, 13,
    -- filter=22 channel=47
    -8, 5, -4, -9, 3, 2, -8, -1, -3,
    -- filter=22 channel=48
    -4, -4, 10, -4, -1, 9, -5, 11, 12,
    -- filter=22 channel=49
    -3, 7, 4, -10, -12, -11, 0, -5, 1,
    -- filter=22 channel=50
    0, 0, 2, 14, 9, 15, 15, 13, 0,
    -- filter=22 channel=51
    0, 0, -12, 3, -13, -14, -13, -14, -5,
    -- filter=22 channel=52
    -5, 6, -8, 9, -6, 3, -4, -9, -4,
    -- filter=22 channel=53
    1, 15, 2, 10, 7, 4, 7, 19, 6,
    -- filter=22 channel=54
    4, 6, -2, -5, -4, 0, 1, -6, 2,
    -- filter=22 channel=55
    -1, -2, -3, -4, 0, -4, -2, -2, -8,
    -- filter=22 channel=56
    0, 11, -8, 7, 6, -5, -6, -3, 1,
    -- filter=22 channel=57
    -5, 0, -2, 8, 6, 7, -9, 0, 8,
    -- filter=22 channel=58
    -1, 10, -6, 14, -5, 8, 0, -5, 11,
    -- filter=22 channel=59
    4, -2, 13, 4, 12, 6, -1, 9, 11,
    -- filter=22 channel=60
    6, -11, -1, -14, -10, 0, -22, -14, -6,
    -- filter=22 channel=61
    3, -1, -11, -17, -14, -8, -12, -18, -8,
    -- filter=22 channel=62
    -7, 15, 9, -3, 13, -3, -6, -7, 4,
    -- filter=22 channel=63
    -2, 1, -4, 0, 9, 3, -7, -1, -4,
    -- filter=23 channel=0
    -4, 5, -3, -1, -4, 7, -13, -2, -3,
    -- filter=23 channel=1
    -16, -5, -1, -15, 3, 16, -12, -6, 14,
    -- filter=23 channel=2
    3, 0, 20, -14, 0, 10, -19, -22, -7,
    -- filter=23 channel=3
    -4, 19, 5, 4, 4, 21, -12, -3, 0,
    -- filter=23 channel=4
    -9, 2, 12, 3, 12, 10, -3, -7, -7,
    -- filter=23 channel=5
    9, 8, 5, 2, 0, 10, 0, -9, 9,
    -- filter=23 channel=6
    -7, -3, 12, 0, 11, 1, -12, -17, -1,
    -- filter=23 channel=7
    -2, 5, 11, -5, -2, 9, 10, 4, 2,
    -- filter=23 channel=8
    3, 19, 36, -6, 10, 25, -14, -17, -12,
    -- filter=23 channel=9
    -3, 31, 26, -4, 33, 37, -1, 2, 20,
    -- filter=23 channel=10
    -5, -17, 1, -9, -4, -5, -4, 4, 9,
    -- filter=23 channel=11
    -12, 2, 7, -5, -2, 18, -14, -3, -7,
    -- filter=23 channel=12
    -3, 6, 4, 8, -3, 9, -7, 4, -5,
    -- filter=23 channel=13
    12, 4, 9, 13, 29, 23, -14, -2, 12,
    -- filter=23 channel=14
    9, 3, 0, -2, -4, 0, -5, 8, -5,
    -- filter=23 channel=15
    4, 31, 16, -9, 21, 32, -16, -22, -3,
    -- filter=23 channel=16
    6, 29, 43, -4, 3, 38, -41, -18, 0,
    -- filter=23 channel=17
    -3, 0, 7, 4, 8, 14, -11, -14, -6,
    -- filter=23 channel=18
    5, 13, 10, -2, 5, 0, -7, 0, 6,
    -- filter=23 channel=19
    -4, 4, 1, 6, -1, 12, 0, -5, -1,
    -- filter=23 channel=20
    8, 18, -1, 9, 7, 5, 10, 19, 8,
    -- filter=23 channel=21
    11, 4, 3, 10, -7, 5, 0, 2, -5,
    -- filter=23 channel=22
    1, 2, 5, 0, 1, 6, 4, -9, 9,
    -- filter=23 channel=23
    -14, -22, 3, -15, -1, -6, 0, -4, -6,
    -- filter=23 channel=24
    -10, -1, 7, 8, 4, 16, -1, -12, -6,
    -- filter=23 channel=25
    1, 2, 13, -2, -11, 19, -29, -25, -1,
    -- filter=23 channel=26
    6, 9, -4, 6, 17, 1, 5, 13, 13,
    -- filter=23 channel=27
    -1, 13, 9, -14, 0, 8, -10, -26, -4,
    -- filter=23 channel=28
    1, 16, 25, 0, 15, 22, -22, -25, -15,
    -- filter=23 channel=29
    13, 32, 42, -1, 27, 39, -35, -16, -4,
    -- filter=23 channel=30
    -4, 6, 7, 6, -7, 3, 17, 0, -6,
    -- filter=23 channel=31
    6, -10, -4, 5, 5, 5, -6, 0, 9,
    -- filter=23 channel=32
    6, -8, -11, -11, -2, 1, -11, -1, -7,
    -- filter=23 channel=33
    -9, -5, 9, -9, -2, -6, -1, -9, 0,
    -- filter=23 channel=34
    4, 0, -1, 12, 9, 6, -3, 3, 5,
    -- filter=23 channel=35
    -2, -2, -2, -13, -9, 0, -24, -21, -5,
    -- filter=23 channel=36
    -2, -12, -13, -2, 7, 5, -4, -2, -8,
    -- filter=23 channel=37
    5, 6, 16, 11, 18, 1, 0, -3, -8,
    -- filter=23 channel=38
    -6, 8, 24, -11, 7, 26, -18, -21, 10,
    -- filter=23 channel=39
    -4, 2, -4, 2, 10, 9, 4, 1, -6,
    -- filter=23 channel=40
    5, -10, -7, 7, -7, 3, -8, -2, -6,
    -- filter=23 channel=41
    2, 14, 35, -10, 5, 22, -31, -25, -11,
    -- filter=23 channel=42
    2, 3, 6, 4, 1, -7, 10, 2, -10,
    -- filter=23 channel=43
    1, -20, -19, 18, 8, 0, 20, 12, 2,
    -- filter=23 channel=44
    4, -3, 8, -11, -13, 10, 2, -2, 0,
    -- filter=23 channel=45
    8, -2, 0, 9, -3, 9, 9, -5, -8,
    -- filter=23 channel=46
    3, 0, 15, 22, 8, -1, -4, 0, 4,
    -- filter=23 channel=47
    -6, 5, 5, -2, -5, 5, -6, -1, -8,
    -- filter=23 channel=48
    12, 6, 20, -2, 18, 19, -3, 1, -2,
    -- filter=23 channel=49
    8, 2, 4, 2, -11, -15, -16, -3, -1,
    -- filter=23 channel=50
    1, -2, -6, 14, 10, -3, 11, 6, -6,
    -- filter=23 channel=51
    4, -9, 0, 0, -12, -14, 13, 0, 7,
    -- filter=23 channel=52
    1, 7, -11, -8, 0, 5, -1, 0, 6,
    -- filter=23 channel=53
    -9, 7, 1, 7, 2, -4, -4, -7, 0,
    -- filter=23 channel=54
    -6, 21, 25, -6, 24, 10, -12, -7, 8,
    -- filter=23 channel=55
    5, -3, 0, 0, -6, -8, 7, -7, -9,
    -- filter=23 channel=56
    -10, 4, -1, -3, 10, 3, 3, 10, -3,
    -- filter=23 channel=57
    -6, 5, -8, 6, -4, 7, 0, 4, 1,
    -- filter=23 channel=58
    -7, 2, 3, 2, 0, -12, -7, 14, 11,
    -- filter=23 channel=59
    0, 17, 31, -4, -7, 18, -27, -24, 0,
    -- filter=23 channel=60
    16, 30, 28, 4, 16, 45, -21, -21, 5,
    -- filter=23 channel=61
    -3, 8, 20, -14, 10, 25, -23, -27, 4,
    -- filter=23 channel=62
    -2, 0, 12, -1, 4, 15, -3, -10, -3,
    -- filter=23 channel=63
    0, -7, -8, 7, -6, 7, 1, 2, -9,
    -- filter=24 channel=0
    1, -9, 2, 0, 6, -4, -7, 8, 9,
    -- filter=24 channel=1
    -8, 5, -7, -7, 4, 0, 2, 1, 6,
    -- filter=24 channel=2
    6, 4, 3, -1, -4, 5, -6, -7, 8,
    -- filter=24 channel=3
    -4, 6, 1, 1, 5, 3, -5, -5, -1,
    -- filter=24 channel=4
    7, -6, 8, 7, -7, 1, 6, 7, -2,
    -- filter=24 channel=5
    -1, -7, -8, 1, -3, 3, 0, 0, 4,
    -- filter=24 channel=6
    -3, -5, -6, 5, -6, 3, 9, 8, -9,
    -- filter=24 channel=7
    5, -4, 6, -6, 6, 9, 7, 0, 1,
    -- filter=24 channel=8
    5, 0, -5, -1, 10, -10, -4, 2, 7,
    -- filter=24 channel=9
    -9, -6, 1, -3, -5, -2, 8, -1, -6,
    -- filter=24 channel=10
    -3, 7, 0, 8, -5, 5, 5, 5, 6,
    -- filter=24 channel=11
    8, -1, 0, -2, 9, -9, -3, 10, 2,
    -- filter=24 channel=12
    3, 0, -9, -2, 0, 1, 0, 2, 1,
    -- filter=24 channel=13
    2, 0, -1, -6, 5, -9, 1, 2, 0,
    -- filter=24 channel=14
    -5, 1, 7, -4, 1, 5, -2, 6, -10,
    -- filter=24 channel=15
    -11, -9, 4, -7, 7, -9, -9, -7, -9,
    -- filter=24 channel=16
    2, 0, -9, 2, -4, -7, -3, 4, 1,
    -- filter=24 channel=17
    5, 8, 9, 2, -5, -8, 10, -7, 1,
    -- filter=24 channel=18
    -9, -2, 8, -6, 4, -5, -1, -7, 7,
    -- filter=24 channel=19
    -7, 9, -6, 1, -8, 6, 6, 2, -4,
    -- filter=24 channel=20
    4, -4, -6, 4, 3, -1, 0, 2, 9,
    -- filter=24 channel=21
    0, 7, 2, 1, 9, -6, 6, 2, -2,
    -- filter=24 channel=22
    -3, -3, -4, -3, 7, -3, -2, -6, 1,
    -- filter=24 channel=23
    -5, -1, 10, 0, 7, 9, 2, -3, 9,
    -- filter=24 channel=24
    -9, -6, -6, 2, 4, -5, -5, -10, 8,
    -- filter=24 channel=25
    -9, -6, 3, -2, -5, -7, 0, -1, 5,
    -- filter=24 channel=26
    8, 6, -7, -5, 8, -1, 3, 10, -4,
    -- filter=24 channel=27
    6, 1, 3, 11, -5, 2, 2, 5, 10,
    -- filter=24 channel=28
    -6, 3, 7, -8, -4, 7, 4, -8, 8,
    -- filter=24 channel=29
    2, -7, -1, -7, 5, 6, -9, -3, 0,
    -- filter=24 channel=30
    -4, 4, -7, -8, 1, -5, 4, -4, 7,
    -- filter=24 channel=31
    2, -7, 0, -9, 0, -6, 7, -5, -1,
    -- filter=24 channel=32
    -5, -7, -1, 9, 5, 10, 0, 0, -1,
    -- filter=24 channel=33
    8, 9, 9, 8, 0, -9, 9, 6, 3,
    -- filter=24 channel=34
    -2, 9, 5, 10, -1, -6, 1, 6, -8,
    -- filter=24 channel=35
    11, -1, 12, 4, 10, -1, 6, 1, 7,
    -- filter=24 channel=36
    4, -5, 10, -6, 7, 1, 0, 1, 8,
    -- filter=24 channel=37
    -1, -7, 6, 2, 1, 1, 0, -2, 1,
    -- filter=24 channel=38
    -6, 3, 9, 10, 10, 2, 3, 7, 12,
    -- filter=24 channel=39
    4, -4, 7, -7, 9, -10, -4, 0, 10,
    -- filter=24 channel=40
    -8, -6, 8, -9, 8, 3, 4, -5, 8,
    -- filter=24 channel=41
    0, -1, 3, 0, -10, -9, 3, 10, -2,
    -- filter=24 channel=42
    9, 4, 4, -6, 0, -4, 10, -5, 1,
    -- filter=24 channel=43
    7, 0, -10, -10, -3, -3, -10, 3, 0,
    -- filter=24 channel=44
    8, -3, 2, -1, 0, 1, 4, -7, 4,
    -- filter=24 channel=45
    -1, 4, 1, -1, -10, -3, -9, 7, 1,
    -- filter=24 channel=46
    9, -4, -5, -6, -9, 1, 7, -7, -5,
    -- filter=24 channel=47
    5, 8, 2, -9, 4, -5, -5, -10, -5,
    -- filter=24 channel=48
    -6, -4, -8, -7, -8, 8, 3, -10, -2,
    -- filter=24 channel=49
    5, -6, -6, 7, 7, -1, -5, 2, -1,
    -- filter=24 channel=50
    8, 0, 7, 5, 0, -1, 5, 10, -4,
    -- filter=24 channel=51
    0, 7, -6, 1, -6, 3, 2, -3, 10,
    -- filter=24 channel=52
    0, -4, 9, 0, -9, 2, 6, 1, 10,
    -- filter=24 channel=53
    10, 7, -1, 4, 7, -7, -7, -5, 8,
    -- filter=24 channel=54
    4, 2, 8, 5, 4, -9, 10, 8, -6,
    -- filter=24 channel=55
    3, 6, -1, -5, -5, -9, 6, 0, 7,
    -- filter=24 channel=56
    0, -7, 5, 0, -5, -2, 3, 6, 0,
    -- filter=24 channel=57
    -10, 5, -3, 8, -6, -9, -9, -2, 1,
    -- filter=24 channel=58
    2, -4, -4, -4, -9, 0, 1, -3, 1,
    -- filter=24 channel=59
    0, 1, 4, 10, -8, -1, 0, 5, -8,
    -- filter=24 channel=60
    -11, -8, 2, -7, 5, 9, 0, -7, -4,
    -- filter=24 channel=61
    -10, -3, -7, -2, -4, -6, -8, -4, 8,
    -- filter=24 channel=62
    1, 0, 10, 5, -9, 9, 7, 2, -2,
    -- filter=24 channel=63
    1, 5, -8, -1, 5, -8, -6, 1, -7,
    -- filter=25 channel=0
    -17, -1, -19, 0, 8, 3, -5, 15, -8,
    -- filter=25 channel=1
    -8, -12, -14, -8, 13, 10, -5, 17, 5,
    -- filter=25 channel=2
    -1, 0, -13, 9, 19, -3, -6, -2, -3,
    -- filter=25 channel=3
    7, 18, 4, 23, 9, 12, 19, 5, 7,
    -- filter=25 channel=4
    -2, -5, -9, -8, 16, -8, -2, 0, 3,
    -- filter=25 channel=5
    4, 13, -2, 6, 11, 1, -3, 8, -4,
    -- filter=25 channel=6
    2, 0, -1, -5, 2, 0, 0, -6, -8,
    -- filter=25 channel=7
    5, 7, 11, -5, 3, 11, 0, -5, -1,
    -- filter=25 channel=8
    0, 13, -3, 10, 22, 8, -9, -2, -9,
    -- filter=25 channel=9
    0, -8, -20, 12, -13, -27, 4, -4, -27,
    -- filter=25 channel=10
    -17, -7, 0, -9, 6, 11, 2, 0, -1,
    -- filter=25 channel=11
    -14, 2, 3, -13, 5, -6, -1, 17, 9,
    -- filter=25 channel=12
    2, 6, 2, 1, -6, -3, 5, -9, 11,
    -- filter=25 channel=13
    -9, -7, -25, 15, -3, -6, 0, -1, -12,
    -- filter=25 channel=14
    -2, -1, 10, 3, 1, 0, -4, 5, 13,
    -- filter=25 channel=15
    -7, 0, -15, 11, 10, 1, -7, 7, -1,
    -- filter=25 channel=16
    10, 0, -17, 24, 13, 7, 9, 2, -2,
    -- filter=25 channel=17
    -2, -4, 5, 7, 23, 5, -3, 7, 3,
    -- filter=25 channel=18
    -7, 6, -3, 2, 5, -5, 0, -6, -12,
    -- filter=25 channel=19
    -8, -1, 5, 8, -6, 9, -6, 6, 0,
    -- filter=25 channel=20
    1, -9, 2, -6, -6, -15, 1, -4, -1,
    -- filter=25 channel=21
    -5, -2, 9, -5, 6, 4, 0, -4, 5,
    -- filter=25 channel=22
    6, -6, 6, -8, 7, 4, -4, -7, -7,
    -- filter=25 channel=23
    -7, -2, 11, -12, 7, 15, -11, 18, 3,
    -- filter=25 channel=24
    -6, -1, -12, -5, 8, 4, -4, 5, 0,
    -- filter=25 channel=25
    -4, 0, -5, 0, 16, 3, -13, 14, -5,
    -- filter=25 channel=26
    -5, 7, 1, -5, -10, -11, 2, -4, 0,
    -- filter=25 channel=27
    -10, 17, -7, 4, 16, 6, 4, 16, 1,
    -- filter=25 channel=28
    -3, 2, -9, 1, 5, -5, -12, -1, 0,
    -- filter=25 channel=29
    13, 4, -31, 20, 18, -7, 17, -4, -25,
    -- filter=25 channel=30
    -1, 12, 0, -8, 12, 15, 9, 2, 10,
    -- filter=25 channel=31
    -4, 3, -3, 7, 5, -5, -3, 10, -3,
    -- filter=25 channel=32
    -15, 1, 3, -15, 0, 10, 2, 9, 17,
    -- filter=25 channel=33
    4, 2, -5, 3, 1, 0, 1, 0, 7,
    -- filter=25 channel=34
    6, 2, 7, -6, 12, -4, 12, 10, -2,
    -- filter=25 channel=35
    -13, 13, 2, -6, 21, 10, -17, -1, 4,
    -- filter=25 channel=36
    3, 1, 12, -8, 8, 0, -4, 7, -7,
    -- filter=25 channel=37
    0, -3, -13, 9, 3, 0, 8, 9, 0,
    -- filter=25 channel=38
    -11, 3, -17, -1, 23, 11, 2, 20, 8,
    -- filter=25 channel=39
    1, -8, -4, 5, 3, -5, -7, -7, 0,
    -- filter=25 channel=40
    1, -3, 6, -6, -7, -2, -10, 8, -8,
    -- filter=25 channel=41
    -5, 13, -11, 7, 33, 12, 1, 1, 0,
    -- filter=25 channel=42
    7, 9, 3, 3, -7, -7, 8, -9, 2,
    -- filter=25 channel=43
    -10, -31, -21, -23, -20, -4, 0, 6, -1,
    -- filter=25 channel=44
    -4, 0, 17, -12, 1, 18, -14, 5, 7,
    -- filter=25 channel=45
    2, 6, 9, -2, -4, -3, -5, -2, 0,
    -- filter=25 channel=46
    13, 3, 6, 0, -8, -9, -4, 2, 4,
    -- filter=25 channel=47
    1, 3, 5, -10, -6, -10, -6, -3, -6,
    -- filter=25 channel=48
    7, -11, -9, 17, -4, -11, 7, 5, -1,
    -- filter=25 channel=49
    -5, 4, -3, 4, 17, 5, -17, 8, -6,
    -- filter=25 channel=50
    -3, -14, 0, 0, -7, 5, -7, 11, 6,
    -- filter=25 channel=51
    -7, -5, 7, -12, -10, -6, 0, 0, -3,
    -- filter=25 channel=52
    -2, 2, -6, -9, 8, 10, 0, -8, -7,
    -- filter=25 channel=53
    -9, 13, 8, -9, 3, 18, -10, -1, 6,
    -- filter=25 channel=54
    -1, 3, -10, 14, -8, -18, 2, -8, -24,
    -- filter=25 channel=55
    -3, 5, 10, 0, 5, -3, -2, 7, 6,
    -- filter=25 channel=56
    1, 3, 0, 11, 6, 1, 0, 9, -7,
    -- filter=25 channel=57
    7, -10, -8, 0, 7, -2, -4, 3, 7,
    -- filter=25 channel=58
    1, 2, 11, -8, -12, 2, 3, 7, 2,
    -- filter=25 channel=59
    -1, 6, -9, 23, 12, 2, 5, 11, 5,
    -- filter=25 channel=60
    3, 12, -28, 4, 36, 4, 19, 31, -8,
    -- filter=25 channel=61
    -3, 3, -15, -1, 24, 14, -10, 23, 16,
    -- filter=25 channel=62
    16, 1, 1, -1, 21, 4, -3, 9, 8,
    -- filter=25 channel=63
    -7, 0, -2, 3, -6, -1, 9, 2, 10,
    -- filter=26 channel=0
    -2, 15, 9, 0, 17, 8, 3, 19, 8,
    -- filter=26 channel=1
    5, -10, 7, 0, -5, 0, -5, -4, 0,
    -- filter=26 channel=2
    -14, -2, -9, -4, 8, -8, -8, 8, 11,
    -- filter=26 channel=3
    5, -2, 6, -2, -6, 7, -1, 5, 8,
    -- filter=26 channel=4
    0, 2, -5, -9, 11, -3, 0, 6, 9,
    -- filter=26 channel=5
    -10, 4, 5, -1, -10, 5, 6, -6, 7,
    -- filter=26 channel=6
    -5, -8, -4, 4, 13, 12, 3, -3, 4,
    -- filter=26 channel=7
    2, -8, 9, -8, -1, 2, 5, 6, -7,
    -- filter=26 channel=8
    0, -7, -2, 0, -1, -8, -4, 4, 4,
    -- filter=26 channel=9
    -13, -11, -12, -19, -24, -8, 0, -13, 0,
    -- filter=26 channel=10
    0, 11, 11, 16, 18, 6, 8, 13, 20,
    -- filter=26 channel=11
    6, -6, -11, 6, 9, -6, -8, 9, 6,
    -- filter=26 channel=12
    7, -8, 5, -8, 10, 6, 5, 1, 9,
    -- filter=26 channel=13
    -1, -13, -5, -1, 7, -10, 0, -3, 7,
    -- filter=26 channel=14
    -2, 8, -10, -3, -2, -1, -3, 5, 2,
    -- filter=26 channel=15
    -10, -4, -9, 8, 0, 5, -1, 8, 13,
    -- filter=26 channel=16
    -15, -13, -1, -9, -20, -15, -12, -8, 0,
    -- filter=26 channel=17
    -15, -8, -6, -13, 10, -5, 2, 2, -6,
    -- filter=26 channel=18
    16, 2, 16, 2, 18, 7, 14, 15, -2,
    -- filter=26 channel=19
    -11, -1, 3, -7, 2, 4, -14, 3, 6,
    -- filter=26 channel=20
    -6, 0, 4, 0, -9, 1, 11, -4, 0,
    -- filter=26 channel=21
    1, 0, 6, 4, -5, 8, 5, 6, -5,
    -- filter=26 channel=22
    -9, 0, 4, 0, -5, -9, 4, 9, -5,
    -- filter=26 channel=23
    1, 18, 8, 19, 18, 5, 2, 23, 21,
    -- filter=26 channel=24
    -11, 4, -3, 3, 1, -2, 4, 1, 3,
    -- filter=26 channel=25
    -10, -9, 0, -11, 5, 9, -7, 4, 11,
    -- filter=26 channel=26
    8, -10, 1, 7, -4, 4, 4, 8, 8,
    -- filter=26 channel=27
    4, -6, -1, 2, 10, 2, 0, 15, 16,
    -- filter=26 channel=28
    -2, -11, -12, -16, -8, -10, -11, -8, 0,
    -- filter=26 channel=29
    -18, -25, -19, -20, -18, -6, -1, -15, -5,
    -- filter=26 channel=30
    -4, -11, -10, 2, -4, 2, -7, 7, 6,
    -- filter=26 channel=31
    7, 5, 13, 12, 9, 13, -1, 6, 4,
    -- filter=26 channel=32
    0, -2, -6, -1, 9, 0, -4, 2, -5,
    -- filter=26 channel=33
    0, 8, -8, -3, 9, 1, -3, 0, -7,
    -- filter=26 channel=34
    -5, -7, 5, -1, -10, 10, 9, 5, -6,
    -- filter=26 channel=35
    18, 16, 12, 1, 24, 14, 14, 7, 3,
    -- filter=26 channel=36
    -2, 0, 6, 13, 9, -4, 0, 11, -3,
    -- filter=26 channel=37
    -3, -5, -10, -10, -12, 4, -13, 6, 4,
    -- filter=26 channel=38
    -4, -4, 7, 5, 8, 5, 8, 10, 10,
    -- filter=26 channel=39
    1, 1, -2, -2, -4, 1, 2, 9, 2,
    -- filter=26 channel=40
    -2, 5, -6, 5, 2, 6, 5, -4, 12,
    -- filter=26 channel=41
    -13, -13, -4, -4, -3, -1, -10, 7, 0,
    -- filter=26 channel=42
    -4, 5, -1, -7, 6, -2, 4, 2, 8,
    -- filter=26 channel=43
    5, 8, 10, -10, -10, 4, -5, -11, -6,
    -- filter=26 channel=44
    2, 0, -1, 0, 3, 8, 8, -3, -7,
    -- filter=26 channel=45
    -7, 6, -3, 0, 3, 8, 1, 3, 0,
    -- filter=26 channel=46
    1, 3, 4, -1, 7, 0, 4, 0, -6,
    -- filter=26 channel=47
    8, 5, -2, -5, -7, -6, 5, -2, -2,
    -- filter=26 channel=48
    6, 4, -5, -8, -2, -9, -5, 3, 3,
    -- filter=26 channel=49
    13, 1, 5, 14, 12, 21, 1, 6, 16,
    -- filter=26 channel=50
    -8, 6, -6, -2, 5, 2, -2, -11, 2,
    -- filter=26 channel=51
    21, 24, 5, 21, 15, 21, 23, 23, 16,
    -- filter=26 channel=52
    7, 10, 8, 11, 0, 10, 1, -9, 6,
    -- filter=26 channel=53
    -9, -7, 0, 7, 8, 0, -5, -2, 6,
    -- filter=26 channel=54
    -16, -1, -9, -14, -8, -19, -1, -2, 0,
    -- filter=26 channel=55
    0, 9, 0, 9, 0, 0, 0, -8, -5,
    -- filter=26 channel=56
    -3, 4, -6, -8, 4, -9, 4, 6, 0,
    -- filter=26 channel=57
    3, -6, 0, 6, -1, -6, 4, -2, -3,
    -- filter=26 channel=58
    1, 12, 2, 11, -3, 5, 16, 6, 13,
    -- filter=26 channel=59
    -8, -6, 5, 1, -6, 10, 0, 10, 0,
    -- filter=26 channel=60
    -10, -1, 1, 5, -10, 11, 5, 2, -1,
    -- filter=26 channel=61
    -3, 0, -3, -12, -5, 1, 6, 1, 17,
    -- filter=26 channel=62
    -7, -10, 2, -7, -7, 5, 2, -4, -1,
    -- filter=26 channel=63
    -9, -3, -9, 6, 5, -2, -9, 1, -9,
    -- filter=27 channel=0
    -19, -8, 0, 1, 1, 1, -9, 13, 6,
    -- filter=27 channel=1
    -15, 5, 2, -7, 10, 23, -2, 12, 17,
    -- filter=27 channel=2
    5, 19, 24, 3, 27, 23, -6, -1, 10,
    -- filter=27 channel=3
    5, 9, 23, 24, 33, 16, 7, 12, 17,
    -- filter=27 channel=4
    -10, 2, -11, -12, 4, -4, -12, -13, 6,
    -- filter=27 channel=5
    0, 9, 9, 0, -4, 7, 3, 3, -4,
    -- filter=27 channel=6
    -8, 1, 0, 0, 5, 2, -9, 1, 9,
    -- filter=27 channel=7
    -5, -10, -8, -3, -10, 0, -8, 2, -10,
    -- filter=27 channel=8
    -3, 5, 0, -12, 11, 30, -19, 4, -4,
    -- filter=27 channel=9
    0, -16, -18, -5, -6, -19, 4, -13, -7,
    -- filter=27 channel=10
    -6, 2, -10, -8, 0, -2, -3, -5, 12,
    -- filter=27 channel=11
    -16, -9, 1, -7, 7, 19, -14, 0, 16,
    -- filter=27 channel=12
    -1, 2, 3, 0, 0, 5, -5, 2, 10,
    -- filter=27 channel=13
    -12, -15, -11, 1, 0, -6, 10, 9, 17,
    -- filter=27 channel=14
    8, -3, -1, -12, 4, 0, -6, 3, -1,
    -- filter=27 channel=15
    3, 4, 7, 2, 23, 10, -15, 8, 1,
    -- filter=27 channel=16
    0, 3, 4, -1, 34, 39, -9, -2, 22,
    -- filter=27 channel=17
    -16, 3, -4, -13, 14, 19, -9, 3, 3,
    -- filter=27 channel=18
    -3, 0, -16, -4, 0, 1, 1, -3, -20,
    -- filter=27 channel=19
    3, 9, -8, 10, 15, -4, 7, 0, -6,
    -- filter=27 channel=20
    -10, -5, -11, 10, 3, -19, 2, 6, -2,
    -- filter=27 channel=21
    -1, 2, 10, 13, 7, 6, 0, -2, -1,
    -- filter=27 channel=22
    6, 3, 0, -6, -10, 8, 0, -1, 0,
    -- filter=27 channel=23
    -15, -9, 6, -10, -14, 9, -17, 8, 12,
    -- filter=27 channel=24
    -23, -3, -13, -9, -7, 3, -9, -5, 11,
    -- filter=27 channel=25
    -3, 24, 22, 5, 27, 23, -10, 10, 19,
    -- filter=27 channel=26
    -3, 3, -3, -4, 1, -4, 8, 0, 7,
    -- filter=27 channel=27
    -8, 13, 6, -11, 14, 28, -20, -2, 7,
    -- filter=27 channel=28
    4, -8, 7, 1, 16, 22, -3, 1, 5,
    -- filter=27 channel=29
    0, 11, -11, 27, 34, 30, 12, 20, 1,
    -- filter=27 channel=30
    4, 0, -16, -7, -22, -3, -7, -18, -12,
    -- filter=27 channel=31
    -7, -7, -4, -8, 6, 4, 9, 11, 0,
    -- filter=27 channel=32
    -22, 0, 2, -5, -1, 13, -11, 0, 8,
    -- filter=27 channel=33
    3, 8, 2, 4, 10, 8, 5, 8, 3,
    -- filter=27 channel=34
    5, -2, -7, 0, -4, 2, 11, -4, 5,
    -- filter=27 channel=35
    -6, -3, 4, -14, 10, 20, -17, 2, 12,
    -- filter=27 channel=36
    0, 0, -1, -11, -2, -6, -8, 10, -2,
    -- filter=27 channel=37
    9, 7, -9, 17, 9, 13, 3, 16, -2,
    -- filter=27 channel=38
    -23, 0, 9, -2, 19, 25, -18, 8, 24,
    -- filter=27 channel=39
    -8, 0, 7, 10, 0, -6, 5, 0, -3,
    -- filter=27 channel=40
    5, 3, 14, -3, 5, -2, 3, -2, 0,
    -- filter=27 channel=41
    9, 10, 14, -3, 21, 29, -6, 3, 9,
    -- filter=27 channel=42
    -2, 4, 3, 1, -6, -4, -3, -9, -5,
    -- filter=27 channel=43
    -26, -34, -28, -12, -22, -18, 15, 4, 2,
    -- filter=27 channel=44
    2, 14, 18, -2, 14, 19, -8, 6, 14,
    -- filter=27 channel=45
    6, 4, 0, -1, 8, 0, 0, -4, 0,
    -- filter=27 channel=46
    0, -7, 4, 12, 1, -2, 3, -7, -5,
    -- filter=27 channel=47
    -7, 0, -7, -3, -8, -5, -7, 9, 4,
    -- filter=27 channel=48
    9, 8, 2, 21, 12, 13, -2, 0, 1,
    -- filter=27 channel=49
    0, -4, 0, -1, -1, 8, -11, -20, -12,
    -- filter=27 channel=50
    -4, -17, -4, -12, -10, 0, 1, -13, 5,
    -- filter=27 channel=51
    -19, -15, -16, -6, -17, -2, -6, 6, 7,
    -- filter=27 channel=52
    7, 6, 0, -4, 9, -6, 9, -8, 2,
    -- filter=27 channel=53
    -4, -13, -6, -4, -14, 3, -13, -17, -7,
    -- filter=27 channel=54
    -4, -7, -16, 11, 3, 1, 4, -1, -9,
    -- filter=27 channel=55
    -7, -10, -4, 2, 1, 2, 10, -4, 0,
    -- filter=27 channel=56
    -6, 0, -5, 0, 7, 0, 0, 0, -4,
    -- filter=27 channel=57
    7, -5, -4, 3, -6, 3, 11, -2, -4,
    -- filter=27 channel=58
    7, 3, -2, 3, -7, -5, 11, 6, 9,
    -- filter=27 channel=59
    2, 6, 10, 6, 21, 32, 7, 11, 19,
    -- filter=27 channel=60
    -16, -12, 1, 13, 31, 21, -8, 10, 18,
    -- filter=27 channel=61
    -22, -7, -16, -15, 8, 12, -4, 3, 18,
    -- filter=27 channel=62
    -3, 2, 5, 8, 20, 25, 0, 3, 15,
    -- filter=27 channel=63
    5, 0, 3, 1, -6, 8, 7, 10, 1,
    -- filter=28 channel=0
    1, 8, 7, 3, 9, 7, -3, -8, -7,
    -- filter=28 channel=1
    -1, -3, 8, -9, -3, 0, 6, -9, 4,
    -- filter=28 channel=2
    6, -9, -9, -2, 2, 2, 1, -9, -9,
    -- filter=28 channel=3
    7, 7, 5, -2, 3, -9, -2, -4, -1,
    -- filter=28 channel=4
    -9, 7, 10, 6, -3, 5, 5, 8, 2,
    -- filter=28 channel=5
    0, 0, 7, 6, 7, -1, 7, 0, -3,
    -- filter=28 channel=6
    8, -1, -2, -5, -5, -3, 9, -7, 0,
    -- filter=28 channel=7
    -10, 3, 3, -5, -8, 1, 5, -8, -6,
    -- filter=28 channel=8
    3, -6, 5, 2, -3, 6, 2, 0, 5,
    -- filter=28 channel=9
    -10, -1, 3, -2, -10, -7, 5, 8, -7,
    -- filter=28 channel=10
    5, 7, -4, -3, -3, 1, 0, -10, -5,
    -- filter=28 channel=11
    -10, 0, 8, -7, -1, -2, -6, 0, 4,
    -- filter=28 channel=12
    -1, 0, 1, -9, -5, 8, -3, 8, 0,
    -- filter=28 channel=13
    -8, -4, 2, -1, -8, 3, 2, -7, 6,
    -- filter=28 channel=14
    6, 1, 8, -3, 10, -8, 3, 7, 5,
    -- filter=28 channel=15
    -8, -1, -10, -1, -1, 1, -1, -7, 3,
    -- filter=28 channel=16
    1, -6, -8, -8, 1, 0, -4, 8, -9,
    -- filter=28 channel=17
    -5, 5, 0, -6, 2, 7, 0, -2, -3,
    -- filter=28 channel=18
    -5, -7, 2, -7, -5, 8, -10, 3, -2,
    -- filter=28 channel=19
    0, -8, 10, -10, 9, 1, 4, -5, -6,
    -- filter=28 channel=20
    -3, -1, -6, 5, 3, -9, 2, 2, 1,
    -- filter=28 channel=21
    6, 0, 0, 8, -1, 3, -6, -6, -1,
    -- filter=28 channel=22
    -8, -3, -4, -7, 6, -6, -1, -4, -1,
    -- filter=28 channel=23
    -4, 5, 6, 8, 2, 10, -2, -2, -9,
    -- filter=28 channel=24
    -8, 5, 3, -2, -9, -5, 0, 9, 1,
    -- filter=28 channel=25
    9, -2, 6, -6, -8, -8, 0, -8, -7,
    -- filter=28 channel=26
    0, -3, 4, 0, -3, -1, 3, -1, -4,
    -- filter=28 channel=27
    -4, -2, 9, -5, -7, -6, -7, -7, 0,
    -- filter=28 channel=28
    4, -7, 8, 0, -5, -2, 9, -9, -7,
    -- filter=28 channel=29
    -9, -10, 10, -5, -1, -8, -5, -5, 9,
    -- filter=28 channel=30
    4, -9, 5, 5, -7, 9, 0, -7, -4,
    -- filter=28 channel=31
    3, -8, -6, 8, 8, 3, 9, 5, 3,
    -- filter=28 channel=32
    -4, -3, -1, -10, 0, -9, 0, -3, 0,
    -- filter=28 channel=33
    1, -5, 6, -8, -3, -4, 8, -9, 2,
    -- filter=28 channel=34
    -8, 1, 6, -3, 7, -9, -9, 10, 0,
    -- filter=28 channel=35
    0, -6, 6, 3, -2, 2, 8, 5, 4,
    -- filter=28 channel=36
    3, 8, -4, -5, -9, 0, 4, 0, 0,
    -- filter=28 channel=37
    6, 0, 2, 4, 0, 6, -10, 9, -10,
    -- filter=28 channel=38
    1, -1, -8, 2, 4, -2, -7, 4, 2,
    -- filter=28 channel=39
    -7, -6, -2, 4, 10, -4, 7, -6, -3,
    -- filter=28 channel=40
    -1, -2, -1, -5, 7, 4, -5, 7, -6,
    -- filter=28 channel=41
    2, 0, -9, -3, 0, -4, -3, 8, 0,
    -- filter=28 channel=42
    -1, -7, 0, 8, -3, -8, 3, -8, -7,
    -- filter=28 channel=43
    3, -6, -5, 1, 0, 0, 0, 7, -6,
    -- filter=28 channel=44
    -1, 9, 7, -9, -4, 1, 0, -5, 8,
    -- filter=28 channel=45
    -5, 9, 2, 7, 2, 4, -2, -6, -1,
    -- filter=28 channel=46
    5, 10, 7, -5, 8, 5, 4, -7, 2,
    -- filter=28 channel=47
    5, 8, -3, 7, -1, 1, 6, 7, 1,
    -- filter=28 channel=48
    -10, 3, 0, -2, 0, 0, 0, 6, -1,
    -- filter=28 channel=49
    -3, 3, -8, 7, -6, 7, 0, 2, -5,
    -- filter=28 channel=50
    -2, 1, 5, 9, 7, 0, -5, 3, 9,
    -- filter=28 channel=51
    -7, 5, 0, -8, 2, -2, 7, 5, 4,
    -- filter=28 channel=52
    -10, 1, -5, 5, 10, -10, 8, -4, 5,
    -- filter=28 channel=53
    -8, 4, -4, 7, 4, -7, -9, -10, -1,
    -- filter=28 channel=54
    -7, 9, -8, -1, 2, -5, 3, -7, 9,
    -- filter=28 channel=55
    2, -2, 2, 9, 7, 0, 1, -10, 8,
    -- filter=28 channel=56
    9, 2, 4, 4, 4, -6, -9, -7, 2,
    -- filter=28 channel=57
    -1, -4, -1, -7, -10, -10, -7, 8, 8,
    -- filter=28 channel=58
    6, -4, 7, -4, -2, 3, 2, -2, 0,
    -- filter=28 channel=59
    -5, 1, 9, -10, -3, -2, -5, 7, -3,
    -- filter=28 channel=60
    -2, -5, 5, 10, 4, -8, -2, 10, 8,
    -- filter=28 channel=61
    -7, -4, 8, 6, 9, -3, -1, -7, -8,
    -- filter=28 channel=62
    4, 3, 8, -2, 10, 3, 2, -3, -5,
    -- filter=28 channel=63
    8, 4, -9, 3, -4, 6, 4, -9, 8,
    -- filter=29 channel=0
    6, -15, -1, 9, -14, -12, 7, -10, -17,
    -- filter=29 channel=1
    -9, -13, 0, -11, -12, 0, -9, -7, 0,
    -- filter=29 channel=2
    -3, -1, -21, 4, 0, -15, -8, -5, -16,
    -- filter=29 channel=3
    7, 0, 15, 5, 1, 19, 11, 13, 0,
    -- filter=29 channel=4
    -1, 4, -2, 4, 2, 9, 3, -5, -4,
    -- filter=29 channel=5
    2, 12, 1, 6, 8, 3, 13, 12, -3,
    -- filter=29 channel=6
    -5, 6, -2, -3, 11, -4, -2, -8, -6,
    -- filter=29 channel=7
    10, 1, -7, 6, -3, -8, -1, -9, -7,
    -- filter=29 channel=8
    -2, 5, -4, 8, -2, 1, 0, 0, -10,
    -- filter=29 channel=9
    25, 41, 51, 45, 66, 58, 43, 68, 71,
    -- filter=29 channel=10
    -2, 1, 0, -7, -12, -11, -9, -15, -6,
    -- filter=29 channel=11
    -7, 0, 3, -12, 4, -7, -3, -4, -12,
    -- filter=29 channel=12
    9, 4, 4, 4, 7, 0, -3, 13, 6,
    -- filter=29 channel=13
    0, 14, -3, 11, 20, 2, 0, 4, -2,
    -- filter=29 channel=14
    -1, 5, -9, -9, -4, 4, 8, -1, -11,
    -- filter=29 channel=15
    -8, 6, 0, 5, 11, -8, -3, 2, 2,
    -- filter=29 channel=16
    -15, -2, 0, 10, 5, 5, -2, 10, 2,
    -- filter=29 channel=17
    -8, 9, -5, 5, 4, 8, 10, -9, 1,
    -- filter=29 channel=18
    7, 19, 5, 16, 9, 11, 12, 21, 2,
    -- filter=29 channel=19
    9, 18, 2, 8, 26, 15, 3, 8, 14,
    -- filter=29 channel=20
    2, 15, 17, 11, 24, 9, 0, 19, 19,
    -- filter=29 channel=21
    -4, -2, 0, 6, 0, 11, -1, 11, 12,
    -- filter=29 channel=22
    5, -5, 2, 0, 0, 1, 1, -2, 7,
    -- filter=29 channel=23
    3, -23, 0, -12, -17, -12, -12, -9, -13,
    -- filter=29 channel=24
    -1, 0, 2, 0, 1, -4, 8, 10, -6,
    -- filter=29 channel=25
    -10, -17, -15, -18, -22, -8, -4, -8, -11,
    -- filter=29 channel=26
    0, 0, -17, 4, 8, -10, 0, 0, -16,
    -- filter=29 channel=27
    -9, -2, -12, -3, -14, -12, -11, -12, -22,
    -- filter=29 channel=28
    2, 2, 12, 8, 12, 15, 0, 6, 7,
    -- filter=29 channel=29
    1, 10, 1, 17, 29, 9, -2, 17, 2,
    -- filter=29 channel=30
    0, -21, -19, -12, -3, -21, 0, -19, -22,
    -- filter=29 channel=31
    -1, 0, 0, -5, 7, -5, 11, 10, 0,
    -- filter=29 channel=32
    8, -5, -7, -10, -16, -11, 8, -4, -2,
    -- filter=29 channel=33
    -5, 0, 1, 4, -8, -8, -1, -5, 6,
    -- filter=29 channel=34
    0, -5, -3, 0, -9, -2, -9, 10, -9,
    -- filter=29 channel=35
    -14, -15, -27, -19, -26, -37, -24, -23, -22,
    -- filter=29 channel=36
    14, 12, -3, 4, -3, 0, -5, 10, -3,
    -- filter=29 channel=37
    1, 1, 0, 3, 20, 8, 14, 22, 8,
    -- filter=29 channel=38
    -19, -18, -6, -17, -18, -14, 3, -15, -21,
    -- filter=29 channel=39
    10, 5, 10, -3, -1, 8, 6, 2, 4,
    -- filter=29 channel=40
    -6, 0, -9, 0, -4, -13, 0, 3, -11,
    -- filter=29 channel=41
    -10, 8, -7, 9, 6, -12, 9, -4, -1,
    -- filter=29 channel=42
    -7, 4, -4, 0, 2, 6, 6, 5, 7,
    -- filter=29 channel=43
    -23, -26, -10, -14, -24, -18, -21, -2, -3,
    -- filter=29 channel=44
    0, 1, -10, -6, -13, -16, 1, -12, -14,
    -- filter=29 channel=45
    -2, -3, 9, 0, 0, 1, 8, -6, 9,
    -- filter=29 channel=46
    -8, 0, -6, 5, 3, -3, -4, 10, 4,
    -- filter=29 channel=47
    2, 11, 0, 7, 0, 2, 0, 10, 9,
    -- filter=29 channel=48
    2, 4, -5, 8, 11, 1, 6, 5, 3,
    -- filter=29 channel=49
    8, -7, -11, 5, 3, -4, 6, -9, -11,
    -- filter=29 channel=50
    -4, -4, -9, 9, -2, -2, 5, 0, -1,
    -- filter=29 channel=51
    5, -7, 2, -8, -4, -14, 3, -3, 9,
    -- filter=29 channel=52
    -6, 1, 0, -8, -1, 2, 11, -2, -8,
    -- filter=29 channel=53
    -17, -17, -5, -7, -15, -13, -18, -9, 0,
    -- filter=29 channel=54
    28, 27, 31, 40, 63, 38, 31, 52, 41,
    -- filter=29 channel=55
    10, 1, 3, 4, -1, 0, 4, -2, -1,
    -- filter=29 channel=56
    6, 4, 6, 3, -7, 8, -4, -4, -2,
    -- filter=29 channel=57
    -5, 9, -5, 3, 0, -8, 0, -3, -7,
    -- filter=29 channel=58
    5, 8, 4, 6, 17, 11, 11, 9, 3,
    -- filter=29 channel=59
    -5, 7, -3, -4, -3, -3, 6, -3, 4,
    -- filter=29 channel=60
    -13, -6, -13, 4, -1, -9, -5, -9, -7,
    -- filter=29 channel=61
    -10, -2, 0, -11, -11, -6, 7, 0, 1,
    -- filter=29 channel=62
    0, 13, 13, 12, -2, 11, -7, 11, 6,
    -- filter=29 channel=63
    -7, -7, 7, -9, 0, -8, -7, 0, -4,
    -- filter=30 channel=0
    -2, -4, 5, -6, 2, 13, -8, 7, -5,
    -- filter=30 channel=1
    -8, -6, -6, 4, 10, 11, 4, 11, 18,
    -- filter=30 channel=2
    5, 17, 1, 9, 13, 7, -10, 7, 10,
    -- filter=30 channel=3
    6, 0, -9, 2, 15, -2, 5, 4, -4,
    -- filter=30 channel=4
    -5, -13, 0, -2, 9, 2, -3, -12, -5,
    -- filter=30 channel=5
    -3, -12, -10, -8, 1, 10, -2, -6, -6,
    -- filter=30 channel=6
    3, 4, 2, 8, 10, -5, -10, 2, 3,
    -- filter=30 channel=7
    -7, -5, -5, -13, -6, 2, 3, -5, 4,
    -- filter=30 channel=8
    -21, -16, -15, -4, 1, 16, -13, 8, 1,
    -- filter=30 channel=9
    0, 0, -12, 9, -12, -1, 12, -4, -9,
    -- filter=30 channel=10
    -1, 9, 10, -1, 11, 1, 5, 2, 1,
    -- filter=30 channel=11
    -11, -8, -1, 5, 13, -3, -6, 4, 6,
    -- filter=30 channel=12
    -3, 9, -4, 4, 1, 2, -8, -7, 7,
    -- filter=30 channel=13
    -5, -12, -6, -1, -1, 3, 0, 9, -6,
    -- filter=30 channel=14
    -5, -12, 0, -2, -9, 1, -6, -3, 9,
    -- filter=30 channel=15
    -4, -6, 0, 8, 12, 0, -10, -11, -11,
    -- filter=30 channel=16
    -4, -8, -14, 7, 16, 10, -9, 0, 6,
    -- filter=30 channel=17
    -6, -1, 0, 8, 10, 17, 5, -4, -5,
    -- filter=30 channel=18
    -4, -13, -7, -1, -1, -9, -7, -10, -6,
    -- filter=30 channel=19
    0, 0, 4, -9, 6, -3, -4, 4, 8,
    -- filter=30 channel=20
    -6, -10, -7, -1, -11, -8, 3, -9, -4,
    -- filter=30 channel=21
    -1, 0, 1, -1, 2, -9, -9, -3, 1,
    -- filter=30 channel=22
    -7, 9, -2, -7, -8, -4, 1, 2, 3,
    -- filter=30 channel=23
    -3, -1, 10, 7, 0, 9, 0, 5, -1,
    -- filter=30 channel=24
    -4, -3, 4, -6, -5, -2, 3, 6, 2,
    -- filter=30 channel=25
    15, 23, 3, 17, 32, 19, -2, 20, 16,
    -- filter=30 channel=26
    2, -9, -6, -4, 1, -7, 12, -6, -4,
    -- filter=30 channel=27
    -3, 0, -6, 13, 29, 16, -5, 21, 4,
    -- filter=30 channel=28
    -6, -12, -8, -1, 0, 9, 3, -4, -7,
    -- filter=30 channel=29
    -9, -17, -22, 6, 9, 6, 0, -8, -9,
    -- filter=30 channel=30
    2, -17, -3, 1, -1, -10, -7, -4, -7,
    -- filter=30 channel=31
    0, 7, 8, 0, -2, -2, -7, 6, 3,
    -- filter=30 channel=32
    6, 5, 3, -1, 13, 5, 8, 4, 1,
    -- filter=30 channel=33
    -3, 0, -1, -4, 9, -6, -4, -7, 5,
    -- filter=30 channel=34
    -5, 1, 0, 2, 1, -1, 0, 5, -3,
    -- filter=30 channel=35
    11, 13, 17, 16, 13, 22, -1, 19, 7,
    -- filter=30 channel=36
    7, 10, 8, 5, 3, -4, 7, 8, 0,
    -- filter=30 channel=37
    2, -7, -11, 4, 4, -1, 12, 9, 0,
    -- filter=30 channel=38
    0, -8, -2, -6, 6, 16, 9, 5, 20,
    -- filter=30 channel=39
    -7, 0, 8, 2, 8, 6, 0, 0, 3,
    -- filter=30 channel=40
    -2, 6, 9, 11, 0, 8, -6, -2, 8,
    -- filter=30 channel=41
    -8, -3, -3, 10, 17, 26, 7, 1, 10,
    -- filter=30 channel=42
    9, 9, 7, -5, 3, 5, -4, -7, -2,
    -- filter=30 channel=43
    -11, -13, 0, -3, -5, 0, 8, 19, 15,
    -- filter=30 channel=44
    14, 4, 4, 10, -2, 3, 7, 1, -1,
    -- filter=30 channel=45
    6, -2, -1, 4, 3, -2, 8, 10, 0,
    -- filter=30 channel=46
    -4, 1, -1, 9, -10, -11, -5, -8, 0,
    -- filter=30 channel=47
    10, -6, -3, -9, -2, 7, -8, -2, 5,
    -- filter=30 channel=48
    7, -12, 1, 14, 9, 6, 1, 3, 0,
    -- filter=30 channel=49
    4, 14, 14, -2, 11, 16, -18, -7, 4,
    -- filter=30 channel=50
    -15, -12, -7, -12, -20, 1, -7, -7, -11,
    -- filter=30 channel=51
    2, -1, -4, 3, -4, 9, -10, -4, -5,
    -- filter=30 channel=52
    4, 6, 2, 7, 5, -1, -9, -6, -5,
    -- filter=30 channel=53
    -10, 6, 4, -4, -13, 1, -2, -2, -5,
    -- filter=30 channel=54
    6, 6, -9, -2, -1, 3, 2, -9, 3,
    -- filter=30 channel=55
    8, -6, 6, -1, -8, 4, 4, -7, 3,
    -- filter=30 channel=56
    7, 0, -3, -5, 0, -4, 7, -3, -5,
    -- filter=30 channel=57
    -9, 10, 8, -1, 8, -4, 10, -6, 6,
    -- filter=30 channel=58
    9, 1, 8, 9, -2, -12, -3, -5, -7,
    -- filter=30 channel=59
    -8, 2, 6, 9, 5, 7, -3, 14, 3,
    -- filter=30 channel=60
    -19, -8, -8, 9, 17, 15, 4, 2, 1,
    -- filter=30 channel=61
    -13, -10, -10, 3, 14, 16, -12, -2, 8,
    -- filter=30 channel=62
    -2, -1, -10, -3, 5, -4, -7, 3, 4,
    -- filter=30 channel=63
    0, -2, 0, -1, 8, 0, -7, -1, 3,
    -- filter=31 channel=0
    -4, 19, 11, 3, 16, 25, 1, 16, 24,
    -- filter=31 channel=1
    0, -23, -7, -21, -13, -24, -17, -23, -11,
    -- filter=31 channel=2
    5, -19, -12, -15, -25, -17, -29, -24, -17,
    -- filter=31 channel=3
    -12, -6, 3, -5, -11, -2, -27, -20, -5,
    -- filter=31 channel=4
    3, 10, 15, 15, 26, 15, -1, 10, 4,
    -- filter=31 channel=5
    -9, -8, 0, -9, -9, -12, -2, -6, -6,
    -- filter=31 channel=6
    5, 1, 0, -10, 10, 0, 0, -4, -8,
    -- filter=31 channel=7
    -7, -5, -5, -14, -1, -2, -4, -3, 5,
    -- filter=31 channel=8
    -6, 23, 17, 3, 34, 38, -18, -2, 19,
    -- filter=31 channel=9
    -2, -25, -18, -14, -18, -30, -17, -17, -30,
    -- filter=31 channel=10
    2, 9, 4, -1, 14, 1, 15, 17, 10,
    -- filter=31 channel=11
    -12, 9, 19, 10, 1, 23, 0, -6, 3,
    -- filter=31 channel=12
    10, -6, -4, 5, -7, -7, 6, -6, 0,
    -- filter=31 channel=13
    0, 21, 18, 17, 27, 19, 12, 26, 12,
    -- filter=31 channel=14
    -16, -11, 0, -14, 1, -6, -4, -2, -10,
    -- filter=31 channel=15
    2, 23, 9, 5, 23, 26, -8, 17, 18,
    -- filter=31 channel=16
    -6, 0, 0, 9, 3, 12, -11, -11, 2,
    -- filter=31 channel=17
    8, 7, 17, 2, 22, 23, 1, 9, 13,
    -- filter=31 channel=18
    12, 26, 22, 17, 33, 37, 13, 34, 12,
    -- filter=31 channel=19
    -17, -11, -21, -21, -20, -28, -17, -19, -26,
    -- filter=31 channel=20
    -2, -2, -16, -6, -23, -11, -3, -6, 0,
    -- filter=31 channel=21
    2, 8, -5, 9, 8, -7, 6, -6, 8,
    -- filter=31 channel=22
    -8, -9, 4, -9, -5, -2, -10, -3, 0,
    -- filter=31 channel=23
    -1, 7, 6, 5, 0, 4, 5, 0, 11,
    -- filter=31 channel=24
    0, 3, 11, 0, 23, 26, -3, 14, 24,
    -- filter=31 channel=25
    -15, -28, -28, -25, -22, -21, -32, -36, -36,
    -- filter=31 channel=26
    -16, -8, -11, -17, -9, -4, -9, -4, -17,
    -- filter=31 channel=27
    -4, 1, 2, 0, -5, -2, -19, -18, -14,
    -- filter=31 channel=28
    0, 10, 12, 0, 1, 20, -12, -1, -5,
    -- filter=31 channel=29
    3, 16, 4, 7, 7, 17, -5, -5, 13,
    -- filter=31 channel=30
    -37, -32, -8, -34, -34, -30, -44, -48, -21,
    -- filter=31 channel=31
    -6, -6, 0, 4, 6, -11, 2, -1, 0,
    -- filter=31 channel=32
    -25, -14, -27, -19, -31, -18, -10, -12, -14,
    -- filter=31 channel=33
    -5, -7, -3, 5, -7, 9, 7, 6, -5,
    -- filter=31 channel=34
    -2, -11, -3, -12, -9, -3, -12, -7, 1,
    -- filter=31 channel=35
    -11, -9, -2, -3, -9, 6, -15, -14, -14,
    -- filter=31 channel=36
    3, -4, 4, -3, 2, -6, 7, 9, -7,
    -- filter=31 channel=37
    -6, -8, -14, -9, -22, -17, -9, -24, -1,
    -- filter=31 channel=38
    -12, 2, 3, -14, -3, -1, -16, 2, 6,
    -- filter=31 channel=39
    -9, -4, 9, 1, -9, 7, 0, 3, 6,
    -- filter=31 channel=40
    -14, 3, 3, -2, -14, 1, -11, 3, -16,
    -- filter=31 channel=41
    3, 5, 22, 9, 16, 20, -24, -7, 10,
    -- filter=31 channel=42
    6, 6, -5, 0, -10, -4, -5, -3, 0,
    -- filter=31 channel=43
    -22, -19, -15, -12, -22, -16, -14, -10, -4,
    -- filter=31 channel=44
    -24, -21, -17, -27, -33, -27, -27, -31, -30,
    -- filter=31 channel=45
    -5, 0, 1, -7, -10, 3, -5, -5, -3,
    -- filter=31 channel=46
    1, -10, -12, 0, -3, -4, -16, -2, -14,
    -- filter=31 channel=47
    8, -7, 3, -7, -3, -3, 0, -3, -2,
    -- filter=31 channel=48
    4, 11, 6, 0, 0, 3, -9, 0, -1,
    -- filter=31 channel=49
    11, 8, 12, 0, 14, 31, 1, 2, 12,
    -- filter=31 channel=50
    -10, -19, -20, -16, -17, -20, -2, -11, -11,
    -- filter=31 channel=51
    15, 11, 17, 7, 30, 20, 18, 31, 22,
    -- filter=31 channel=52
    11, 8, -5, 9, 3, 0, 11, 4, -1,
    -- filter=31 channel=53
    -25, -28, -15, -32, -41, -20, -33, -34, -24,
    -- filter=31 channel=54
    -14, -10, -11, -18, -28, -18, -19, -32, -23,
    -- filter=31 channel=55
    7, -4, 9, -1, 4, 4, 0, -7, -7,
    -- filter=31 channel=56
    3, -6, -12, -4, -11, 6, 0, 3, 9,
    -- filter=31 channel=57
    4, 3, 6, 0, 9, -9, -2, -1, -2,
    -- filter=31 channel=58
    7, -1, 6, -8, 2, 3, 2, 8, 4,
    -- filter=31 channel=59
    -12, -8, 0, -8, -2, -8, -28, -10, -7,
    -- filter=31 channel=60
    9, 31, 16, 12, 43, 35, -6, 24, 28,
    -- filter=31 channel=61
    2, 19, 32, 7, 26, 24, -6, 18, 21,
    -- filter=31 channel=62
    -15, -4, -3, -9, -5, 0, -16, -13, -12,
    -- filter=31 channel=63
    -1, -2, -3, 1, 2, -6, 5, 8, -4,
    -- filter=32 channel=0
    -14, -15, -2, 8, 5, -9, -6, 0, 6,
    -- filter=32 channel=1
    -3, 6, -4, -10, 23, 14, -10, 21, 15,
    -- filter=32 channel=2
    -17, 1, -3, -12, 19, 12, -24, 4, -10,
    -- filter=32 channel=3
    20, 16, 2, 18, 31, 11, 20, 29, 3,
    -- filter=32 channel=4
    -7, -1, -10, 6, 0, 5, -10, 1, 3,
    -- filter=32 channel=5
    -2, 11, 14, -2, 21, 1, -1, 9, 0,
    -- filter=32 channel=6
    0, 5, -6, 1, -5, 6, -4, 2, -12,
    -- filter=32 channel=7
    1, 10, -1, 2, 0, -7, -5, 9, -4,
    -- filter=32 channel=8
    -4, -7, -3, -2, 21, -5, -19, 5, -5,
    -- filter=32 channel=9
    2, 26, 13, 10, 17, 16, 14, 21, 13,
    -- filter=32 channel=10
    -18, -7, 1, -8, -11, 6, -3, -6, 11,
    -- filter=32 channel=11
    -6, -8, 3, -10, 15, 4, 2, 7, -3,
    -- filter=32 channel=12
    11, 1, 0, 10, 2, 0, 8, 7, 0,
    -- filter=32 channel=13
    -8, -14, -4, 0, 7, -8, 0, 4, 2,
    -- filter=32 channel=14
    2, 3, -3, -2, 12, 9, 3, -3, -8,
    -- filter=32 channel=15
    1, 6, -21, 1, 12, -6, -14, -11, -15,
    -- filter=32 channel=16
    -8, 14, 2, -3, 29, 7, -1, -7, -9,
    -- filter=32 channel=17
    5, 7, -6, -5, 9, 14, -2, -4, -7,
    -- filter=32 channel=18
    7, -11, -3, -5, 4, -3, 5, -3, -18,
    -- filter=32 channel=19
    10, 8, -7, 4, 17, 5, -8, 5, 1,
    -- filter=32 channel=20
    5, 15, 10, 7, 19, 0, -2, 9, -4,
    -- filter=32 channel=21
    -3, -6, -5, 0, -6, -8, 0, -10, 4,
    -- filter=32 channel=22
    -10, 9, 7, 6, 3, 4, 7, 8, -2,
    -- filter=32 channel=23
    -10, -1, 8, -6, -8, 7, 2, 10, -1,
    -- filter=32 channel=24
    -9, 0, -15, -12, 5, -7, 4, -5, -6,
    -- filter=32 channel=25
    -3, 22, 6, -12, 23, 8, -3, 11, 10,
    -- filter=32 channel=26
    13, 5, 9, 7, 8, 7, 0, 11, 7,
    -- filter=32 channel=27
    -3, 6, 0, 0, 9, 8, -16, 0, 8,
    -- filter=32 channel=28
    -9, 14, -2, -9, 8, -5, -21, -7, -16,
    -- filter=32 channel=29
    7, -5, -23, 19, 31, -8, 0, 8, -6,
    -- filter=32 channel=30
    -2, 22, 11, 8, 16, -1, -5, 6, 7,
    -- filter=32 channel=31
    0, 0, 1, 10, -10, 5, -8, -6, -4,
    -- filter=32 channel=32
    0, -4, 2, 2, -2, 21, -12, 14, 22,
    -- filter=32 channel=33
    -9, -4, -9, -3, 8, -7, -1, -6, -1,
    -- filter=32 channel=34
    9, 5, -7, 13, 10, -10, 9, 0, -7,
    -- filter=32 channel=35
    -7, -2, -1, -16, 16, 7, -10, 4, -1,
    -- filter=32 channel=36
    3, -2, 6, -7, -7, 6, 4, 9, 3,
    -- filter=32 channel=37
    18, 9, -5, 22, 26, 10, 12, 20, -1,
    -- filter=32 channel=38
    -2, 9, 0, 4, 8, 11, -17, 16, 7,
    -- filter=32 channel=39
    6, 9, -9, -5, 5, 11, -8, -9, -9,
    -- filter=32 channel=40
    2, 12, -4, 1, 2, 7, 7, -4, 0,
    -- filter=32 channel=41
    -3, 8, 5, 8, 22, 3, 0, 9, -12,
    -- filter=32 channel=42
    -6, 8, 8, 7, 9, 6, 4, -2, -3,
    -- filter=32 channel=43
    -4, -7, -4, 13, 5, 1, 14, 15, 19,
    -- filter=32 channel=44
    9, 20, 23, -8, 9, 22, 7, 0, 12,
    -- filter=32 channel=45
    7, -5, 1, 0, 10, -2, 6, -9, -1,
    -- filter=32 channel=46
    -1, 10, -8, 4, 15, 6, 12, 0, -9,
    -- filter=32 channel=47
    3, -6, -8, -9, 6, -7, 3, -3, 0,
    -- filter=32 channel=48
    4, 0, 2, 1, 18, 0, 5, 0, -13,
    -- filter=32 channel=49
    -5, 7, 8, -15, -6, 8, -18, -8, -15,
    -- filter=32 channel=50
    3, 3, 4, 4, 5, 4, -4, 0, 2,
    -- filter=32 channel=51
    -2, -20, -2, -4, -3, -5, -5, -14, 8,
    -- filter=32 channel=52
    -3, 8, 1, 5, -6, 3, -5, 0, -5,
    -- filter=32 channel=53
    -8, 17, 9, -2, 20, 14, -2, 17, 3,
    -- filter=32 channel=54
    6, 26, 14, 16, 22, 6, 12, 12, 5,
    -- filter=32 channel=55
    10, -3, -7, -6, -6, 0, 2, -5, -6,
    -- filter=32 channel=56
    -1, -2, -3, -3, 9, 5, 11, -6, -3,
    -- filter=32 channel=57
    -5, 0, -10, -5, -2, -1, 0, 11, -9,
    -- filter=32 channel=58
    -6, 1, 1, 12, 5, -11, 1, -6, -6,
    -- filter=32 channel=59
    16, 18, 14, 6, 28, 4, 11, 21, 0,
    -- filter=32 channel=60
    8, 10, -15, 4, 9, 8, 4, 12, -6,
    -- filter=32 channel=61
    -9, 0, -17, -10, 11, -5, 0, 10, 5,
    -- filter=32 channel=62
    15, 14, 15, 17, 23, 5, -3, 19, -1,
    -- filter=32 channel=63
    8, -4, 1, -4, 6, -6, 6, -9, -9,
    -- filter=33 channel=0
    -3, 9, -4, 7, 9, 4, 4, 5, -7,
    -- filter=33 channel=1
    -8, 5, 18, -4, 24, 20, -4, 17, 10,
    -- filter=33 channel=2
    16, 16, 8, -2, 8, 10, -8, 3, 0,
    -- filter=33 channel=3
    21, 10, 2, 13, 10, -2, 3, 7, 11,
    -- filter=33 channel=4
    8, -3, -7, -8, -8, 3, -18, -6, -16,
    -- filter=33 channel=5
    3, 0, -4, 9, 7, 1, 2, 1, 2,
    -- filter=33 channel=6
    -3, 4, 0, -9, -6, -8, -7, -10, 5,
    -- filter=33 channel=7
    9, -6, -9, -8, -7, -7, -9, -8, -3,
    -- filter=33 channel=8
    10, 25, 9, 2, 4, -5, -25, -6, -17,
    -- filter=33 channel=9
    -3, 4, -10, 9, 2, -11, 0, 3, -13,
    -- filter=33 channel=10
    -10, -1, 0, 3, 8, -5, 8, 3, 5,
    -- filter=33 channel=11
    7, 2, 10, 2, 10, 11, -13, -10, -13,
    -- filter=33 channel=12
    5, -2, -9, -5, 10, -2, 0, -1, -3,
    -- filter=33 channel=13
    3, 10, 1, -1, 8, 9, 4, -6, -16,
    -- filter=33 channel=14
    -11, -4, 9, -7, 7, -5, 1, 1, 6,
    -- filter=33 channel=15
    20, 21, 9, 0, 3, -8, -25, -15, -5,
    -- filter=33 channel=16
    25, 27, 22, 11, 13, 2, -8, -2, -13,
    -- filter=33 channel=17
    -2, 13, 14, -3, 5, 6, -4, -11, -16,
    -- filter=33 channel=18
    -3, -3, -15, -9, -9, -3, -1, 0, -13,
    -- filter=33 channel=19
    -8, 7, 7, 0, 11, 15, -8, 2, 6,
    -- filter=33 channel=20
    -7, 5, -12, 2, 0, 3, 0, 7, -2,
    -- filter=33 channel=21
    6, -5, -5, 1, 4, 0, 9, 0, -2,
    -- filter=33 channel=22
    6, -8, -3, -3, -1, 8, 8, -7, 9,
    -- filter=33 channel=23
    -16, -10, -2, -11, 0, -3, 1, 3, 1,
    -- filter=33 channel=24
    -12, -2, 9, -10, 14, 13, -7, -11, -16,
    -- filter=33 channel=25
    16, 27, 11, -3, 12, 19, -8, 8, 15,
    -- filter=33 channel=26
    11, 3, -12, -2, -4, -7, 6, 13, 7,
    -- filter=33 channel=27
    10, 30, 21, -14, 5, 0, -12, 1, 9,
    -- filter=33 channel=28
    1, 1, 12, -9, 1, 6, -21, -6, -13,
    -- filter=33 channel=29
    22, 33, 1, 14, 18, -2, -17, -15, -17,
    -- filter=33 channel=30
    0, 3, -2, 0, 9, 9, -8, -3, 8,
    -- filter=33 channel=31
    -2, -1, -6, 10, -7, 0, 0, 0, 3,
    -- filter=33 channel=32
    0, 5, -4, -9, 6, -1, -4, 8, 5,
    -- filter=33 channel=33
    -8, -7, 5, 2, 6, 0, -2, -6, 1,
    -- filter=33 channel=34
    2, 6, 5, 7, -3, 4, -7, -8, 5,
    -- filter=33 channel=35
    8, 21, 0, 0, 0, 4, -17, 9, 9,
    -- filter=33 channel=36
    -4, -7, -11, -2, 2, 8, 7, 2, 1,
    -- filter=33 channel=37
    8, 5, 2, 14, 15, 6, 5, 0, 3,
    -- filter=33 channel=38
    -1, 9, 4, 0, 23, 1, -16, -8, -11,
    -- filter=33 channel=39
    10, -8, -6, -6, 5, -3, 10, 1, -1,
    -- filter=33 channel=40
    10, 0, 9, -6, 0, 8, 7, -8, 3,
    -- filter=33 channel=41
    8, 29, 22, 5, 3, 0, -6, -8, -4,
    -- filter=33 channel=42
    -5, 2, 9, 9, 3, 8, -8, 8, -8,
    -- filter=33 channel=43
    -9, 2, 0, 9, 8, 17, -7, 3, 1,
    -- filter=33 channel=44
    2, -3, 3, -1, 8, -2, -3, -2, 9,
    -- filter=33 channel=45
    -2, 7, -7, -9, 4, -7, 10, -5, 8,
    -- filter=33 channel=46
    1, 6, 0, 1, -6, -8, -5, -6, -10,
    -- filter=33 channel=47
    8, 3, 0, 1, 6, -2, -10, 6, -4,
    -- filter=33 channel=48
    10, 2, 2, -3, 4, 8, -3, 5, -4,
    -- filter=33 channel=49
    -1, -6, 0, -13, 1, -4, -15, -8, 0,
    -- filter=33 channel=50
    -7, -5, -5, 0, -2, -2, -6, -8, -2,
    -- filter=33 channel=51
    2, -15, -7, -11, 4, 4, -4, -9, 2,
    -- filter=33 channel=52
    -1, 1, -2, 9, 5, -3, 4, 5, -8,
    -- filter=33 channel=53
    -15, -7, 13, -5, 5, -2, -15, -6, -7,
    -- filter=33 channel=54
    -9, 0, -13, -4, -8, -1, -15, 1, -4,
    -- filter=33 channel=55
    -10, -2, 7, -6, -9, 1, -5, -6, -9,
    -- filter=33 channel=56
    5, -10, 0, -10, 10, 6, 8, 1, 3,
    -- filter=33 channel=57
    -9, 1, 6, 5, -9, 0, 4, 8, 10,
    -- filter=33 channel=58
    -1, 0, 5, -4, 0, 0, 9, 4, 1,
    -- filter=33 channel=59
    17, 25, 25, 4, 15, 1, -11, 5, -5,
    -- filter=33 channel=60
    28, 28, -3, 6, 4, 5, -26, -17, -12,
    -- filter=33 channel=61
    8, 16, 13, 4, 16, 1, -12, -19, -14,
    -- filter=33 channel=62
    9, 21, 15, 11, 18, 2, -7, 1, -5,
    -- filter=33 channel=63
    -2, -5, 2, -9, -6, 1, 6, -10, 0,
    -- filter=34 channel=0
    -5, 10, 2, -11, 20, 9, -13, 4, 20,
    -- filter=34 channel=1
    2, -19, 4, -15, -19, 10, -8, -14, 15,
    -- filter=34 channel=2
    -15, -9, 20, -17, -1, 16, -19, -10, -3,
    -- filter=34 channel=3
    -15, 12, 15, -11, 16, 23, -9, -6, 19,
    -- filter=34 channel=4
    -10, 7, 11, -10, -11, 17, -1, -8, 16,
    -- filter=34 channel=5
    9, -5, 6, 22, -10, 11, 10, 1, 17,
    -- filter=34 channel=6
    -14, 5, -5, -9, 0, 6, -11, 0, -7,
    -- filter=34 channel=7
    15, 0, 8, 10, 13, 21, 27, 19, 16,
    -- filter=34 channel=8
    -16, 2, 28, -15, -9, 45, -14, -17, 10,
    -- filter=34 channel=9
    -4, -5, 7, 2, -8, -1, -1, 1, 0,
    -- filter=34 channel=10
    -12, -8, 7, -16, 5, -4, -19, 4, -1,
    -- filter=34 channel=11
    -3, -13, 5, -8, -5, 26, -7, -7, 15,
    -- filter=34 channel=12
    8, 6, -2, -7, 6, 3, 5, -7, 8,
    -- filter=34 channel=13
    -13, 15, 10, -10, 16, 18, -23, -6, 20,
    -- filter=34 channel=14
    9, 7, 7, 16, 6, 23, 17, 0, 11,
    -- filter=34 channel=15
    -26, 5, 12, -38, 1, 33, -15, -3, 16,
    -- filter=34 channel=16
    -14, -14, 19, -21, -14, 26, -22, -18, 9,
    -- filter=34 channel=17
    -12, -4, 17, 6, -24, 36, 1, -12, 3,
    -- filter=34 channel=18
    -2, 1, -6, -5, 13, 5, -8, 11, -4,
    -- filter=34 channel=19
    0, -9, 3, 15, -31, 19, 24, -18, 15,
    -- filter=34 channel=20
    -6, 24, 12, 5, 25, 15, -10, 22, 13,
    -- filter=34 channel=21
    2, 7, 0, -3, 4, -7, -3, 0, -3,
    -- filter=34 channel=22
    -9, 2, 0, 8, 9, -10, 0, -8, 1,
    -- filter=34 channel=23
    -9, -8, 4, -16, -7, 0, 1, -15, 7,
    -- filter=34 channel=24
    9, -17, 12, 0, -20, 14, -6, -3, 5,
    -- filter=34 channel=25
    -17, -6, 18, -26, 3, 14, -21, -16, 11,
    -- filter=34 channel=26
    4, 25, 10, -2, 37, 24, 8, 16, 29,
    -- filter=34 channel=27
    -12, 0, 20, -34, -19, 31, -11, -16, 11,
    -- filter=34 channel=28
    2, -17, 0, -7, -17, 28, 2, -12, 1,
    -- filter=34 channel=29
    -23, 0, 23, -37, 13, 28, -33, -2, 20,
    -- filter=34 channel=30
    48, 31, 41, 66, 15, 58, 47, 31, 47,
    -- filter=34 channel=31
    4, 8, -6, -10, 7, 0, -3, 3, 0,
    -- filter=34 channel=32
    7, -3, 5, 6, -16, 12, 6, -8, 10,
    -- filter=34 channel=33
    6, -2, -10, -9, 8, 8, 7, -10, -3,
    -- filter=34 channel=34
    14, 2, 2, 11, 14, 6, 14, 7, 10,
    -- filter=34 channel=35
    -12, -7, 11, -25, 3, 18, -25, -11, 1,
    -- filter=34 channel=36
    3, -2, -1, 10, 9, 0, 5, -7, 6,
    -- filter=34 channel=37
    8, 4, 2, 5, -14, 16, -1, -11, 16,
    -- filter=34 channel=38
    -26, -3, 19, -34, -3, 32, -17, -20, 26,
    -- filter=34 channel=39
    0, -6, -9, 8, -10, 4, -10, -3, 7,
    -- filter=34 channel=40
    -2, -4, 2, -4, 8, 7, 8, -10, 2,
    -- filter=34 channel=41
    -15, 3, 35, -35, -5, 37, -13, -19, 15,
    -- filter=34 channel=42
    0, 0, -3, -2, -8, 3, -8, 3, -5,
    -- filter=34 channel=43
    18, 4, -17, -2, 3, 3, -16, -6, -2,
    -- filter=34 channel=44
    3, 1, 21, 21, 0, 7, 25, -5, 1,
    -- filter=34 channel=45
    0, 5, -4, -5, 0, -3, 4, -9, -9,
    -- filter=34 channel=46
    4, 10, 20, 2, 34, 26, 9, 14, 17,
    -- filter=34 channel=47
    3, -7, 8, 9, -4, -5, 3, 9, -7,
    -- filter=34 channel=48
    -19, 19, 5, -14, 25, 5, -4, 4, 16,
    -- filter=34 channel=49
    -4, 7, 6, -13, -6, 21, 8, -14, -1,
    -- filter=34 channel=50
    38, 1, 8, 28, -2, 22, 29, 0, 22,
    -- filter=34 channel=51
    5, 6, 7, -10, 12, 2, 2, 6, 6,
    -- filter=34 channel=52
    -7, 10, -7, 6, 7, -6, 3, -1, -1,
    -- filter=34 channel=53
    21, 23, 36, 42, 4, 39, 39, 8, 36,
    -- filter=34 channel=54
    14, 1, 12, 0, -11, 7, 0, -17, 2,
    -- filter=34 channel=55
    7, 0, -7, 3, 4, 8, 8, 8, -5,
    -- filter=34 channel=56
    16, 11, -4, 20, 8, 13, 8, 0, 3,
    -- filter=34 channel=57
    1, 5, 3, 2, 9, 2, 6, 2, 7,
    -- filter=34 channel=58
    3, -2, -4, -3, 2, -14, 2, 9, -3,
    -- filter=34 channel=59
    -12, 5, 2, -32, 16, 25, -13, 5, 2,
    -- filter=34 channel=60
    -20, -3, 34, -46, 15, 61, -31, -6, 40,
    -- filter=34 channel=61
    -12, -6, 16, -14, -8, 42, -5, -16, 30,
    -- filter=34 channel=62
    -9, -13, 4, 5, -7, 18, -6, -8, 5,
    -- filter=34 channel=63
    9, 0, -7, 1, 6, -7, -3, -8, 4,
    -- filter=35 channel=0
    -2, -8, -10, -9, -9, 0, 4, -8, 0,
    -- filter=35 channel=1
    9, -8, 7, -9, 8, 2, 9, 9, 1,
    -- filter=35 channel=2
    1, 4, 0, 9, -8, -5, 0, -2, -8,
    -- filter=35 channel=3
    -3, 9, -3, -9, 6, 3, -3, 8, -8,
    -- filter=35 channel=4
    -8, 2, 0, 9, 3, 3, 1, 2, 5,
    -- filter=35 channel=5
    7, -6, 0, -4, 0, -10, -6, 9, -9,
    -- filter=35 channel=6
    8, 10, -3, -1, -3, -10, 2, -2, -8,
    -- filter=35 channel=7
    10, 7, 4, -3, -8, -4, -5, 7, 3,
    -- filter=35 channel=8
    8, 2, 9, -3, -1, -1, -6, -2, 9,
    -- filter=35 channel=9
    10, -5, -5, 7, 6, -6, 4, -3, -9,
    -- filter=35 channel=10
    -8, -2, -8, -8, 6, 10, -1, -5, 1,
    -- filter=35 channel=11
    2, 8, -9, 9, 7, -4, -8, -5, 3,
    -- filter=35 channel=12
    -8, -2, 8, 3, 1, -1, 9, -6, 9,
    -- filter=35 channel=13
    2, -5, 7, 8, 3, -2, 8, -1, -9,
    -- filter=35 channel=14
    7, 0, -9, 6, 7, 9, -5, -1, 1,
    -- filter=35 channel=15
    -8, -10, 2, 0, 0, -4, -4, -4, 10,
    -- filter=35 channel=16
    -7, -5, 7, -9, -8, 2, -2, 4, 8,
    -- filter=35 channel=17
    0, -3, 5, 0, 9, -2, 9, 6, 8,
    -- filter=35 channel=18
    -8, 7, -4, 7, -8, 5, 10, -2, 0,
    -- filter=35 channel=19
    1, -6, -2, 6, 9, 10, 2, -1, -7,
    -- filter=35 channel=20
    -4, -7, -10, -10, -2, -3, 4, 6, -7,
    -- filter=35 channel=21
    8, 10, 6, 0, 2, -6, -7, 1, 10,
    -- filter=35 channel=22
    -3, 0, -1, 9, -3, 1, 2, 4, -6,
    -- filter=35 channel=23
    3, 8, -6, 0, 8, -2, -10, -4, -7,
    -- filter=35 channel=24
    5, 1, 3, -3, -10, -6, 7, 9, 0,
    -- filter=35 channel=25
    -1, 1, -3, -2, 5, -2, 7, -2, -4,
    -- filter=35 channel=26
    3, 9, 8, 0, -5, 6, -4, 4, -5,
    -- filter=35 channel=27
    -4, 1, -10, 2, -2, -10, -3, -4, 6,
    -- filter=35 channel=28
    7, 6, -7, 0, 0, -9, 2, 5, 6,
    -- filter=35 channel=29
    8, -7, -2, -2, -7, -3, -3, 7, 2,
    -- filter=35 channel=30
    0, -6, 10, 0, -10, -10, -3, 9, -2,
    -- filter=35 channel=31
    5, 7, 3, -10, -7, 1, 10, 7, 10,
    -- filter=35 channel=32
    0, 4, -7, -6, 7, 1, 9, 0, 4,
    -- filter=35 channel=33
    0, -4, -9, 7, -4, 9, -6, 6, -6,
    -- filter=35 channel=34
    6, -9, 8, 6, 8, 4, -4, 0, 9,
    -- filter=35 channel=35
    -1, -2, -6, 9, -7, 1, -3, -4, 1,
    -- filter=35 channel=36
    5, 9, 1, 5, 0, -8, 9, -9, -4,
    -- filter=35 channel=37
    -9, 0, -9, -6, -10, 1, 8, 1, -6,
    -- filter=35 channel=38
    10, -8, -10, 4, -8, 5, -6, 5, 0,
    -- filter=35 channel=39
    -8, -5, 10, 1, 0, 4, 0, -10, -7,
    -- filter=35 channel=40
    0, 1, -2, 2, 0, -2, -4, -8, 0,
    -- filter=35 channel=41
    -9, -1, 1, -7, 7, -6, -7, -6, -5,
    -- filter=35 channel=42
    -3, -10, 9, -3, -6, 3, -8, 4, -3,
    -- filter=35 channel=43
    6, 4, -7, 2, 6, 6, 1, 3, 10,
    -- filter=35 channel=44
    -8, 0, 5, -8, -4, -3, 8, -3, -7,
    -- filter=35 channel=45
    -3, 1, -7, 0, -1, -4, 7, 0, 7,
    -- filter=35 channel=46
    2, -4, -7, 2, 7, -5, -8, 0, 4,
    -- filter=35 channel=47
    3, 9, 8, 7, 8, -6, -6, 4, -1,
    -- filter=35 channel=48
    -9, -6, 5, -4, 0, 0, -10, 1, -7,
    -- filter=35 channel=49
    -7, -4, -9, -9, -3, -2, -6, 10, -3,
    -- filter=35 channel=50
    4, 0, 3, 9, -8, -7, -2, -4, 8,
    -- filter=35 channel=51
    -4, 0, -1, -4, 0, 2, 6, -2, 4,
    -- filter=35 channel=52
    6, -1, 0, -1, 3, -1, 4, 2, 8,
    -- filter=35 channel=53
    7, 4, 4, 3, -2, -3, 0, -9, 4,
    -- filter=35 channel=54
    -8, 7, 1, -4, 10, -5, -5, -4, 5,
    -- filter=35 channel=55
    -10, 4, 3, -10, -7, 0, 3, -5, 5,
    -- filter=35 channel=56
    8, -3, -3, -7, -3, 7, 5, 1, -7,
    -- filter=35 channel=57
    9, -5, -3, -6, -4, 3, -5, 5, -5,
    -- filter=35 channel=58
    -3, 4, -9, 1, -2, 0, -8, 3, 8,
    -- filter=35 channel=59
    1, -3, -7, -2, -9, -9, 6, -6, -3,
    -- filter=35 channel=60
    -10, 5, -10, 3, -2, -6, 0, 7, 8,
    -- filter=35 channel=61
    0, -4, 4, 9, 4, -6, 9, -1, -2,
    -- filter=35 channel=62
    5, 5, 8, -9, -9, -6, -5, -9, -10,
    -- filter=35 channel=63
    -4, 0, 9, 10, -8, 2, -4, -6, 0,
    -- filter=36 channel=0
    4, 4, -7, 2, -1, 0, 10, 1, 0,
    -- filter=36 channel=1
    -5, -8, -9, -8, -18, -7, -13, -12, -19,
    -- filter=36 channel=2
    -7, -5, -13, -7, -13, -14, 3, -10, -14,
    -- filter=36 channel=3
    -12, -4, -19, -2, -11, -8, -3, -15, -8,
    -- filter=36 channel=4
    13, 3, 12, 1, 15, 3, 14, 6, 17,
    -- filter=36 channel=5
    -6, -6, -3, -8, 8, 1, 2, -3, 10,
    -- filter=36 channel=6
    10, -9, 2, 0, -3, 5, 10, 12, 10,
    -- filter=36 channel=7
    8, 12, 16, -4, 10, 16, 12, 2, 11,
    -- filter=36 channel=8
    -6, -4, 2, 9, 8, 13, 5, 23, 22,
    -- filter=36 channel=9
    -4, -3, -10, 7, 0, -11, 12, 13, -8,
    -- filter=36 channel=10
    12, -3, 0, 11, -3, 1, 14, 6, 13,
    -- filter=36 channel=11
    5, 5, -9, -3, 10, -1, -3, 12, -4,
    -- filter=36 channel=12
    10, 2, -7, -2, -7, 6, 0, 8, -9,
    -- filter=36 channel=13
    8, 8, 1, 11, 1, -2, 8, 21, 9,
    -- filter=36 channel=14
    0, -1, -2, 1, 0, 1, -7, 14, 13,
    -- filter=36 channel=15
    -6, 8, 4, 19, 6, 17, 2, 22, 18,
    -- filter=36 channel=16
    -7, -3, -5, -8, 5, -2, 3, 0, 8,
    -- filter=36 channel=17
    2, 9, -4, 14, 19, 3, 15, 1, 14,
    -- filter=36 channel=18
    23, 22, 9, 22, 33, 25, 10, 22, 20,
    -- filter=36 channel=19
    3, -11, -8, -9, -9, 3, -9, -13, 7,
    -- filter=36 channel=20
    11, 13, 0, 7, -1, 15, 13, 14, 0,
    -- filter=36 channel=21
    7, -4, 1, 2, 10, 2, -7, 3, 3,
    -- filter=36 channel=22
    6, 4, 0, 6, -2, 0, -8, 4, -7,
    -- filter=36 channel=23
    -1, -2, -5, 10, -3, 11, 1, 1, 0,
    -- filter=36 channel=24
    8, 3, -6, 0, -2, -2, 10, 19, 2,
    -- filter=36 channel=25
    -24, -29, -15, -11, -33, -29, -19, -29, -20,
    -- filter=36 channel=26
    -5, 0, 13, 9, 2, 11, -2, 2, 0,
    -- filter=36 channel=27
    -15, -16, -14, -6, -2, -22, -16, -15, -19,
    -- filter=36 channel=28
    -1, 12, 12, 7, 1, 6, 5, 21, 12,
    -- filter=36 channel=29
    -5, -6, -15, 4, -4, -9, 15, 10, 0,
    -- filter=36 channel=30
    3, 0, 11, 1, 14, 6, 1, -4, 18,
    -- filter=36 channel=31
    1, 12, -7, 5, 1, 8, 3, -10, -6,
    -- filter=36 channel=32
    0, -4, -16, -3, -19, -14, -6, -17, -12,
    -- filter=36 channel=33
    4, 8, -2, -9, -5, 4, 0, 1, -6,
    -- filter=36 channel=34
    -5, 7, 12, -4, 7, -1, -3, 0, 9,
    -- filter=36 channel=35
    -11, -12, -15, -1, -7, -13, -18, -17, -16,
    -- filter=36 channel=36
    2, 10, 2, -3, 0, -1, -9, 9, -8,
    -- filter=36 channel=37
    -1, -10, -10, -5, -7, -4, -7, -7, 3,
    -- filter=36 channel=38
    -16, -15, -7, 2, -17, -11, -7, -4, -4,
    -- filter=36 channel=39
    0, 6, -9, -8, -7, 1, -8, 1, 7,
    -- filter=36 channel=40
    4, -12, -11, 0, 2, -13, 0, -14, -9,
    -- filter=36 channel=41
    -3, -12, -9, 7, -4, -2, 6, 15, -4,
    -- filter=36 channel=42
    -6, -5, 3, 9, 3, -6, -3, 4, 3,
    -- filter=36 channel=43
    0, 7, -8, -10, -8, -16, -1, -1, -2,
    -- filter=36 channel=44
    -8, -16, -4, -13, -19, -2, 3, -16, -14,
    -- filter=36 channel=45
    -1, 1, 9, 5, -9, 9, 1, 7, -6,
    -- filter=36 channel=46
    -4, 13, 14, 9, 12, 14, 3, 1, 11,
    -- filter=36 channel=47
    8, 9, -2, -1, 0, 7, 2, 0, -9,
    -- filter=36 channel=48
    -7, 1, 2, 1, -3, 6, 13, 7, -5,
    -- filter=36 channel=49
    7, 13, 0, 22, 2, 14, 5, 13, 18,
    -- filter=36 channel=50
    12, 3, 19, -1, 14, -3, 13, 3, 12,
    -- filter=36 channel=51
    7, 7, 12, 22, 22, 22, 14, 20, 4,
    -- filter=36 channel=52
    2, -3, 10, -4, -9, -1, -3, 3, 3,
    -- filter=36 channel=53
    10, -10, 4, -6, -3, 4, 2, 0, 2,
    -- filter=36 channel=54
    -15, 1, 0, 0, -6, 3, -2, -8, 0,
    -- filter=36 channel=55
    2, -10, -3, -9, 7, -3, 2, -1, 9,
    -- filter=36 channel=56
    -4, 12, 1, 4, 4, 2, 5, 1, 0,
    -- filter=36 channel=57
    -7, 7, -4, 4, 5, 6, 1, -8, 10,
    -- filter=36 channel=58
    1, 7, 11, 11, 12, 15, 7, 12, 2,
    -- filter=36 channel=59
    -21, -10, -5, -13, -6, -8, -8, -13, -17,
    -- filter=36 channel=60
    -10, -5, -8, 0, 14, 12, 21, 16, 6,
    -- filter=36 channel=61
    -4, 4, 8, 5, 7, 14, 7, 18, 12,
    -- filter=36 channel=62
    -17, -3, -5, -4, -2, -6, -8, -9, 4,
    -- filter=36 channel=63
    -9, -5, 8, -8, 3, 2, -5, -8, -5,
    -- filter=37 channel=0
    1, -8, 1, 8, 1, -1, 7, 2, 4,
    -- filter=37 channel=1
    12, 27, 4, 8, 31, 13, 18, 19, 22,
    -- filter=37 channel=2
    19, 27, 24, 16, 37, 14, 21, 25, 19,
    -- filter=37 channel=3
    -1, 12, 1, -4, 10, 3, 9, -2, 4,
    -- filter=37 channel=4
    -16, 2, -12, -4, -12, -3, -9, -1, -11,
    -- filter=37 channel=5
    -4, 2, 3, -17, -2, 0, -4, 5, 6,
    -- filter=37 channel=6
    11, -2, 5, 15, 0, 13, 4, 8, 12,
    -- filter=37 channel=7
    2, 1, 13, -10, -7, 4, 9, 8, 0,
    -- filter=37 channel=8
    -9, -17, -18, -18, -17, -7, -14, -10, -9,
    -- filter=37 channel=9
    -32, -36, -21, -39, -48, -28, -25, -27, -24,
    -- filter=37 channel=10
    10, 9, 4, 24, 27, 19, 17, 14, 22,
    -- filter=37 channel=11
    5, -1, 0, -1, 1, -2, 8, 15, 0,
    -- filter=37 channel=12
    -3, 2, 10, -7, 0, 0, -1, -9, 4,
    -- filter=37 channel=13
    0, -1, 6, -17, -20, -14, 4, -1, -11,
    -- filter=37 channel=14
    -11, -2, 4, -9, 9, 9, -4, 4, 0,
    -- filter=37 channel=15
    -5, -16, 1, -9, -4, 4, 6, -8, 2,
    -- filter=37 channel=16
    -12, -1, 11, -6, -5, 12, -2, 11, 10,
    -- filter=37 channel=17
    -20, -19, 1, -13, -4, -7, 3, -1, -10,
    -- filter=37 channel=18
    -5, -4, 4, -7, -14, -2, -13, -17, -11,
    -- filter=37 channel=19
    4, 12, 17, 2, 8, 16, 0, 4, 17,
    -- filter=37 channel=20
    7, -1, 1, -12, 1, 4, 1, 2, -2,
    -- filter=37 channel=21
    -6, -2, -6, -5, 0, 6, 8, -8, -6,
    -- filter=37 channel=22
    -6, 6, 3, -5, 3, 5, -8, 3, 9,
    -- filter=37 channel=23
    3, 20, 2, 10, 29, 11, 21, 22, 7,
    -- filter=37 channel=24
    -21, -9, 4, -3, -3, -11, -5, -7, -3,
    -- filter=37 channel=25
    28, 20, 13, 29, 40, 34, 16, 23, 20,
    -- filter=37 channel=26
    0, 12, 16, 10, 0, 0, 18, 15, 6,
    -- filter=37 channel=27
    10, 11, 1, 22, 24, 8, 22, 26, 8,
    -- filter=37 channel=28
    -7, -1, 0, -8, -6, -7, -11, 0, 0,
    -- filter=37 channel=29
    -20, -11, -6, -24, -13, 4, -5, -11, 12,
    -- filter=37 channel=30
    15, 15, 14, 4, 23, 21, -2, 15, 24,
    -- filter=37 channel=31
    11, 4, 3, 10, 3, 1, -2, -7, 6,
    -- filter=37 channel=32
    20, 11, 8, 5, 22, 10, 22, 25, 3,
    -- filter=37 channel=33
    -3, 6, -3, 2, -4, 10, 9, -3, 2,
    -- filter=37 channel=34
    -9, -9, 10, -2, -10, -3, 0, -10, 4,
    -- filter=37 channel=35
    32, 32, 11, 33, 51, 21, 27, 25, 14,
    -- filter=37 channel=36
    -4, 0, -4, 10, 14, -3, 0, 11, 11,
    -- filter=37 channel=37
    -17, 1, 3, -14, 0, 7, -13, -6, 0,
    -- filter=37 channel=38
    -7, 15, 4, -3, 5, 14, 16, 25, 8,
    -- filter=37 channel=39
    -5, -4, 4, 1, 2, 9, 9, -4, 3,
    -- filter=37 channel=40
    3, 8, 3, 12, 4, 8, 9, 0, 9,
    -- filter=37 channel=41
    -10, -5, 10, -1, -2, 15, -4, 17, -3,
    -- filter=37 channel=42
    -4, -2, -7, 10, 0, 4, -2, 5, -7,
    -- filter=37 channel=43
    30, 22, 32, 26, 20, 24, 29, 26, 38,
    -- filter=37 channel=44
    4, 4, 10, 7, 25, 23, 12, 22, 14,
    -- filter=37 channel=45
    0, 9, 2, -7, 0, 0, -5, 0, 0,
    -- filter=37 channel=46
    -8, -4, -3, 4, -3, 2, -12, -6, 3,
    -- filter=37 channel=47
    -10, 2, -5, -4, 4, -9, -3, 0, 6,
    -- filter=37 channel=48
    -4, 7, -3, 8, 0, -7, -7, -1, 7,
    -- filter=37 channel=49
    18, 0, 2, 9, 22, 13, 2, 17, 4,
    -- filter=37 channel=50
    6, 5, 5, 2, 10, 10, 5, 15, 9,
    -- filter=37 channel=51
    11, -2, -3, 1, 6, -3, -1, 13, 5,
    -- filter=37 channel=52
    -7, -7, 1, -5, 4, 0, -8, -6, -7,
    -- filter=37 channel=53
    18, 17, 2, 18, 20, 18, 0, 8, 16,
    -- filter=37 channel=54
    -16, -19, -22, -33, -31, -25, -22, -35, -26,
    -- filter=37 channel=55
    2, 7, 0, 0, 3, -7, 9, 4, -6,
    -- filter=37 channel=56
    7, -4, 10, 3, -6, 2, 2, 0, -5,
    -- filter=37 channel=57
    2, 10, 1, 10, -7, 1, -7, 0, -4,
    -- filter=37 channel=58
    1, 4, 15, 10, 7, 14, 3, 15, 6,
    -- filter=37 channel=59
    0, 13, -5, -1, 8, 4, 13, 2, 18,
    -- filter=37 channel=60
    -11, -24, -8, -12, -2, -9, -16, 1, 0,
    -- filter=37 channel=61
    -10, -22, -9, -17, -15, -13, 0, 3, 0,
    -- filter=37 channel=62
    6, -4, 3, 7, 7, -6, -3, 2, 10,
    -- filter=37 channel=63
    -6, 5, -6, 9, 1, 8, -1, 5, -10,
    -- filter=38 channel=0
    4, -1, 9, -9, 13, -3, -11, -1, 5,
    -- filter=38 channel=1
    -5, -4, 7, 0, 4, 15, -14, -9, -5,
    -- filter=38 channel=2
    -1, 0, -1, 0, -5, 11, -14, 1, -1,
    -- filter=38 channel=3
    -8, 0, 3, -7, 13, -5, 3, -8, -3,
    -- filter=38 channel=4
    -6, -6, -6, -8, 11, 5, -8, -7, -7,
    -- filter=38 channel=5
    -5, 0, -5, -2, -2, 0, 7, 7, -9,
    -- filter=38 channel=6
    0, 12, 6, -5, 2, -8, -5, -13, -9,
    -- filter=38 channel=7
    0, -13, -9, 7, 4, 4, -3, 6, -11,
    -- filter=38 channel=8
    -7, 7, 11, -8, 15, 8, -21, -4, -5,
    -- filter=38 channel=9
    4, 9, 5, 1, 8, 4, -1, 1, -13,
    -- filter=38 channel=10
    -6, 1, 8, -5, 0, 6, -9, -6, 14,
    -- filter=38 channel=11
    -5, 7, 5, 2, 4, 15, -4, 7, -3,
    -- filter=38 channel=12
    9, 4, 3, 3, 5, -3, 5, -5, 0,
    -- filter=38 channel=13
    9, -5, -11, 8, 3, -7, 1, 2, 4,
    -- filter=38 channel=14
    -11, -6, 0, 4, 2, 1, 7, -6, -5,
    -- filter=38 channel=15
    14, 3, -5, -6, 8, 2, 0, 0, -9,
    -- filter=38 channel=16
    -5, 13, -2, 3, 7, 9, -21, -1, -19,
    -- filter=38 channel=17
    4, 10, 3, -12, 11, -2, -5, -5, -5,
    -- filter=38 channel=18
    3, 5, 0, 8, -3, -7, 9, -5, -6,
    -- filter=38 channel=19
    2, -6, -4, -4, 2, -3, -4, 3, 6,
    -- filter=38 channel=20
    6, -13, -4, 6, -10, -7, -8, 0, -7,
    -- filter=38 channel=21
    0, 8, 10, -4, -10, 4, 0, 5, -7,
    -- filter=38 channel=22
    -1, 9, 6, -10, -6, 4, 2, 3, -9,
    -- filter=38 channel=23
    -15, 8, 6, 1, 3, 10, -9, 7, 12,
    -- filter=38 channel=24
    0, 6, 2, -5, 10, 4, -1, 0, 5,
    -- filter=38 channel=25
    8, 16, 18, -9, -1, 7, -4, -5, -2,
    -- filter=38 channel=26
    2, 1, -8, 7, 4, -3, -2, -2, 5,
    -- filter=38 channel=27
    7, 12, 5, 0, -3, 4, -19, 1, 3,
    -- filter=38 channel=28
    7, 10, 2, 0, 6, 4, -17, -9, -15,
    -- filter=38 channel=29
    18, 12, 6, 1, 15, -1, -10, 0, -23,
    -- filter=38 channel=30
    -12, -13, -6, -10, -21, -6, -12, -17, -14,
    -- filter=38 channel=31
    0, 8, -6, 3, 1, 8, -3, 11, 1,
    -- filter=38 channel=32
    -16, -10, 4, -3, 2, 0, 1, -1, 2,
    -- filter=38 channel=33
    -5, -4, 4, -3, 6, 7, 0, 0, -2,
    -- filter=38 channel=34
    4, -4, -8, -9, 1, -4, -6, -7, 7,
    -- filter=38 channel=35
    1, 6, 19, -8, -7, 7, -13, 1, 7,
    -- filter=38 channel=36
    2, 4, 9, 1, -2, 10, 0, 5, 3,
    -- filter=38 channel=37
    5, -7, 6, 8, 9, 6, -3, 0, -6,
    -- filter=38 channel=38
    10, -1, 3, -7, 12, 6, -9, -11, 4,
    -- filter=38 channel=39
    3, 6, 7, -9, 7, 4, 8, 2, 10,
    -- filter=38 channel=40
    -4, 1, -4, -4, 9, 10, 2, -4, 9,
    -- filter=38 channel=41
    -1, 16, 19, 3, 9, 10, -14, -1, -4,
    -- filter=38 channel=42
    -4, 2, 6, 2, -1, -5, 4, 2, -4,
    -- filter=38 channel=43
    -20, -14, -6, 0, -9, -10, 2, -10, -3,
    -- filter=38 channel=44
    4, -1, 1, -8, 4, -8, -2, 8, 1,
    -- filter=38 channel=45
    6, -4, 0, -2, -9, 6, -10, 1, 8,
    -- filter=38 channel=46
    -8, 1, -3, -1, -1, -3, 0, -8, -4,
    -- filter=38 channel=47
    -3, -7, -4, -7, 3, 4, 7, -1, -7,
    -- filter=38 channel=48
    7, -1, 3, 13, 5, -1, -13, -12, -3,
    -- filter=38 channel=49
    0, 0, 0, -9, -5, -3, -1, -1, -6,
    -- filter=38 channel=50
    -6, -13, -6, -5, -1, -11, -8, 0, 5,
    -- filter=38 channel=51
    -5, -3, 3, 6, -8, 0, 0, 13, -4,
    -- filter=38 channel=52
    3, 4, -7, -2, -2, 1, -5, 9, 5,
    -- filter=38 channel=53
    -8, -16, 4, 0, -9, 4, -3, -5, 3,
    -- filter=38 channel=54
    6, -2, 9, 11, -6, -8, -4, -4, 0,
    -- filter=38 channel=55
    3, 10, -4, -7, 3, -4, 2, 7, 2,
    -- filter=38 channel=56
    -11, -2, 1, 6, -7, 7, 4, -6, -10,
    -- filter=38 channel=57
    0, 7, 7, 0, 5, -2, -8, 5, -9,
    -- filter=38 channel=58
    -5, 9, 1, -3, -4, -11, 5, 10, -3,
    -- filter=38 channel=59
    1, 19, 0, 0, 10, 11, 2, -6, -12,
    -- filter=38 channel=60
    12, 23, 0, 14, 14, 12, -6, 1, -4,
    -- filter=38 channel=61
    -8, 10, 6, 8, 16, 13, 0, 0, -5,
    -- filter=38 channel=62
    -3, 3, 3, -10, 14, 6, -9, -2, -9,
    -- filter=38 channel=63
    6, -3, -8, -2, 3, -7, -9, -6, 9,
    -- filter=39 channel=0
    4, -9, 0, -1, -7, 2, -6, -2, -4,
    -- filter=39 channel=1
    -10, -11, 0, 6, -5, -4, 9, -5, -6,
    -- filter=39 channel=2
    -8, -7, -9, 6, 0, -13, -10, -5, -15,
    -- filter=39 channel=3
    3, 3, 5, -1, -5, 0, 4, -8, -5,
    -- filter=39 channel=4
    9, 8, -10, -4, 10, -6, -4, 0, -6,
    -- filter=39 channel=5
    -6, 8, 5, 9, 1, -5, 5, 7, 2,
    -- filter=39 channel=6
    -6, 0, 1, 7, 1, 1, -3, -5, 0,
    -- filter=39 channel=7
    -1, -10, 3, 8, 0, -2, -1, -4, 4,
    -- filter=39 channel=8
    -12, -1, 0, -5, 14, -5, -1, -9, 1,
    -- filter=39 channel=9
    -1, 14, 20, 25, 31, 38, 13, 32, 24,
    -- filter=39 channel=10
    5, 8, -9, 8, -6, 0, 11, 9, -3,
    -- filter=39 channel=11
    -13, -4, 6, 6, -9, 5, -6, -7, -9,
    -- filter=39 channel=12
    9, -9, -1, 2, 4, 7, 12, 4, 11,
    -- filter=39 channel=13
    -7, 9, -2, 5, -2, 0, -5, 5, 1,
    -- filter=39 channel=14
    -1, -9, 0, 4, 8, 0, -11, 8, -4,
    -- filter=39 channel=15
    -5, 10, -4, 15, 6, 0, 1, 5, 0,
    -- filter=39 channel=16
    -5, -6, -11, -8, 12, 10, -4, 4, -10,
    -- filter=39 channel=17
    -8, -6, -8, 10, 5, 4, 4, 5, 1,
    -- filter=39 channel=18
    0, 9, 12, 5, 18, 15, 12, 12, -1,
    -- filter=39 channel=19
    -9, 12, 3, 6, 6, 5, 7, 5, 5,
    -- filter=39 channel=20
    0, 14, 14, 5, 13, 6, 15, 16, 1,
    -- filter=39 channel=21
    8, 4, 7, 11, -6, 3, -4, 7, 10,
    -- filter=39 channel=22
    6, -6, 2, 8, -4, -5, 0, 6, 9,
    -- filter=39 channel=23
    1, 3, -4, 5, -3, -4, -2, -3, 2,
    -- filter=39 channel=24
    6, 3, -1, 0, -3, 0, -7, 1, -6,
    -- filter=39 channel=25
    4, -8, -16, 7, 0, 1, 1, 2, -3,
    -- filter=39 channel=26
    2, -8, -7, -6, -1, -4, -10, -3, -2,
    -- filter=39 channel=27
    5, -13, -8, 0, -8, -1, 1, -10, -14,
    -- filter=39 channel=28
    5, 11, 6, 5, 17, 18, 5, 10, 4,
    -- filter=39 channel=29
    4, 8, -5, 10, 19, 0, 7, 14, 4,
    -- filter=39 channel=30
    -13, -11, -5, -5, -13, -2, -19, -8, -14,
    -- filter=39 channel=31
    13, 6, 4, 11, 8, 0, 6, 11, -2,
    -- filter=39 channel=32
    3, 1, 0, -1, -10, -1, 3, 0, -5,
    -- filter=39 channel=33
    -9, -1, 8, 5, -1, -8, -4, -8, 3,
    -- filter=39 channel=34
    -8, -3, -4, -7, -4, 0, -10, -2, 4,
    -- filter=39 channel=35
    -1, 1, -7, 0, -14, -10, -4, -19, -7,
    -- filter=39 channel=36
    -4, -6, 4, 11, 3, -7, 8, 1, -5,
    -- filter=39 channel=37
    -7, 3, 3, 11, 5, 4, 10, 3, 10,
    -- filter=39 channel=38
    -11, -14, -14, -8, 1, 0, -7, -2, -10,
    -- filter=39 channel=39
    -8, -6, -8, 9, 4, 8, -1, -9, 6,
    -- filter=39 channel=40
    9, 8, -10, -5, 5, -9, 8, 6, 7,
    -- filter=39 channel=41
    -1, -7, 5, 7, -7, 8, 2, -9, 1,
    -- filter=39 channel=42
    3, 7, 8, 0, -1, 9, 2, -9, -6,
    -- filter=39 channel=43
    -1, -1, -9, -9, -15, -12, 2, -8, -2,
    -- filter=39 channel=44
    2, 7, -5, 4, -8, 7, -2, -8, -5,
    -- filter=39 channel=45
    6, -2, -2, -10, 6, -3, -4, -5, -5,
    -- filter=39 channel=46
    7, -1, -9, 4, 1, -5, 5, -1, -8,
    -- filter=39 channel=47
    0, -5, 10, 3, 0, 2, 3, -7, -9,
    -- filter=39 channel=48
    -7, 8, -3, -3, 0, 9, 3, -7, -3,
    -- filter=39 channel=49
    6, 2, -2, 0, -5, 4, -8, 3, 1,
    -- filter=39 channel=50
    3, 4, 6, -10, -5, -7, -6, -8, -4,
    -- filter=39 channel=51
    -1, 8, 11, 4, 11, -5, 6, -1, 8,
    -- filter=39 channel=52
    6, 7, 4, 10, 8, -1, 8, -4, -1,
    -- filter=39 channel=53
    -11, -6, -7, -11, -7, -6, -3, 0, 0,
    -- filter=39 channel=54
    2, 6, 15, 14, 32, 12, 5, 11, 22,
    -- filter=39 channel=55
    6, 1, -1, -6, -8, -2, 10, 10, 8,
    -- filter=39 channel=56
    -3, -3, -10, 1, -2, 2, 8, -4, 5,
    -- filter=39 channel=57
    -5, 10, -2, 5, -6, -7, 7, 1, 3,
    -- filter=39 channel=58
    4, 9, 5, 9, -4, 11, 3, 9, 12,
    -- filter=39 channel=59
    5, -11, 1, -4, 8, 4, -1, 3, -9,
    -- filter=39 channel=60
    -10, -2, -15, 0, -2, 1, 3, -1, -7,
    -- filter=39 channel=61
    -1, 7, -13, 7, 6, -2, 8, 6, 1,
    -- filter=39 channel=62
    -5, 0, -10, 2, -8, 0, -2, -5, 2,
    -- filter=39 channel=63
    0, 5, -1, -8, 4, 8, 7, -4, 2,
    -- filter=40 channel=0
    4, 5, -5, 5, -11, -11, 1, -6, -6,
    -- filter=40 channel=1
    1, 7, 2, 1, -5, 8, 5, 10, 0,
    -- filter=40 channel=2
    4, 12, 12, -1, -6, 2, 0, 3, 0,
    -- filter=40 channel=3
    -11, 4, 4, 1, -10, -6, -10, -18, -5,
    -- filter=40 channel=4
    0, 3, -5, -7, 1, 6, 0, -8, -9,
    -- filter=40 channel=5
    -5, -1, 0, 4, -4, -12, -12, -8, -7,
    -- filter=40 channel=6
    0, 9, 14, 13, 10, 1, 8, 9, 7,
    -- filter=40 channel=7
    -4, 2, 1, 0, 0, 0, -6, 1, -2,
    -- filter=40 channel=8
    0, 1, -2, -2, 6, -8, -11, 0, -9,
    -- filter=40 channel=9
    22, 14, 13, 10, 13, 27, 7, 9, 24,
    -- filter=40 channel=10
    14, -3, 0, 13, -5, -4, 2, -2, -5,
    -- filter=40 channel=11
    -7, 0, 12, -6, 0, -4, -4, -7, 0,
    -- filter=40 channel=12
    0, -8, 5, -3, 1, -2, 2, 9, -3,
    -- filter=40 channel=13
    11, 14, 0, 5, -3, 16, 14, 8, -6,
    -- filter=40 channel=14
    4, 6, 9, -3, 1, -8, 2, -6, -10,
    -- filter=40 channel=15
    12, 14, 3, 10, -6, 8, 8, 7, 2,
    -- filter=40 channel=16
    2, 10, 17, 8, -7, -6, 0, 1, -1,
    -- filter=40 channel=17
    3, 2, 10, 3, 4, -8, -10, -9, -7,
    -- filter=40 channel=18
    9, 5, 9, 15, 15, 0, 19, 20, 13,
    -- filter=40 channel=19
    10, 22, 10, 14, 21, 1, 5, 11, 6,
    -- filter=40 channel=20
    17, 11, 4, 14, 16, 14, 13, 0, 4,
    -- filter=40 channel=21
    -4, -7, 8, -6, -8, -2, 1, 1, -7,
    -- filter=40 channel=22
    -7, 9, 3, 5, -9, -3, -9, -1, 6,
    -- filter=40 channel=23
    4, 7, 10, 1, 3, 4, 1, -5, 1,
    -- filter=40 channel=24
    8, 7, 3, -8, 5, 7, 3, 2, 4,
    -- filter=40 channel=25
    -3, 13, 7, 0, 0, -3, -12, 1, 4,
    -- filter=40 channel=26
    -3, -6, 3, 4, -5, 9, 3, -6, 9,
    -- filter=40 channel=27
    -4, 0, 5, -10, -15, -11, -6, 0, -8,
    -- filter=40 channel=28
    10, 10, 16, 4, 10, 11, -4, 9, 0,
    -- filter=40 channel=29
    12, 4, 0, -3, 7, 10, 8, 2, -5,
    -- filter=40 channel=30
    -13, 6, -5, 2, 10, -6, -9, 0, 1,
    -- filter=40 channel=31
    -7, -4, -8, -6, -3, -3, 1, 8, -3,
    -- filter=40 channel=32
    -10, -8, 5, -12, -6, -1, -5, -6, -6,
    -- filter=40 channel=33
    -7, 2, 10, 10, 6, -4, -3, 1, -10,
    -- filter=40 channel=34
    9, 10, 7, 7, -9, -3, -1, 6, -8,
    -- filter=40 channel=35
    -10, -5, 4, -4, 2, -10, -9, -15, 1,
    -- filter=40 channel=36
    8, 0, -5, 10, -6, 0, 2, 0, -7,
    -- filter=40 channel=37
    -7, -6, -9, -11, -5, -11, -3, -17, -16,
    -- filter=40 channel=38
    -2, 7, -8, -9, 1, 5, 1, -13, 7,
    -- filter=40 channel=39
    6, 0, -6, 3, 6, 1, 6, -5, 4,
    -- filter=40 channel=40
    -9, -6, 1, -2, -5, 4, -4, -11, -8,
    -- filter=40 channel=41
    0, 0, 3, -2, -17, 1, -9, -17, -5,
    -- filter=40 channel=42
    -6, -3, -1, -4, -3, -1, -2, -2, 0,
    -- filter=40 channel=43
    0, 1, -9, -2, -2, -4, 10, 1, 6,
    -- filter=40 channel=44
    2, -1, -3, 5, -2, -2, -5, 8, -4,
    -- filter=40 channel=45
    1, 1, 3, -6, -3, 10, -7, -4, -2,
    -- filter=40 channel=46
    2, -3, 0, -5, 0, 0, 0, -5, -10,
    -- filter=40 channel=47
    10, 6, -2, 10, 6, 0, -5, -10, 10,
    -- filter=40 channel=48
    6, 10, 3, 13, -3, 12, 5, -5, -5,
    -- filter=40 channel=49
    6, 1, 0, 3, -3, -1, 5, -2, 0,
    -- filter=40 channel=50
    6, 1, 8, -2, 8, 8, 4, -2, -6,
    -- filter=40 channel=51
    1, 0, 5, 3, 7, -5, 9, 6, 0,
    -- filter=40 channel=52
    8, -8, 10, -7, -9, 6, 9, 5, -1,
    -- filter=40 channel=53
    -8, -1, 7, -8, 0, 5, -10, 0, -3,
    -- filter=40 channel=54
    3, 11, 5, 1, 4, 0, -2, 3, 4,
    -- filter=40 channel=55
    -8, 6, 8, 0, 5, 9, -6, 3, 7,
    -- filter=40 channel=56
    -8, -3, -7, -7, -9, 8, 3, -5, 5,
    -- filter=40 channel=57
    1, 0, -4, 8, -3, 0, -9, -4, -4,
    -- filter=40 channel=58
    12, 13, 17, 12, 8, 0, 13, 13, 5,
    -- filter=40 channel=59
    0, -2, 1, -13, -4, 1, -19, -11, -4,
    -- filter=40 channel=60
    -6, -11, 2, 7, 1, -14, -5, 1, 0,
    -- filter=40 channel=61
    -5, -9, -5, 3, -8, -4, -4, -4, -12,
    -- filter=40 channel=62
    -13, -5, -6, -3, -1, 1, -18, -15, 0,
    -- filter=40 channel=63
    4, 10, -3, 2, 7, 7, 3, 4, 1,
    -- filter=41 channel=0
    9, -8, -3, 23, -21, 2, 23, 3, 0,
    -- filter=41 channel=1
    -3, 6, -33, 4, 4, -41, -6, 7, -18,
    -- filter=41 channel=2
    22, -8, -22, 25, -2, -19, 9, -8, 4,
    -- filter=41 channel=3
    28, -13, -17, 16, 5, -5, 7, -7, 5,
    -- filter=41 channel=4
    4, -4, -8, 13, 1, -12, 2, -4, 5,
    -- filter=41 channel=5
    9, 24, -10, 2, 27, 0, -1, 18, 1,
    -- filter=41 channel=6
    16, -8, -3, 11, -19, -14, 13, -5, 2,
    -- filter=41 channel=7
    7, 31, 15, 3, 30, 18, 16, 29, 16,
    -- filter=41 channel=8
    37, 0, -42, 28, -3, -43, 13, 11, -17,
    -- filter=41 channel=9
    12, -9, 1, 19, -1, -3, -5, -16, 3,
    -- filter=41 channel=10
    1, -12, 0, -1, -14, 0, 1, -12, 11,
    -- filter=41 channel=11
    10, 11, -31, 21, 17, -27, -1, 19, -16,
    -- filter=41 channel=12
    6, 1, -9, -7, -1, 1, -4, -9, -2,
    -- filter=41 channel=13
    14, -27, 14, 9, -22, 2, 13, -1, -1,
    -- filter=41 channel=14
    20, 36, 2, 16, 22, 11, 14, 26, 9,
    -- filter=41 channel=15
    42, -25, -14, 47, -33, -15, 27, -4, -1,
    -- filter=41 channel=16
    38, -5, -37, 44, -25, -44, 18, 2, -11,
    -- filter=41 channel=17
    10, 10, -31, 14, 25, -32, 18, 12, -7,
    -- filter=41 channel=18
    -5, -14, -1, 0, -6, 5, 5, 1, 0,
    -- filter=41 channel=19
    -1, 22, -27, -13, 33, -20, -6, 17, -14,
    -- filter=41 channel=20
    3, 4, 21, 10, -1, 22, 10, 7, 11,
    -- filter=41 channel=21
    -5, 3, 1, 2, -6, 8, -8, -6, 8,
    -- filter=41 channel=22
    5, 10, 7, -9, -7, 8, -3, 5, -2,
    -- filter=41 channel=23
    9, -2, -18, 3, 7, -22, 9, 9, -20,
    -- filter=41 channel=24
    5, 19, -22, 7, 27, -30, 0, 22, -6,
    -- filter=41 channel=25
    22, -19, -20, 14, -29, -20, 4, -16, -21,
    -- filter=41 channel=26
    32, 11, 28, 30, 10, 32, 34, 21, 30,
    -- filter=41 channel=27
    25, -1, -30, 27, 1, -43, 20, 15, -19,
    -- filter=41 channel=28
    10, 18, -40, 12, 6, -38, -7, 14, -12,
    -- filter=41 channel=29
    45, -37, -19, 34, -28, -26, 26, -17, -9,
    -- filter=41 channel=30
    51, 92, 0, 47, 101, 16, 37, 97, 23,
    -- filter=41 channel=31
    -12, 5, 3, 4, 5, -6, 5, -12, -3,
    -- filter=41 channel=32
    9, 13, -8, 12, 7, -9, 13, 11, 0,
    -- filter=41 channel=33
    -9, -4, 2, 3, 1, 0, 2, 7, 0,
    -- filter=41 channel=34
    17, 13, 14, 20, 2, 10, 4, 19, 19,
    -- filter=41 channel=35
    22, 0, -29, 35, 4, -20, 22, -1, -8,
    -- filter=41 channel=36
    0, 6, 6, -7, 0, -7, 6, 3, 9,
    -- filter=41 channel=37
    2, -2, 0, 10, 2, -14, 7, 6, -21,
    -- filter=41 channel=38
    21, -10, -24, 41, -9, -41, 19, 9, -29,
    -- filter=41 channel=39
    0, -3, 3, -7, -4, 5, -1, 9, -4,
    -- filter=41 channel=40
    -1, -2, -8, 11, 3, 7, -5, 0, -5,
    -- filter=41 channel=41
    51, -10, -36, 44, -9, -45, 31, 18, -5,
    -- filter=41 channel=42
    2, -6, 3, -8, 2, 8, -7, 5, 6,
    -- filter=41 channel=43
    -6, 12, 23, 10, 3, -3, 7, -7, -8,
    -- filter=41 channel=44
    -2, 28, -12, 6, 16, -8, -3, 31, -9,
    -- filter=41 channel=45
    7, -7, 8, 8, 2, -9, -6, -10, 0,
    -- filter=41 channel=46
    29, 12, 27, 40, 11, 19, 21, 15, 20,
    -- filter=41 channel=47
    -5, -4, 9, 1, 5, -1, -5, -7, 1,
    -- filter=41 channel=48
    20, -18, 13, 20, -19, -9, 21, -8, 0,
    -- filter=41 channel=49
    22, -6, -11, 20, 6, -14, 0, 14, 10,
    -- filter=41 channel=50
    19, 39, 21, 16, 58, 0, 24, 28, -4,
    -- filter=41 channel=51
    -9, -7, 10, 9, 5, 4, 1, -5, 3,
    -- filter=41 channel=52
    -9, 4, 1, 9, -9, -7, -3, -2, 4,
    -- filter=41 channel=53
    11, 60, -4, 26, 78, 1, 25, 56, 5,
    -- filter=41 channel=54
    14, 4, -18, 15, 8, -8, -1, 5, -14,
    -- filter=41 channel=55
    5, 5, -4, -5, 9, -3, 5, 2, -4,
    -- filter=41 channel=56
    8, 7, 20, 1, 3, 20, 9, 3, 19,
    -- filter=41 channel=57
    -3, 0, 5, -4, -6, -3, -8, -2, -6,
    -- filter=41 channel=58
    2, -11, 5, -11, -3, 5, -13, 1, 11,
    -- filter=41 channel=59
    29, -23, 2, 37, -18, -19, 24, 3, -11,
    -- filter=41 channel=60
    44, -25, -25, 70, -16, -43, 46, 5, -18,
    -- filter=41 channel=61
    29, 12, -32, 43, 23, -49, 28, 14, -13,
    -- filter=41 channel=62
    18, 4, -26, 14, 5, -22, -5, 20, -12,
    -- filter=41 channel=63
    -1, -4, 8, 4, 0, -9, 0, 6, 9,
    -- filter=42 channel=0
    -6, 3, -2, 12, 0, -5, 9, 7, 7,
    -- filter=42 channel=1
    16, 4, 8, 4, 0, 2, 16, 15, -1,
    -- filter=42 channel=2
    7, 14, 7, 19, 5, -1, 14, 5, 4,
    -- filter=42 channel=3
    3, 10, -6, -6, -2, -9, 12, -4, -11,
    -- filter=42 channel=4
    -7, -6, -5, -9, -2, 8, -9, 0, -2,
    -- filter=42 channel=5
    -9, -13, -2, 0, 0, -9, 6, -2, -8,
    -- filter=42 channel=6
    6, 0, -1, 2, -3, 7, 7, 8, -2,
    -- filter=42 channel=7
    -10, -5, -1, -2, -3, 1, -2, 3, 2,
    -- filter=42 channel=8
    8, 0, 2, -5, -7, 12, 1, 7, -3,
    -- filter=42 channel=9
    -3, 3, 6, -17, -10, -5, -13, 1, 6,
    -- filter=42 channel=10
    9, 11, 3, 5, 9, 1, 8, 13, -3,
    -- filter=42 channel=11
    8, -5, -10, 1, 13, 11, -2, -7, -7,
    -- filter=42 channel=12
    -10, -6, 0, -9, 9, -9, -9, -6, -3,
    -- filter=42 channel=13
    -14, -14, 5, -3, -7, -10, -8, -5, 2,
    -- filter=42 channel=14
    3, -5, -11, -13, -6, 4, -7, 0, -6,
    -- filter=42 channel=15
    -8, -10, -6, 5, -5, 5, -7, 2, -7,
    -- filter=42 channel=16
    0, -5, 0, -5, 8, -3, 5, 1, 4,
    -- filter=42 channel=17
    0, -6, 2, 0, 1, -3, 0, -5, 0,
    -- filter=42 channel=18
    -13, 0, 2, -4, -3, -3, -12, -12, -7,
    -- filter=42 channel=19
    -7, 1, 8, 3, 8, -5, 9, -5, 2,
    -- filter=42 channel=20
    2, 0, -10, -5, -4, -6, -4, -9, -1,
    -- filter=42 channel=21
    10, 7, -4, 2, -6, 9, -2, -3, -5,
    -- filter=42 channel=22
    2, 0, -3, 6, 3, 5, 5, -2, 5,
    -- filter=42 channel=23
    13, 7, -12, 7, 1, -6, 3, 7, 0,
    -- filter=42 channel=24
    -1, -6, -2, 7, 0, -1, 8, 3, 0,
    -- filter=42 channel=25
    11, 5, 5, 8, 20, 11, 3, 3, 8,
    -- filter=42 channel=26
    -7, -12, -12, 5, 0, -7, -8, -4, 0,
    -- filter=42 channel=27
    12, 8, -12, 21, 9, 10, 7, 10, 10,
    -- filter=42 channel=28
    8, -5, 13, -2, 3, 13, 6, -2, -8,
    -- filter=42 channel=29
    5, -9, 8, -6, -1, 0, -1, 6, -2,
    -- filter=42 channel=30
    -5, -13, -15, -22, -24, -18, -12, -11, -12,
    -- filter=42 channel=31
    11, 9, 8, -3, 8, -10, 10, -10, -1,
    -- filter=42 channel=32
    11, -3, 3, 13, -3, -2, -2, 9, 0,
    -- filter=42 channel=33
    -5, 3, -3, 0, -3, -10, -8, -3, 3,
    -- filter=42 channel=34
    -11, 0, -8, 6, 0, -5, 0, 0, -11,
    -- filter=42 channel=35
    5, 6, -4, 12, 7, -1, 16, 16, 0,
    -- filter=42 channel=36
    11, -7, 8, -1, -6, 7, 11, -1, -4,
    -- filter=42 channel=37
    -6, 9, 2, -4, -6, -1, -9, -4, 5,
    -- filter=42 channel=38
    12, -1, -7, 11, 5, 6, 9, 16, -2,
    -- filter=42 channel=39
    -5, -7, 6, 0, 0, 10, -2, 7, 2,
    -- filter=42 channel=40
    7, -7, -5, -7, 3, -1, 0, 0, 0,
    -- filter=42 channel=41
    5, 10, 2, 1, 15, 9, 0, 7, -2,
    -- filter=42 channel=42
    8, -6, 3, -8, 5, -9, -7, 6, 2,
    -- filter=42 channel=43
    5, -6, -2, -9, 0, 11, 7, 11, 14,
    -- filter=42 channel=44
    8, -2, 0, 0, 12, -1, 0, -6, -11,
    -- filter=42 channel=45
    3, 8, 2, -1, 7, 8, -6, 1, 0,
    -- filter=42 channel=46
    -17, -12, -5, -9, -2, -1, 0, -7, -17,
    -- filter=42 channel=47
    -1, -3, 6, -10, -1, 3, -4, -1, 8,
    -- filter=42 channel=48
    -9, -3, -1, 2, -5, -5, 4, -9, 5,
    -- filter=42 channel=49
    11, 10, -5, 3, 11, 4, 5, 0, -7,
    -- filter=42 channel=50
    -15, -9, -2, -16, -15, -9, -18, -9, -10,
    -- filter=42 channel=51
    -4, 4, -12, 11, -3, -12, 11, -3, 8,
    -- filter=42 channel=52
    3, 1, 5, 8, 9, -3, 7, 8, 5,
    -- filter=42 channel=53
    -16, -15, -9, -8, -2, -15, 2, 2, -7,
    -- filter=42 channel=54
    2, -8, 8, -9, -16, 4, -12, -8, 0,
    -- filter=42 channel=55
    -8, 2, 9, 0, -4, 9, -3, 4, -1,
    -- filter=42 channel=56
    -9, -13, 3, -12, -9, -8, 2, 4, -13,
    -- filter=42 channel=57
    -9, 2, 10, 0, 8, -3, 0, -7, -4,
    -- filter=42 channel=58
    -6, 3, 5, 0, -8, -3, -5, 4, -9,
    -- filter=42 channel=59
    0, 1, 1, 16, 0, 4, -3, -4, 3,
    -- filter=42 channel=60
    2, -7, 0, 0, -5, 0, 8, -10, -11,
    -- filter=42 channel=61
    6, -12, -6, -3, -2, 7, 10, -3, -1,
    -- filter=42 channel=62
    -3, 5, -9, 12, -2, 4, -6, -7, -4,
    -- filter=42 channel=63
    -2, 5, -1, 6, -3, -8, -9, -3, 8,
    -- filter=43 channel=0
    0, -3, 6, -10, -2, -6, -16, -15, -5,
    -- filter=43 channel=1
    9, 18, 7, 15, 11, 13, 4, 10, 8,
    -- filter=43 channel=2
    0, 12, 13, 3, -7, 4, -8, -5, -4,
    -- filter=43 channel=3
    4, 10, 16, 13, -2, 8, 9, 5, 1,
    -- filter=43 channel=4
    9, -1, 8, -6, -3, 4, -9, -2, -14,
    -- filter=43 channel=5
    2, 3, 11, 0, 13, -1, 5, 3, 1,
    -- filter=43 channel=6
    -2, 7, 3, 6, 3, 2, -10, -9, 0,
    -- filter=43 channel=7
    0, 2, 10, 10, 11, 5, 1, 10, 10,
    -- filter=43 channel=8
    14, 9, 22, -15, 1, -7, -19, -29, -11,
    -- filter=43 channel=9
    12, 25, 18, 11, 21, 25, 5, 6, 17,
    -- filter=43 channel=10
    -3, -8, -2, 2, 0, 10, 7, 1, -1,
    -- filter=43 channel=11
    9, 17, 11, -5, -2, -1, -5, -7, -10,
    -- filter=43 channel=12
    -5, 3, 7, 0, -3, 9, -5, 5, 10,
    -- filter=43 channel=13
    -1, 5, 13, 0, 16, 13, -14, -3, -14,
    -- filter=43 channel=14
    -7, 8, -8, 9, -6, -4, 5, 1, -5,
    -- filter=43 channel=15
    7, 13, 13, -12, 1, -4, -21, -11, -20,
    -- filter=43 channel=16
    4, 18, 29, -12, 10, 9, -21, -13, -12,
    -- filter=43 channel=17
    -3, 9, 1, -12, -14, -3, 0, -23, -17,
    -- filter=43 channel=18
    -4, 2, -8, -7, -13, -4, 4, -4, -4,
    -- filter=43 channel=19
    -3, 11, 7, 0, 19, 5, 15, 11, 10,
    -- filter=43 channel=20
    16, 16, 16, 6, 19, 7, -5, 9, 19,
    -- filter=43 channel=21
    -8, -6, -2, -5, -8, 1, -7, 2, 0,
    -- filter=43 channel=22
    -8, 9, 4, -1, 10, -4, -3, 7, 0,
    -- filter=43 channel=23
    -1, -5, 2, 0, 6, -5, 3, 1, -6,
    -- filter=43 channel=24
    8, -6, -1, 5, -10, 9, 0, -17, -17,
    -- filter=43 channel=25
    0, 9, 7, 0, 12, 19, -7, -7, -1,
    -- filter=43 channel=26
    14, 12, 9, 18, 9, 9, 9, 19, -3,
    -- filter=43 channel=27
    16, 22, 11, -10, -2, 1, -11, -18, -5,
    -- filter=43 channel=28
    11, 17, -1, -5, 3, -8, -12, -14, 0,
    -- filter=43 channel=29
    12, 25, 9, -2, 3, 1, -23, -21, -10,
    -- filter=43 channel=30
    -2, 18, 7, 22, 10, 4, 17, 12, -4,
    -- filter=43 channel=31
    -6, -5, -2, -8, 2, 6, 10, 9, 10,
    -- filter=43 channel=32
    -2, 5, 0, 0, 12, 6, 17, 11, 6,
    -- filter=43 channel=33
    4, -4, 9, -9, -4, 3, -1, 9, -5,
    -- filter=43 channel=34
    6, -1, -5, -1, 0, 1, 10, 7, 7,
    -- filter=43 channel=35
    9, 12, 8, -9, 11, 8, 2, 5, -2,
    -- filter=43 channel=36
    0, 0, -6, 6, -3, 1, 4, -5, 0,
    -- filter=43 channel=37
    4, 19, -1, -3, 21, 3, 11, 1, 7,
    -- filter=43 channel=38
    13, 8, 19, 2, 6, 0, -19, -4, -5,
    -- filter=43 channel=39
    3, 6, 2, 7, 5, -8, -3, 2, 4,
    -- filter=43 channel=40
    -2, 2, 0, -3, -6, -3, 8, -4, 8,
    -- filter=43 channel=41
    15, 23, 21, -8, -13, -10, -13, -23, -12,
    -- filter=43 channel=42
    -6, -5, 6, 6, 2, -5, -10, -6, 7,
    -- filter=43 channel=43
    11, 22, 14, 27, 37, 31, 19, 17, 14,
    -- filter=43 channel=44
    -5, 11, 15, 3, -1, 0, 13, 19, 9,
    -- filter=43 channel=45
    -8, 5, -7, -3, -10, 0, 3, -5, -3,
    -- filter=43 channel=46
    11, 6, 13, 7, 4, -1, -1, 5, 6,
    -- filter=43 channel=47
    1, -8, 0, -4, 0, 4, -9, 5, 9,
    -- filter=43 channel=48
    11, 13, -3, 3, -4, -2, -5, -5, 6,
    -- filter=43 channel=49
    1, 9, 10, -1, -6, -18, -9, -12, -2,
    -- filter=43 channel=50
    9, 4, 18, 17, 10, 13, 6, 0, 6,
    -- filter=43 channel=51
    -6, -11, -11, 6, -12, 4, -5, -12, 1,
    -- filter=43 channel=52
    8, 4, -10, 0, 0, -1, 1, 3, -3,
    -- filter=43 channel=53
    7, 1, 2, 0, 22, 14, 21, 21, 6,
    -- filter=43 channel=54
    12, 8, 18, 2, 18, 9, 0, 4, 7,
    -- filter=43 channel=55
    -8, -2, -9, -3, -1, 5, 9, -1, 1,
    -- filter=43 channel=56
    -5, -6, 5, 13, -6, 3, 11, -7, -8,
    -- filter=43 channel=57
    2, -6, -9, 3, -2, 4, -9, 10, -6,
    -- filter=43 channel=58
    11, -8, 1, 11, 11, 2, 1, 9, 6,
    -- filter=43 channel=59
    19, 14, 16, 3, 3, -4, -6, -13, -9,
    -- filter=43 channel=60
    0, 15, 1, -4, -8, 2, -21, -25, -28,
    -- filter=43 channel=61
    2, 16, 15, -1, -1, -1, -3, -26, -14,
    -- filter=43 channel=62
    0, 12, 18, 4, 7, -1, 3, 4, 0,
    -- filter=43 channel=63
    -6, -4, 0, -7, -3, 5, 4, 2, -5,
    -- filter=44 channel=0
    2, 9, 4, 5, 3, 12, 6, 12, 1,
    -- filter=44 channel=1
    -6, 5, -8, 4, 8, 14, 0, 1, 7,
    -- filter=44 channel=2
    2, 4, 12, 10, 12, 14, 7, 0, 3,
    -- filter=44 channel=3
    1, -5, 8, 4, -2, -7, 3, -5, 5,
    -- filter=44 channel=4
    -12, -6, -8, -8, -4, -4, 5, 12, -6,
    -- filter=44 channel=5
    -12, -12, -6, -6, 2, -9, -13, -12, 4,
    -- filter=44 channel=6
    2, -3, -3, -1, 15, 1, -3, -2, 14,
    -- filter=44 channel=7
    -2, 6, 5, 0, -9, 9, -6, 5, -7,
    -- filter=44 channel=8
    -2, 10, 12, -11, 11, 11, 2, 5, 7,
    -- filter=44 channel=9
    -15, -29, -38, -40, -48, -46, -31, -41, -21,
    -- filter=44 channel=10
    6, 10, -1, -6, 9, 2, 0, 8, 9,
    -- filter=44 channel=11
    -10, -9, -2, 5, -3, -4, -10, 8, 2,
    -- filter=44 channel=12
    9, 0, -6, 0, 10, 9, 8, -9, 5,
    -- filter=44 channel=13
    0, -12, 1, -4, -11, 8, -2, 0, -1,
    -- filter=44 channel=14
    -13, -10, 11, 2, 0, 0, -4, 0, 7,
    -- filter=44 channel=15
    -8, 0, 10, 2, -6, 5, -6, 7, 8,
    -- filter=44 channel=16
    -15, 2, -6, -8, 11, 5, -4, -2, -4,
    -- filter=44 channel=17
    -5, 8, 4, -1, -3, 12, -4, 7, -2,
    -- filter=44 channel=18
    1, 3, -7, 9, 2, 0, -9, -10, 4,
    -- filter=44 channel=19
    -5, -4, 2, -10, 0, -14, -1, -2, 0,
    -- filter=44 channel=20
    4, -12, -5, -6, -13, -6, -3, -11, -9,
    -- filter=44 channel=21
    0, 7, -4, 0, -5, 8, 11, -8, 10,
    -- filter=44 channel=22
    -8, 6, 8, 4, 9, 0, -8, -10, 3,
    -- filter=44 channel=23
    10, 8, 6, -4, 8, 14, 3, 16, 15,
    -- filter=44 channel=24
    -6, -2, -8, -1, 4, -6, -3, 9, -2,
    -- filter=44 channel=25
    -8, 4, 12, 6, 9, 19, 3, 4, 4,
    -- filter=44 channel=26
    -4, -3, 12, 1, -8, 3, -3, 4, 10,
    -- filter=44 channel=27
    0, 5, 0, 8, 2, 18, -5, 5, 6,
    -- filter=44 channel=28
    1, 0, 2, -12, 2, -4, -13, 4, 4,
    -- filter=44 channel=29
    -5, 0, -3, -4, -10, 14, 6, -2, -5,
    -- filter=44 channel=30
    -15, -10, 1, -4, -7, 5, 0, -8, 7,
    -- filter=44 channel=31
    6, -6, 0, 4, 7, -3, 12, 9, 2,
    -- filter=44 channel=32
    -2, -10, 9, -13, 2, 7, 3, 11, 3,
    -- filter=44 channel=33
    -5, 0, 8, -5, -8, -10, -7, 5, -8,
    -- filter=44 channel=34
    7, 1, -3, -6, 1, 6, 4, 6, -3,
    -- filter=44 channel=35
    2, 20, 8, 15, 27, 14, 0, 21, 2,
    -- filter=44 channel=36
    -6, 2, -1, -4, -2, -7, -1, 2, -1,
    -- filter=44 channel=37
    -15, -15, -7, -10, -8, -3, -15, -4, -10,
    -- filter=44 channel=38
    6, -1, 11, 10, 2, 18, 3, 18, 10,
    -- filter=44 channel=39
    5, 0, 10, 8, -3, -6, -8, 4, -1,
    -- filter=44 channel=40
    8, -4, -3, -2, -6, 13, 1, 6, 4,
    -- filter=44 channel=41
    -5, 4, 17, -2, 5, 16, -1, 18, 7,
    -- filter=44 channel=42
    9, 4, 0, -9, 2, 3, 6, 7, 1,
    -- filter=44 channel=43
    0, 8, 1, 10, 15, 9, 14, 2, 17,
    -- filter=44 channel=44
    -4, -10, 8, -5, 8, 1, -1, 1, 5,
    -- filter=44 channel=45
    3, -9, -9, -9, 0, 2, -10, 5, 9,
    -- filter=44 channel=46
    1, 5, 10, -7, 2, -2, 7, 7, 1,
    -- filter=44 channel=47
    -1, 4, 4, 2, 8, -2, -5, -4, -5,
    -- filter=44 channel=48
    6, -5, 9, -8, -3, 3, 4, -4, -11,
    -- filter=44 channel=49
    -7, 19, 12, 5, 19, 17, 0, 13, -1,
    -- filter=44 channel=50
    -5, -6, 4, -11, -8, 13, -6, 1, 6,
    -- filter=44 channel=51
    -7, 17, 7, 0, 6, 5, -1, 10, 15,
    -- filter=44 channel=52
    3, -3, -3, 10, -4, -6, 0, -1, 6,
    -- filter=44 channel=53
    -12, -5, 11, -13, -5, 3, -1, 5, 12,
    -- filter=44 channel=54
    -27, -28, -21, -29, -29, -26, -31, -29, -28,
    -- filter=44 channel=55
    -4, 10, -1, 8, -7, -3, -3, 8, -4,
    -- filter=44 channel=56
    -10, 1, -1, -9, 6, -6, 6, 2, 5,
    -- filter=44 channel=57
    8, 4, -5, 5, 8, 10, -1, 5, -6,
    -- filter=44 channel=58
    11, 4, -7, -6, 10, 9, 0, -4, 8,
    -- filter=44 channel=59
    -6, 4, 0, -2, 10, 19, 1, 8, 5,
    -- filter=44 channel=60
    -5, 7, 9, -10, 5, 11, -6, 8, 15,
    -- filter=44 channel=61
    -7, -4, 0, 4, 12, 12, 0, 18, 14,
    -- filter=44 channel=62
    -12, 4, 1, -5, 7, 6, -2, 9, -2,
    -- filter=44 channel=63
    -4, -1, -8, -3, -9, 2, -1, 3, -9,
    -- filter=45 channel=0
    5, -11, -9, -2, -6, 5, -5, 0, -1,
    -- filter=45 channel=1
    0, 5, 6, 5, 15, 13, 0, 0, 5,
    -- filter=45 channel=2
    11, 19, 13, 13, 5, 12, 6, 1, 8,
    -- filter=45 channel=3
    -1, -3, -9, -7, -2, -10, -8, -7, 6,
    -- filter=45 channel=4
    -10, 3, 7, 2, -11, -1, 9, -1, 6,
    -- filter=45 channel=5
    1, 2, -12, -1, -16, -2, -12, -1, -11,
    -- filter=45 channel=6
    7, 8, 8, 8, 12, 3, -1, -4, 12,
    -- filter=45 channel=7
    0, -5, -6, -4, -8, 4, 4, -4, 0,
    -- filter=45 channel=8
    -5, -12, 0, -1, -1, -4, 1, -7, 2,
    -- filter=45 channel=9
    13, 18, 8, 4, 5, 1, 10, 0, -1,
    -- filter=45 channel=10
    0, 1, 0, 6, 6, -6, -3, 6, -1,
    -- filter=45 channel=11
    1, 1, -4, -6, 3, 2, 7, 5, -2,
    -- filter=45 channel=12
    -3, -8, 0, -3, 9, 0, -5, -6, -1,
    -- filter=45 channel=13
    -1, -5, -8, 5, -7, 0, 10, 9, 6,
    -- filter=45 channel=14
    3, 0, 6, 0, -17, -11, -11, -1, -10,
    -- filter=45 channel=15
    3, -10, 0, 3, 5, -5, 4, -7, -9,
    -- filter=45 channel=16
    -1, 8, 4, -1, 11, 1, 3, 2, 4,
    -- filter=45 channel=17
    -2, -2, -8, -10, -14, 5, -10, -11, -1,
    -- filter=45 channel=18
    -1, 4, 13, 5, 0, 3, 14, -1, 8,
    -- filter=45 channel=19
    5, -2, 4, -2, 6, 1, 10, 0, 15,
    -- filter=45 channel=20
    5, 0, -1, 4, -3, 7, 0, 2, 3,
    -- filter=45 channel=21
    7, 11, 9, 6, -1, 3, -5, -8, 4,
    -- filter=45 channel=22
    -8, 3, 8, -5, -2, 7, -6, 0, 8,
    -- filter=45 channel=23
    4, 13, 12, 2, -5, 11, -5, 3, 13,
    -- filter=45 channel=24
    -10, -4, 0, -1, -9, 7, -9, -4, -4,
    -- filter=45 channel=25
    4, 15, 10, 7, 22, 9, 12, 5, 0,
    -- filter=45 channel=26
    -5, -11, -6, 6, -12, -7, -5, -5, 3,
    -- filter=45 channel=27
    -3, 13, 7, 9, -1, 11, 4, 6, -4,
    -- filter=45 channel=28
    9, 3, 4, -4, -9, 5, 9, 8, 5,
    -- filter=45 channel=29
    9, 9, -10, -8, -9, 6, 4, -1, 8,
    -- filter=45 channel=30
    -24, -21, -7, -25, -13, -15, -27, -29, -12,
    -- filter=45 channel=31
    7, 4, -8, 10, 1, -8, 9, -4, 7,
    -- filter=45 channel=32
    11, -1, 13, -3, -1, 7, 8, 2, 11,
    -- filter=45 channel=33
    4, -1, -1, -5, -2, 1, 2, 5, -5,
    -- filter=45 channel=34
    -6, -1, -3, 5, -3, -11, -3, -9, -10,
    -- filter=45 channel=35
    8, 5, 5, -4, 1, 3, 8, -1, 10,
    -- filter=45 channel=36
    -6, 5, -7, 12, 4, 6, 8, 3, 11,
    -- filter=45 channel=37
    3, 8, 5, -1, 0, -11, -13, -6, -7,
    -- filter=45 channel=38
    5, 10, 1, -1, 6, 2, 6, -1, -3,
    -- filter=45 channel=39
    -1, 5, -4, 6, -8, -3, 2, 3, -3,
    -- filter=45 channel=40
    -2, -9, -4, -11, 3, 9, -3, 9, -5,
    -- filter=45 channel=41
    -10, -10, -8, -13, -2, -5, -6, 1, -6,
    -- filter=45 channel=42
    5, -3, 3, 0, 5, 1, 7, 6, 10,
    -- filter=45 channel=43
    7, -5, 1, 5, -4, -2, 5, -1, 8,
    -- filter=45 channel=44
    4, -7, 8, 2, 3, -7, 10, 8, -4,
    -- filter=45 channel=45
    -4, 7, 5, -6, 0, -5, -8, -5, -4,
    -- filter=45 channel=46
    -14, -13, -10, -14, -12, -3, -7, -8, -3,
    -- filter=45 channel=47
    -2, -3, -2, 4, 3, 0, -4, 6, -2,
    -- filter=45 channel=48
    -1, 0, 10, -5, -4, 9, 9, 9, -5,
    -- filter=45 channel=49
    -2, 0, -2, -5, 11, 6, 7, 12, 6,
    -- filter=45 channel=50
    -9, -7, -11, -7, -10, 5, -9, -1, -12,
    -- filter=45 channel=51
    3, 3, 10, 9, 11, -1, 2, 10, -7,
    -- filter=45 channel=52
    -7, -7, -1, -10, 6, -1, -8, -5, 0,
    -- filter=45 channel=53
    1, -11, 0, -4, -2, -7, -1, -17, 1,
    -- filter=45 channel=54
    6, 7, 10, -14, -5, 2, -9, -11, 0,
    -- filter=45 channel=55
    4, 3, 2, 1, 4, -8, -6, -6, 8,
    -- filter=45 channel=56
    -4, -9, 7, -8, 0, -1, 5, 5, -11,
    -- filter=45 channel=57
    -3, -1, -5, -6, 3, 1, -1, 5, -7,
    -- filter=45 channel=58
    8, 11, -2, 5, 2, 12, 6, 8, 8,
    -- filter=45 channel=59
    7, 9, 4, -6, -4, -3, 4, 11, 7,
    -- filter=45 channel=60
    -8, 0, -15, -1, -6, -7, -4, -14, -1,
    -- filter=45 channel=61
    -5, -3, -7, -5, 1, -2, -15, -5, 7,
    -- filter=45 channel=62
    5, -6, -5, 1, 3, 0, -12, -12, 8,
    -- filter=45 channel=63
    6, 0, 7, 10, 4, -1, -3, 2, -6,
    -- filter=46 channel=0
    3, -9, -3, 1, -10, -5, 3, -6, 1,
    -- filter=46 channel=1
    3, -3, 3, 8, 0, 9, -2, 4, 8,
    -- filter=46 channel=2
    0, -10, 0, 1, -8, 12, 3, 8, 8,
    -- filter=46 channel=3
    -6, -7, 7, 10, -6, -7, -6, 1, -2,
    -- filter=46 channel=4
    12, 9, 4, 11, -1, 7, -5, 0, 4,
    -- filter=46 channel=5
    5, -6, 9, -4, -6, -10, 1, -1, 2,
    -- filter=46 channel=6
    2, 5, 6, 2, -6, 6, 6, 0, -6,
    -- filter=46 channel=7
    6, 8, 0, -7, 10, 9, -7, 5, -3,
    -- filter=46 channel=8
    1, -8, 2, 8, -7, -12, 6, 3, -4,
    -- filter=46 channel=9
    -2, 5, -10, 0, -8, -5, 12, -3, 0,
    -- filter=46 channel=10
    -2, -4, -4, -7, 11, 6, -3, 1, 8,
    -- filter=46 channel=11
    6, -9, -10, -2, 8, -11, 10, 3, 0,
    -- filter=46 channel=12
    -10, 5, -8, 0, 5, -2, 9, -6, -10,
    -- filter=46 channel=13
    -3, -5, -7, -1, 0, -7, 0, 0, -8,
    -- filter=46 channel=14
    -8, -7, -8, 0, 5, 2, -1, 7, -3,
    -- filter=46 channel=15
    -7, -9, 8, 2, -10, -11, 6, -2, 6,
    -- filter=46 channel=16
    -5, 3, 3, 9, -7, -3, 12, -6, 6,
    -- filter=46 channel=17
    4, -9, -8, 4, 6, -13, 2, 8, 3,
    -- filter=46 channel=18
    -1, -4, -9, -6, -7, 4, 10, 4, 0,
    -- filter=46 channel=19
    -4, -8, 0, 9, -4, 5, 14, 1, 7,
    -- filter=46 channel=20
    -4, -8, 3, -2, -6, -1, 6, 8, 13,
    -- filter=46 channel=21
    -5, -7, -6, 0, 10, 2, -6, 4, -5,
    -- filter=46 channel=22
    9, 1, 8, -2, 7, 8, 2, 9, -8,
    -- filter=46 channel=23
    4, 6, 3, 8, 4, -8, 0, -5, -3,
    -- filter=46 channel=24
    -2, 9, -8, -1, -6, 0, 6, -6, 7,
    -- filter=46 channel=25
    9, 1, 3, -1, 0, 0, 1, -8, -4,
    -- filter=46 channel=26
    8, 6, 14, -6, 1, 10, 6, 4, -6,
    -- filter=46 channel=27
    0, -12, 3, 0, 3, 0, -4, -3, -1,
    -- filter=46 channel=28
    14, -2, 3, 6, 3, 0, 9, 4, -2,
    -- filter=46 channel=29
    11, 3, 4, -3, -13, -2, -1, -11, 0,
    -- filter=46 channel=30
    15, 15, 6, 10, 19, -6, 5, 4, 1,
    -- filter=46 channel=31
    0, -8, 4, -3, 3, 4, -6, 8, -6,
    -- filter=46 channel=32
    -9, 0, 10, 9, 3, 10, 0, 1, 10,
    -- filter=46 channel=33
    -10, 1, 1, -4, -6, -6, 2, 2, 7,
    -- filter=46 channel=34
    -9, -4, 9, 1, 10, -5, -5, 10, -2,
    -- filter=46 channel=35
    -4, -9, -6, 3, 0, 0, 3, -6, -4,
    -- filter=46 channel=36
    -5, 5, 4, 4, -8, -4, -5, 8, 6,
    -- filter=46 channel=37
    6, -8, 9, 9, 9, 0, -1, 7, -4,
    -- filter=46 channel=38
    10, -4, 10, -3, -4, 1, -3, 1, 3,
    -- filter=46 channel=39
    0, 5, 6, -8, 9, -1, -3, 8, 0,
    -- filter=46 channel=40
    0, -7, -6, -1, 3, 5, 1, 1, -10,
    -- filter=46 channel=41
    -3, 1, -4, 11, -5, 3, -4, -8, -4,
    -- filter=46 channel=42
    8, -9, -1, 8, -8, -1, 10, 10, 4,
    -- filter=46 channel=43
    5, 12, 13, -6, 8, -4, 3, 9, -5,
    -- filter=46 channel=44
    7, 0, 10, -3, 13, 9, 9, 10, 0,
    -- filter=46 channel=45
    6, 2, 3, 4, -10, -5, 4, -1, -3,
    -- filter=46 channel=46
    -8, 7, 12, 8, 5, -6, 0, 8, 1,
    -- filter=46 channel=47
    -7, 8, -1, 3, 3, 2, 8, 0, 4,
    -- filter=46 channel=48
    -9, 0, 3, -3, -8, 9, -7, -5, -3,
    -- filter=46 channel=49
    9, -7, -6, -1, 0, 5, 10, 7, 4,
    -- filter=46 channel=50
    -3, 16, 7, 5, 6, -2, 16, 15, -9,
    -- filter=46 channel=51
    7, -7, 3, 7, -5, 0, -8, 8, -8,
    -- filter=46 channel=52
    0, 6, -9, -9, 4, 7, -7, 9, 1,
    -- filter=46 channel=53
    11, 11, 0, 15, 0, 5, 2, 2, 0,
    -- filter=46 channel=54
    -2, -7, -6, 12, 6, -12, 0, -10, -3,
    -- filter=46 channel=55
    -1, -1, -8, 0, 6, 1, 9, 10, -10,
    -- filter=46 channel=56
    4, -2, 11, 10, 3, 0, 9, -3, -7,
    -- filter=46 channel=57
    -7, -10, 9, 0, 9, -9, -7, 2, -3,
    -- filter=46 channel=58
    -8, 2, 12, -7, 4, -2, 5, 3, 2,
    -- filter=46 channel=59
    0, 1, -3, -4, -1, 2, 0, -1, 4,
    -- filter=46 channel=60
    -7, -2, 4, 13, -5, -3, -3, -10, 7,
    -- filter=46 channel=61
    -6, 2, 2, -2, -5, 4, 10, 5, -8,
    -- filter=46 channel=62
    -2, 0, 9, -2, -4, -8, 11, 7, -8,
    -- filter=46 channel=63
    -6, 7, 6, -7, 9, 6, -10, 6, -2,
    -- filter=47 channel=0
    13, 23, 15, 7, 33, 12, 4, 22, 15,
    -- filter=47 channel=1
    -18, -3, -10, -3, 0, 3, -12, -1, 1,
    -- filter=47 channel=2
    -8, -7, -2, -2, -7, -14, -22, -21, -14,
    -- filter=47 channel=3
    -13, -11, 6, -10, -4, 0, -12, -3, 7,
    -- filter=47 channel=4
    1, 12, -3, 19, 8, 10, 0, -1, 3,
    -- filter=47 channel=5
    2, -16, -1, -5, -15, -1, -2, -11, 2,
    -- filter=47 channel=6
    8, 8, 1, -6, -1, 0, -2, 4, 5,
    -- filter=47 channel=7
    -3, -5, -5, -13, 1, 2, 0, -2, 9,
    -- filter=47 channel=8
    17, 4, 0, 14, 17, 0, 9, 16, 0,
    -- filter=47 channel=9
    -12, -44, -33, -21, -54, -30, -19, -40, -36,
    -- filter=47 channel=10
    7, 12, 3, 15, 27, 17, 14, 7, 19,
    -- filter=47 channel=11
    1, 10, -4, 4, 4, 3, 10, 3, -4,
    -- filter=47 channel=12
    7, 4, 0, 7, 5, -5, -8, 10, 5,
    -- filter=47 channel=13
    -7, -5, -11, 5, -1, -4, 7, -7, -9,
    -- filter=47 channel=14
    -13, -10, -7, -14, 1, -7, -11, -2, -7,
    -- filter=47 channel=15
    9, 3, -4, 7, 6, 9, -7, 1, 0,
    -- filter=47 channel=16
    1, 0, -4, 2, -12, -1, 0, -2, -3,
    -- filter=47 channel=17
    5, 15, 13, 5, 21, 17, 2, 12, 13,
    -- filter=47 channel=18
    9, 10, -2, 23, 7, 0, 14, 6, 3,
    -- filter=47 channel=19
    -21, -21, -12, -16, -19, -9, -18, -10, -7,
    -- filter=47 channel=20
    -11, 0, -10, -19, -19, -18, -4, -15, -9,
    -- filter=47 channel=21
    -2, 1, -1, -6, -1, -8, 6, -2, 12,
    -- filter=47 channel=22
    -7, 6, 4, -4, 0, 6, -3, -5, 0,
    -- filter=47 channel=23
    2, 9, 7, 9, 16, 13, 9, 14, 17,
    -- filter=47 channel=24
    -8, 0, 5, -1, 5, 9, 11, 13, 3,
    -- filter=47 channel=25
    -20, -16, -3, -18, -7, -12, -4, -6, -4,
    -- filter=47 channel=26
    -14, -11, -8, -1, -1, 8, -11, -11, 4,
    -- filter=47 channel=27
    -1, 1, 7, -4, 22, 12, -4, 9, -2,
    -- filter=47 channel=28
    1, -6, -15, 9, -15, 0, 7, -16, -12,
    -- filter=47 channel=29
    -8, -10, 0, -2, -7, -9, -18, -21, -17,
    -- filter=47 channel=30
    -22, -2, 7, -14, -3, 7, -27, -10, 4,
    -- filter=47 channel=31
    -4, 13, 1, -6, 12, -7, 14, 10, 12,
    -- filter=47 channel=32
    -8, 8, -3, -17, -8, 14, -5, -2, 5,
    -- filter=47 channel=33
    0, -1, 10, 2, 7, 10, -10, -4, 5,
    -- filter=47 channel=34
    -14, 5, 0, 5, -7, -8, 3, 0, 3,
    -- filter=47 channel=35
    13, 14, 20, 6, 24, 26, 10, 27, 11,
    -- filter=47 channel=36
    4, 11, 2, -6, 5, 12, -8, -4, -4,
    -- filter=47 channel=37
    -4, -22, -19, -11, -21, -11, -3, -14, -9,
    -- filter=47 channel=38
    2, -2, -5, 11, 20, 20, -6, 0, -6,
    -- filter=47 channel=39
    -9, -6, 0, -8, 0, 1, -6, -2, 3,
    -- filter=47 channel=40
    -4, 11, 4, 8, 9, -3, -11, -6, -1,
    -- filter=47 channel=41
    14, 15, 17, 9, 14, 8, 7, 6, 14,
    -- filter=47 channel=42
    0, -6, -5, 9, 10, 7, -9, 5, 4,
    -- filter=47 channel=43
    -24, -12, -7, 1, 7, 8, -8, 7, 17,
    -- filter=47 channel=44
    4, 3, 1, -3, -6, 0, -11, -6, -3,
    -- filter=47 channel=45
    10, 9, -8, 0, 9, 7, 0, 1, -5,
    -- filter=47 channel=46
    -6, -12, -2, -8, -12, -7, -6, -4, -3,
    -- filter=47 channel=47
    9, -8, -10, 0, 7, -9, -7, 4, 9,
    -- filter=47 channel=48
    -6, -13, -11, 0, -18, 3, 0, -15, -15,
    -- filter=47 channel=49
    17, 34, 12, 22, 28, 22, 1, 7, 18,
    -- filter=47 channel=50
    -10, -2, -5, -21, -4, 5, -13, -13, 12,
    -- filter=47 channel=51
    16, 26, 14, 27, 28, 19, 9, 29, 26,
    -- filter=47 channel=52
    -9, -4, 6, 6, 8, 10, 0, -6, 4,
    -- filter=47 channel=53
    -17, -2, 7, -15, -17, 2, -7, -3, -3,
    -- filter=47 channel=54
    -17, -31, -16, -14, -38, -37, -23, -29, -24,
    -- filter=47 channel=55
    -8, 2, 0, -5, -5, 7, 2, -6, -4,
    -- filter=47 channel=56
    -4, -3, 7, -11, -4, -2, -4, -9, 7,
    -- filter=47 channel=57
    6, 8, 0, 9, -8, -1, -8, -2, 4,
    -- filter=47 channel=58
    -2, 7, 3, -8, -8, 9, 9, -3, 4,
    -- filter=47 channel=59
    -6, 3, 9, 0, 3, -1, 4, 8, 6,
    -- filter=47 channel=60
    10, 14, 10, 17, 24, 12, 12, 5, 2,
    -- filter=47 channel=61
    4, 18, 15, 22, 19, 15, 0, 26, 19,
    -- filter=47 channel=62
    -3, -2, -2, -4, -9, -6, 0, -6, -7,
    -- filter=47 channel=63
    -10, -7, 0, 9, 1, -6, 6, -9, -10,
    -- filter=48 channel=0
    -13, -6, 0, -2, 1, 15, 0, 8, 15,
    -- filter=48 channel=1
    0, -3, -9, -7, -12, -3, 10, -3, -6,
    -- filter=48 channel=2
    0, -13, -6, 8, -2, 8, -6, 0, -7,
    -- filter=48 channel=3
    -8, 2, 3, 7, 13, 0, 0, 0, 10,
    -- filter=48 channel=4
    -11, -8, -2, 4, 6, -4, 6, 14, 8,
    -- filter=48 channel=5
    2, -17, -8, -1, 3, -5, 0, -13, -12,
    -- filter=48 channel=6
    -1, -12, -3, 3, 7, 13, 4, 1, 6,
    -- filter=48 channel=7
    1, 0, 0, -2, -4, 0, -4, -10, 3,
    -- filter=48 channel=8
    -2, -10, -9, 5, 17, 14, 15, 24, 0,
    -- filter=48 channel=9
    -11, -19, -28, -27, -33, -34, -21, -39, -38,
    -- filter=48 channel=10
    1, 3, 9, -15, 3, 5, 5, 8, 11,
    -- filter=48 channel=11
    -5, -11, 3, 3, -5, 14, 9, 13, 20,
    -- filter=48 channel=12
    -6, 5, 0, -8, -1, 3, 0, 5, -2,
    -- filter=48 channel=13
    -14, -17, -8, 7, -6, -2, 12, -2, -5,
    -- filter=48 channel=14
    -12, -4, -8, -13, -11, 3, -4, -10, -6,
    -- filter=48 channel=15
    -2, -18, -15, 19, 14, 13, 0, 6, -2,
    -- filter=48 channel=16
    -19, -25, -19, 11, 12, 12, 22, 16, -4,
    -- filter=48 channel=17
    -6, -18, 2, -1, 10, 9, 18, 6, 3,
    -- filter=48 channel=18
    -4, 10, -2, 0, 5, -3, 4, 6, -4,
    -- filter=48 channel=19
    -9, -9, -3, -10, -8, -2, 4, -1, -10,
    -- filter=48 channel=20
    -13, -1, -13, -8, -4, -2, -3, -7, -15,
    -- filter=48 channel=21
    12, -7, 5, -1, 10, 6, -1, -8, 11,
    -- filter=48 channel=22
    -7, 3, -1, 5, 7, 1, 3, 4, 4,
    -- filter=48 channel=23
    -9, 8, 1, -4, 6, 19, 8, 14, 19,
    -- filter=48 channel=24
    -2, -18, -14, 7, -6, 7, 16, 9, 11,
    -- filter=48 channel=25
    -13, -12, -5, 0, 8, 5, 5, 5, 8,
    -- filter=48 channel=26
    -4, -9, 0, -7, -8, -7, -7, -10, 5,
    -- filter=48 channel=27
    2, 5, -12, 7, 14, 8, 2, 10, 17,
    -- filter=48 channel=28
    -11, -5, -10, 15, 11, 7, 9, -2, -11,
    -- filter=48 channel=29
    -8, -24, -9, 13, 10, 7, 24, 7, 2,
    -- filter=48 channel=30
    -8, -11, -7, -7, -23, -15, -23, -22, 2,
    -- filter=48 channel=31
    4, -3, 5, 3, 9, 2, 8, 0, -5,
    -- filter=48 channel=32
    -15, -6, -4, -6, -13, 3, -13, 0, 11,
    -- filter=48 channel=33
    -8, -1, -2, -9, -10, -10, 10, -4, -7,
    -- filter=48 channel=34
    -4, -5, -6, 1, -6, 1, -2, -14, 0,
    -- filter=48 channel=35
    -9, 12, 0, -5, 10, 13, 4, 9, 7,
    -- filter=48 channel=36
    8, 7, 9, -6, -9, -10, 1, 0, 10,
    -- filter=48 channel=37
    -16, -20, -1, 3, -1, -9, -8, 2, -2,
    -- filter=48 channel=38
    -12, -3, -7, 0, 5, 9, 22, 26, 17,
    -- filter=48 channel=39
    -9, -5, 4, 4, 0, 10, -6, -8, -3,
    -- filter=48 channel=40
    6, -1, -7, 10, 5, -2, 0, 2, 8,
    -- filter=48 channel=41
    -9, -5, 0, 21, 24, 27, 26, 11, 9,
    -- filter=48 channel=42
    5, -4, 0, 0, -2, -7, 1, -6, 7,
    -- filter=48 channel=43
    -4, -21, -3, -28, -25, -16, 4, -2, 0,
    -- filter=48 channel=44
    1, -14, 8, -9, 1, 0, -3, -9, 0,
    -- filter=48 channel=45
    -9, 9, -7, 2, 0, 5, 0, -2, 9,
    -- filter=48 channel=46
    2, -10, 5, -13, 4, -3, -7, 0, -13,
    -- filter=48 channel=47
    1, -5, -2, -7, 4, -7, 1, -9, -4,
    -- filter=48 channel=48
    -14, -15, -1, -4, 0, 0, 1, -5, -11,
    -- filter=48 channel=49
    -2, 11, 2, 7, 23, 27, -1, 4, 10,
    -- filter=48 channel=50
    -5, -15, -9, -15, -29, -10, -8, -12, -5,
    -- filter=48 channel=51
    7, 14, 2, -8, 6, 18, -5, 5, 20,
    -- filter=48 channel=52
    -7, 11, -6, 5, -3, 1, 0, 2, -8,
    -- filter=48 channel=53
    -13, -7, -3, -6, -5, -14, -5, -16, 7,
    -- filter=48 channel=54
    -7, -31, -23, -9, -20, -30, -9, -22, -30,
    -- filter=48 channel=55
    -9, -7, -2, -5, -8, 7, -1, 10, 5,
    -- filter=48 channel=56
    -2, 0, 6, -6, -1, -8, 8, -1, 1,
    -- filter=48 channel=57
    -6, 0, 6, 5, 2, 3, 5, -8, 3,
    -- filter=48 channel=58
    6, 11, 7, 0, 7, -4, -4, 3, -10,
    -- filter=48 channel=59
    -9, 5, -6, 15, 15, 6, 9, 7, 2,
    -- filter=48 channel=60
    -9, -17, -21, 13, 11, 11, 19, 27, 9,
    -- filter=48 channel=61
    -19, -8, -15, -1, 21, 22, 17, 33, 24,
    -- filter=48 channel=62
    -2, -9, -1, 7, 1, 8, 9, 13, 9,
    -- filter=48 channel=63
    1, 1, 9, -7, 4, 10, -7, 0, 8,
    -- filter=49 channel=0
    2, -1, -6, -11, 2, -8, 6, -11, -11,
    -- filter=49 channel=1
    0, 6, 9, 1, 5, 0, 0, 15, 7,
    -- filter=49 channel=2
    -13, 5, -6, 4, 9, 16, 4, 12, 21,
    -- filter=49 channel=3
    -6, 10, 1, 2, 21, 10, 16, 12, 19,
    -- filter=49 channel=4
    2, -17, -13, -5, 0, 4, -6, -4, 6,
    -- filter=49 channel=5
    4, 3, 5, 15, 3, 10, 0, -3, 2,
    -- filter=49 channel=6
    -2, -12, -1, -8, 2, 4, -8, 6, -4,
    -- filter=49 channel=7
    0, -8, -12, -5, -2, 8, -8, 4, -4,
    -- filter=49 channel=8
    -23, -23, -22, -6, -7, 9, 6, 10, 14,
    -- filter=49 channel=9
    0, 15, 14, -7, 12, 20, 14, 14, 24,
    -- filter=49 channel=10
    0, -12, 0, 0, 1, -18, -8, -3, -6,
    -- filter=49 channel=11
    -13, -11, -9, -2, -9, 0, 11, 3, 2,
    -- filter=49 channel=12
    -6, -6, 5, 1, 7, -7, -4, 0, -4,
    -- filter=49 channel=13
    -19, -2, -4, -2, -1, -12, 14, 17, 7,
    -- filter=49 channel=14
    5, 3, -6, -11, 5, -7, 8, -5, 0,
    -- filter=49 channel=15
    -23, -7, -24, -7, 3, 6, -2, 16, -1,
    -- filter=49 channel=16
    -16, -10, -28, 13, 5, 15, 22, 15, 27,
    -- filter=49 channel=17
    0, -4, -24, -1, 6, 2, 15, 11, 16,
    -- filter=49 channel=18
    -1, -10, -15, 8, -2, -3, 7, 5, -14,
    -- filter=49 channel=19
    13, 15, 9, 7, 16, 13, 1, 16, 14,
    -- filter=49 channel=20
    -9, 4, 0, -8, 11, -9, 2, 0, -10,
    -- filter=49 channel=21
    12, -7, 1, 6, -5, 3, 1, 0, -1,
    -- filter=49 channel=22
    -4, -4, -3, -10, 1, 7, 8, 2, 9,
    -- filter=49 channel=23
    4, -10, -10, -4, -18, -11, 5, 0, 1,
    -- filter=49 channel=24
    -10, -1, -4, 2, -15, -9, 5, 0, 11,
    -- filter=49 channel=25
    -12, -6, 1, 13, 22, 23, 7, 26, 21,
    -- filter=49 channel=26
    -13, 0, -1, 1, 1, -5, -3, 5, 6,
    -- filter=49 channel=27
    3, -10, -15, -4, 9, 11, 18, 8, 15,
    -- filter=49 channel=28
    -9, 0, -11, 7, 16, 10, -2, 7, 21,
    -- filter=49 channel=29
    -12, -22, -21, 0, 1, 13, 25, 17, 25,
    -- filter=49 channel=30
    0, -4, -17, -2, -14, -8, -9, -1, -7,
    -- filter=49 channel=31
    13, 6, 11, 10, 9, -9, 8, 7, -8,
    -- filter=49 channel=32
    5, 4, 7, -6, -1, -7, 1, 3, 10,
    -- filter=49 channel=33
    -8, 6, 6, -6, 8, 8, 10, -2, 7,
    -- filter=49 channel=34
    -9, -8, -3, -6, -5, -2, -4, -6, 0,
    -- filter=49 channel=35
    -5, -4, -10, 2, 8, 9, 0, -3, -3,
    -- filter=49 channel=36
    -2, 9, 6, -7, 4, 7, -7, -6, 0,
    -- filter=49 channel=37
    4, 3, 8, 8, 4, 0, 2, 6, 4,
    -- filter=49 channel=38
    -19, -15, -16, -5, -10, -4, 14, 16, 13,
    -- filter=49 channel=39
    2, -6, 4, 1, -6, 0, 9, 8, 7,
    -- filter=49 channel=40
    9, -2, 7, -7, 0, 13, 0, 0, 0,
    -- filter=49 channel=41
    -1, -9, -28, 4, 15, -1, 4, 17, 1,
    -- filter=49 channel=42
    0, -1, -2, 3, -5, -8, 3, 5, 5,
    -- filter=49 channel=43
    4, 4, -1, -3, -12, 1, 0, 11, 5,
    -- filter=49 channel=44
    -4, 0, -6, 10, 14, 14, -6, 10, 13,
    -- filter=49 channel=45
    2, -4, -3, 0, 7, -2, 5, -6, 0,
    -- filter=49 channel=46
    -7, -4, -1, 4, -7, 3, -8, 3, -6,
    -- filter=49 channel=47
    -9, 8, -8, -8, -4, 0, 4, 6, -2,
    -- filter=49 channel=48
    2, -7, -14, 1, 1, 12, -6, 0, 7,
    -- filter=49 channel=49
    -9, -13, -14, -5, -5, 2, -1, -12, 3,
    -- filter=49 channel=50
    9, -10, -12, 6, -10, -12, 0, 2, 4,
    -- filter=49 channel=51
    1, -7, -3, -16, -12, -5, 0, -15, -13,
    -- filter=49 channel=52
    -4, -4, 7, 8, 0, 2, 3, -7, 5,
    -- filter=49 channel=53
    5, 3, -9, -12, -2, -9, 0, -10, -6,
    -- filter=49 channel=54
    -7, 2, 0, 2, 21, 24, 8, 16, 10,
    -- filter=49 channel=55
    4, -1, 0, -1, -2, 7, -7, -6, -5,
    -- filter=49 channel=56
    -6, -9, 3, 6, -9, -1, -7, 4, 3,
    -- filter=49 channel=57
    1, 9, -2, 5, 6, -3, 4, 0, 0,
    -- filter=49 channel=58
    -4, 3, 8, 4, 14, 5, 1, 11, 8,
    -- filter=49 channel=59
    -4, -3, 0, 17, 9, 16, 14, 25, 13,
    -- filter=49 channel=60
    -13, -30, -36, 2, 2, -12, 17, 13, 12,
    -- filter=49 channel=61
    -1, -18, -30, -2, -17, -16, -1, -2, 9,
    -- filter=49 channel=62
    -7, -7, 2, 1, 1, 0, 9, 9, 15,
    -- filter=49 channel=63
    -6, 4, 7, 10, -6, -3, -2, 5, 2,
    -- filter=50 channel=0
    -8, -2, 9, 0, -6, 0, -17, 6, 3,
    -- filter=50 channel=1
    2, 0, 8, 12, -3, -4, 7, -2, 13,
    -- filter=50 channel=2
    16, 7, -2, 12, 9, 15, -5, 0, -2,
    -- filter=50 channel=3
    -5, 7, 6, -6, 12, -9, -12, 9, 3,
    -- filter=50 channel=4
    1, -11, 8, -8, -4, 6, -14, 7, -7,
    -- filter=50 channel=5
    9, 2, 8, -4, -4, 0, -5, -10, -7,
    -- filter=50 channel=6
    0, -5, 10, -4, 4, 5, 0, -7, 0,
    -- filter=50 channel=7
    6, 4, -15, -6, -2, -16, 0, -4, -14,
    -- filter=50 channel=8
    -8, 0, 11, -12, 13, 2, -15, -8, 15,
    -- filter=50 channel=9
    2, 3, -10, 2, 5, -8, 6, -5, -7,
    -- filter=50 channel=10
    -8, 2, -4, -8, -8, -9, 5, 6, 8,
    -- filter=50 channel=11
    -1, -5, -5, 7, 10, 7, -3, 1, 1,
    -- filter=50 channel=12
    0, 6, 8, 4, 3, 10, -8, 0, -6,
    -- filter=50 channel=13
    -1, -6, 6, 11, 11, -2, -8, 3, 0,
    -- filter=50 channel=14
    -10, -1, -2, -5, 0, -8, 0, -17, -14,
    -- filter=50 channel=15
    -3, 2, 11, 0, -2, 21, -14, -4, 14,
    -- filter=50 channel=16
    17, 8, 5, 14, 21, 8, 0, 3, 6,
    -- filter=50 channel=17
    5, -7, 6, -8, 9, 8, -16, -7, -1,
    -- filter=50 channel=18
    -4, -1, -5, 1, 0, 10, -11, -1, 13,
    -- filter=50 channel=19
    17, -6, -6, 12, 0, -6, 14, 3, 5,
    -- filter=50 channel=20
    2, -13, -18, 2, -15, -8, -4, -12, -16,
    -- filter=50 channel=21
    -1, -4, -3, 8, -5, 1, 6, 2, 0,
    -- filter=50 channel=22
    3, 0, -4, -10, 5, -6, -6, 0, -2,
    -- filter=50 channel=23
    2, -11, 11, -9, 3, 0, 3, -4, 13,
    -- filter=50 channel=24
    2, 3, -2, -8, 0, 8, -3, 3, 13,
    -- filter=50 channel=25
    10, 1, 15, 14, 11, 15, 9, 12, 7,
    -- filter=50 channel=26
    -10, -8, -11, -7, -11, -9, 3, 3, -3,
    -- filter=50 channel=27
    5, -4, 6, 1, 9, 8, -8, -3, 0,
    -- filter=50 channel=28
    7, 1, 16, 7, 13, 6, 0, 0, 11,
    -- filter=50 channel=29
    -4, 5, 2, 14, 6, 9, 3, 1, 13,
    -- filter=50 channel=30
    -10, -26, -15, -20, -30, -26, -26, -24, -19,
    -- filter=50 channel=31
    -2, -1, 4, -10, -8, 1, -8, 10, 2,
    -- filter=50 channel=32
    6, -4, 2, -12, 0, -11, 0, -10, -8,
    -- filter=50 channel=33
    8, 8, 10, 0, -6, 7, 8, -8, 2,
    -- filter=50 channel=34
    -12, 0, -14, 4, 0, 1, 1, 3, -11,
    -- filter=50 channel=35
    -2, 1, -4, 1, 2, 1, -2, -3, 3,
    -- filter=50 channel=36
    8, 8, -1, 3, -6, -1, -7, 0, -5,
    -- filter=50 channel=37
    -8, -5, 2, 1, 7, -11, -1, -7, 0,
    -- filter=50 channel=38
    -4, 4, 2, 0, 13, 14, -9, 0, 15,
    -- filter=50 channel=39
    -5, -2, -8, 6, 3, 5, 0, -7, 3,
    -- filter=50 channel=40
    -8, 3, -8, -12, 3, -6, -1, -12, 1,
    -- filter=50 channel=41
    -3, -8, 14, -8, 16, 14, -12, -7, 13,
    -- filter=50 channel=42
    -4, 7, 3, 2, -5, -5, -10, -6, 4,
    -- filter=50 channel=43
    -16, -23, -16, 5, -17, -9, 5, -1, -6,
    -- filter=50 channel=44
    3, 2, -3, 6, 5, 0, 2, -15, -7,
    -- filter=50 channel=45
    -9, -5, -6, 1, 7, -7, -9, -1, 0,
    -- filter=50 channel=46
    -17, 0, -13, -1, 0, -19, -15, -10, -16,
    -- filter=50 channel=47
    5, -6, 10, -8, -2, 8, 0, 5, -6,
    -- filter=50 channel=48
    -4, -1, -6, 9, 13, 2, 5, 3, 6,
    -- filter=50 channel=49
    1, 3, 11, -8, 9, 6, -11, -3, -4,
    -- filter=50 channel=50
    -4, -26, -6, -17, -26, -8, 2, -16, -9,
    -- filter=50 channel=51
    2, 0, 9, -2, -1, -4, -14, -2, 8,
    -- filter=50 channel=52
    5, -8, 9, 7, 6, 3, 11, 2, -6,
    -- filter=50 channel=53
    -16, -26, -19, -6, -27, -5, -22, -27, -6,
    -- filter=50 channel=54
    -3, 0, -17, -13, -16, -15, 0, -16, -16,
    -- filter=50 channel=55
    -2, 2, -2, -3, 5, -9, 2, 3, 0,
    -- filter=50 channel=56
    2, 0, -2, -11, -11, -9, 0, 2, 3,
    -- filter=50 channel=57
    -3, -5, -3, -2, 0, -8, 4, -1, -5,
    -- filter=50 channel=58
    -3, 12, -5, 0, 9, -2, 1, 9, 2,
    -- filter=50 channel=59
    6, -4, -9, 0, 5, 2, -4, -7, 4,
    -- filter=50 channel=60
    -8, 6, 14, 0, 8, 15, -16, 2, 13,
    -- filter=50 channel=61
    -3, 0, 12, 1, 3, 7, -11, -8, 4,
    -- filter=50 channel=62
    -4, -11, 2, -7, 9, 4, -13, 3, 2,
    -- filter=50 channel=63
    -7, -3, -1, -6, 5, 0, -6, 2, 0,
    -- filter=51 channel=0
    -8, -2, 8, -10, -5, -5, -7, -2, -10,
    -- filter=51 channel=1
    -4, 2, 7, 5, 0, -3, -6, -8, -8,
    -- filter=51 channel=2
    9, -7, -7, -8, 9, 2, -8, 1, -4,
    -- filter=51 channel=3
    0, -8, -5, 3, 5, -3, -3, 9, 4,
    -- filter=51 channel=4
    -3, 6, 7, 6, 3, 4, 8, -3, 7,
    -- filter=51 channel=5
    -7, -9, 3, 6, 8, 6, 2, 2, -9,
    -- filter=51 channel=6
    -6, 10, -2, 3, -6, -5, 5, -5, -4,
    -- filter=51 channel=7
    10, 5, -8, -8, -9, 5, 1, -2, 0,
    -- filter=51 channel=8
    -5, -6, 2, 7, -5, -1, 2, -1, 4,
    -- filter=51 channel=9
    -7, 6, 3, 8, 9, -5, 7, -4, -7,
    -- filter=51 channel=10
    -5, 9, 2, -8, 0, 5, -6, 5, -3,
    -- filter=51 channel=11
    -8, -6, 7, 6, -3, 0, 5, -8, -8,
    -- filter=51 channel=12
    -2, 1, -1, -1, 3, 8, 8, -4, 4,
    -- filter=51 channel=13
    3, 7, 1, -4, -2, 8, 2, 2, 4,
    -- filter=51 channel=14
    8, 4, 8, 2, -4, 5, 7, 5, 1,
    -- filter=51 channel=15
    -6, 1, -5, -3, 0, -6, -3, -2, 0,
    -- filter=51 channel=16
    -6, -7, 3, 7, -8, 10, -4, -1, 4,
    -- filter=51 channel=17
    -3, 4, -8, -6, 7, -5, -10, -8, -9,
    -- filter=51 channel=18
    0, -1, -9, 2, 4, 1, -8, -3, 5,
    -- filter=51 channel=19
    -5, 6, 5, 1, 2, -9, -6, -5, 5,
    -- filter=51 channel=20
    0, -1, 3, 0, 8, 10, 7, 7, 3,
    -- filter=51 channel=21
    10, 3, 1, 7, -2, 10, 0, 8, -7,
    -- filter=51 channel=22
    9, -3, -1, -10, 7, -2, -1, -10, 0,
    -- filter=51 channel=23
    1, 8, -5, 9, -10, 5, -7, 0, 0,
    -- filter=51 channel=24
    -9, 0, 7, 0, -7, 5, -1, 6, 10,
    -- filter=51 channel=25
    8, -10, -3, -10, 10, 4, -3, -8, -5,
    -- filter=51 channel=26
    3, 6, 1, 0, -3, 5, 0, 3, -5,
    -- filter=51 channel=27
    3, 5, -5, 5, 9, 2, 1, -8, 10,
    -- filter=51 channel=28
    9, -4, 3, 7, 9, 5, 2, -6, 11,
    -- filter=51 channel=29
    -8, -9, 2, -9, -7, 0, 4, 5, 3,
    -- filter=51 channel=30
    -5, -1, -3, -5, 0, 5, -3, 7, -10,
    -- filter=51 channel=31
    0, -8, -2, -1, 5, -2, -3, 5, 4,
    -- filter=51 channel=32
    -9, 5, -2, -4, -4, 0, -8, 5, -1,
    -- filter=51 channel=33
    -1, -8, -4, 8, 6, -1, 7, -7, 0,
    -- filter=51 channel=34
    7, -9, 5, -1, 9, 2, 0, 10, -7,
    -- filter=51 channel=35
    3, 1, 8, -1, -3, -6, 9, -9, 9,
    -- filter=51 channel=36
    5, -2, 0, -10, 1, -1, 0, 7, -7,
    -- filter=51 channel=37
    -8, 0, -5, 3, 10, 2, 5, -6, 3,
    -- filter=51 channel=38
    -2, 5, 2, 3, -1, 2, -10, 1, -4,
    -- filter=51 channel=39
    7, -3, 4, -3, -3, 1, 6, -7, -1,
    -- filter=51 channel=40
    0, 1, -1, -9, -2, -8, -5, 5, -4,
    -- filter=51 channel=41
    -2, -3, 2, -6, 0, 6, 4, 8, -1,
    -- filter=51 channel=42
    6, -2, 3, -9, 7, 1, 1, -5, -8,
    -- filter=51 channel=43
    10, 10, 2, 4, -7, -2, 0, 3, 0,
    -- filter=51 channel=44
    0, 2, -1, 3, -6, 2, -8, 2, 10,
    -- filter=51 channel=45
    -7, -5, -1, 6, 7, -6, -4, -7, -6,
    -- filter=51 channel=46
    7, -4, 0, -5, 7, 7, -3, 2, 8,
    -- filter=51 channel=47
    9, -8, -5, 0, 9, -4, -7, -3, -10,
    -- filter=51 channel=48
    0, 9, 9, 1, -5, 4, 3, 2, 4,
    -- filter=51 channel=49
    -9, 3, -9, 2, 8, -9, 7, 0, -8,
    -- filter=51 channel=50
    7, 9, -7, -1, 7, 2, -1, 2, -9,
    -- filter=51 channel=51
    10, 0, -5, -9, 8, 1, 2, -7, 3,
    -- filter=51 channel=52
    -8, -3, 6, -3, 8, -9, -6, 3, 5,
    -- filter=51 channel=53
    5, -3, 7, -7, 3, -8, 5, -5, 9,
    -- filter=51 channel=54
    3, 5, 2, -1, 11, 11, -5, 4, 5,
    -- filter=51 channel=55
    9, 6, 0, -2, 4, 10, -4, 3, -6,
    -- filter=51 channel=56
    4, -10, -8, -8, -2, 4, -9, 3, 3,
    -- filter=51 channel=57
    5, -6, -6, 1, -4, -3, 1, 9, -4,
    -- filter=51 channel=58
    -9, -10, -3, -6, 4, -9, 6, 2, -9,
    -- filter=51 channel=59
    5, -8, -3, -8, -9, -5, 8, 0, 9,
    -- filter=51 channel=60
    -8, 10, -7, -6, -6, 3, 0, -6, -8,
    -- filter=51 channel=61
    10, 0, 3, -7, 1, -6, -6, 0, 2,
    -- filter=51 channel=62
    1, -3, 4, 8, -8, -3, 2, -9, 0,
    -- filter=51 channel=63
    4, -5, 6, 10, 5, 3, -3, -4, 7,
    -- filter=52 channel=0
    -3, -2, -1, -9, -5, 16, 0, 2, 5,
    -- filter=52 channel=1
    -16, 0, 1, -21, -15, -3, -17, -17, -1,
    -- filter=52 channel=2
    -15, -10, 6, -22, -18, 6, -7, 3, 7,
    -- filter=52 channel=3
    -6, -6, 3, -7, 13, 0, 0, -5, -6,
    -- filter=52 channel=4
    2, -2, 2, -12, 9, 14, 8, 0, -4,
    -- filter=52 channel=5
    -4, 11, 14, 2, 15, 12, 7, 11, 10,
    -- filter=52 channel=6
    -9, -2, 0, 0, 7, -5, -13, 9, -4,
    -- filter=52 channel=7
    14, 8, 7, 1, 18, 18, 10, 14, 18,
    -- filter=52 channel=8
    -15, -3, -4, -5, 11, 3, -10, 8, 18,
    -- filter=52 channel=9
    3, 10, 4, 10, 9, 0, 9, 13, 1,
    -- filter=52 channel=10
    5, -7, 5, -3, 6, -7, 4, -8, -3,
    -- filter=52 channel=11
    3, -11, -7, -7, 2, -5, -11, 6, 2,
    -- filter=52 channel=12
    -1, 4, 5, 5, 8, 10, 10, 1, 6,
    -- filter=52 channel=13
    0, 7, 2, -11, 7, 6, -12, 3, 11,
    -- filter=52 channel=14
    15, 20, 5, 4, 14, 2, 1, 6, 4,
    -- filter=52 channel=15
    -13, -4, 14, -1, 4, 17, -13, 0, 4,
    -- filter=52 channel=16
    0, 2, 8, -6, -6, 5, -14, 3, 6,
    -- filter=52 channel=17
    -12, -7, -1, -6, -8, 2, -10, 12, 1,
    -- filter=52 channel=18
    9, 4, 6, 4, 6, 5, 6, 16, -1,
    -- filter=52 channel=19
    -8, 10, -10, 4, -7, 4, 2, -2, -4,
    -- filter=52 channel=20
    5, 14, 16, 20, 7, 7, 16, 22, 6,
    -- filter=52 channel=21
    8, -3, 5, 6, -4, -6, 9, -9, -8,
    -- filter=52 channel=22
    3, 0, -7, -1, -1, 5, 1, 3, -2,
    -- filter=52 channel=23
    1, 6, 1, 3, -9, 5, 2, -4, 11,
    -- filter=52 channel=24
    -4, 9, 5, -16, -9, 14, -1, 11, 13,
    -- filter=52 channel=25
    -8, -4, 0, -13, 0, 6, -13, -16, 0,
    -- filter=52 channel=26
    22, 6, 5, 5, 8, 11, 2, 23, 13,
    -- filter=52 channel=27
    -14, -14, 0, -25, 3, -3, -16, -11, 9,
    -- filter=52 channel=28
    -1, 3, -12, -18, 10, -5, -8, 9, -7,
    -- filter=52 channel=29
    -4, 8, 10, -15, 15, 11, -9, 16, -2,
    -- filter=52 channel=30
    33, 25, 23, 35, 37, 35, 26, 37, 24,
    -- filter=52 channel=31
    -7, 6, -8, -4, 4, 2, -2, -10, 7,
    -- filter=52 channel=32
    -1, 8, -6, -1, 1, 4, 6, -9, 7,
    -- filter=52 channel=33
    0, -4, -5, 0, 4, -6, -9, 5, -8,
    -- filter=52 channel=34
    0, 13, 10, 17, 0, 6, -1, 9, 1,
    -- filter=52 channel=35
    -12, 1, 6, -14, 0, -3, 0, 0, 6,
    -- filter=52 channel=36
    10, -10, -3, 5, 0, -1, -9, -7, 5,
    -- filter=52 channel=37
    7, -8, -2, -2, 11, 10, 2, -3, 5,
    -- filter=52 channel=38
    -5, -2, 0, -11, 0, 5, -22, 0, 0,
    -- filter=52 channel=39
    5, -4, -9, 2, 5, 0, -1, -10, 6,
    -- filter=52 channel=40
    0, 0, 2, 6, 5, 7, 4, -6, 4,
    -- filter=52 channel=41
    -4, -1, -2, -20, -4, 12, 1, 3, 12,
    -- filter=52 channel=42
    -3, -7, 1, -4, 3, -3, -3, 0, 1,
    -- filter=52 channel=43
    17, 16, 12, 10, 8, 5, 11, 0, 8,
    -- filter=52 channel=44
    8, 12, 13, -1, -4, 8, -5, 3, 18,
    -- filter=52 channel=45
    -5, -7, 0, 1, 1, 7, 9, 8, 2,
    -- filter=52 channel=46
    11, 13, 23, 19, 16, 20, 24, 6, 8,
    -- filter=52 channel=47
    -1, 5, 10, 0, 9, -6, 9, -8, 2,
    -- filter=52 channel=48
    11, 9, 4, 2, -2, 13, 8, -1, -7,
    -- filter=52 channel=49
    -16, -5, 6, 2, -9, 5, -4, 6, 6,
    -- filter=52 channel=50
    13, 28, 16, 15, 25, 11, 12, 7, 12,
    -- filter=52 channel=51
    1, 11, -4, -3, 1, -5, 0, 8, 5,
    -- filter=52 channel=52
    0, -3, 3, 0, 0, -2, 8, 5, -1,
    -- filter=52 channel=53
    17, 17, 17, 7, 10, 24, 7, 23, 22,
    -- filter=52 channel=54
    -1, 0, 6, -7, 10, 2, -5, 1, 10,
    -- filter=52 channel=55
    -9, -5, -6, -9, 8, -8, 2, 2, 10,
    -- filter=52 channel=56
    13, -4, 11, 1, 13, 0, 11, 7, 6,
    -- filter=52 channel=57
    6, 2, 8, -2, -2, -6, -1, -6, 1,
    -- filter=52 channel=58
    7, -7, 3, 0, 0, 4, 3, 6, -11,
    -- filter=52 channel=59
    -5, -1, 5, -12, 9, 3, -7, 1, 13,
    -- filter=52 channel=60
    4, 11, 13, -17, 11, 16, -7, 9, 12,
    -- filter=52 channel=61
    7, 0, -7, -5, -3, 16, -13, 5, 6,
    -- filter=52 channel=62
    -1, 11, -3, -3, 0, 13, -10, -5, -5,
    -- filter=52 channel=63
    1, 0, -1, 8, 3, 7, 6, -3, 9,
    -- filter=53 channel=0
    -7, -3, -7, -8, 0, 8, -2, 4, -8,
    -- filter=53 channel=1
    -3, -4, -14, 0, 4, -14, -4, 0, -4,
    -- filter=53 channel=2
    -4, -1, -10, -12, -5, 3, -6, -11, -10,
    -- filter=53 channel=3
    0, 9, 8, -6, 6, -4, -7, -4, 2,
    -- filter=53 channel=4
    0, 3, 4, -8, 10, 0, 7, 6, 2,
    -- filter=53 channel=5
    -8, 2, 7, 12, 8, 12, 0, -6, -5,
    -- filter=53 channel=6
    -9, -1, 6, 6, 6, -2, 4, -6, -5,
    -- filter=53 channel=7
    -10, -2, 3, -1, 10, -2, 9, 7, 2,
    -- filter=53 channel=8
    -7, 3, 0, -3, 8, 8, -6, 7, 3,
    -- filter=53 channel=9
    16, 17, 20, 21, 31, 15, 9, 15, 11,
    -- filter=53 channel=10
    4, 2, 8, -3, -5, -11, 10, -10, -1,
    -- filter=53 channel=11
    1, 1, 3, 3, -9, 4, 0, 0, -6,
    -- filter=53 channel=12
    -4, -6, 2, -7, 3, 5, 3, -3, 9,
    -- filter=53 channel=13
    3, 0, 5, 7, 0, 8, 10, 5, 13,
    -- filter=53 channel=14
    10, -7, 3, -4, 7, -1, -4, 0, 9,
    -- filter=53 channel=15
    9, 7, -4, -6, 6, 15, -9, 9, 0,
    -- filter=53 channel=16
    -3, 1, 8, -5, -1, -1, -1, -2, 6,
    -- filter=53 channel=17
    3, 0, -2, 3, 12, 0, -5, 1, 7,
    -- filter=53 channel=18
    7, 17, -4, 14, 8, 4, 7, 5, 14,
    -- filter=53 channel=19
    -3, -5, 10, -6, 10, 4, -9, -1, -6,
    -- filter=53 channel=20
    5, 1, -2, 10, 5, 15, 7, -2, -4,
    -- filter=53 channel=21
    -1, 0, -6, 10, 6, 0, 2, 1, 11,
    -- filter=53 channel=22
    -3, 2, -8, 0, -10, -6, 10, -6, -9,
    -- filter=53 channel=23
    -5, -8, -11, 5, -16, -4, -4, -12, -11,
    -- filter=53 channel=24
    7, 2, 9, -10, -1, 3, -3, 11, 5,
    -- filter=53 channel=25
    -11, 0, 2, 0, -4, -8, -8, -18, -13,
    -- filter=53 channel=26
    8, -9, 4, -6, -3, 8, -7, -7, 2,
    -- filter=53 channel=27
    -10, -13, -5, 5, -10, -15, -10, 2, -14,
    -- filter=53 channel=28
    -8, 5, -1, 0, 1, 11, -3, 11, 9,
    -- filter=53 channel=29
    6, 3, -5, 7, -2, 7, -2, 8, 1,
    -- filter=53 channel=30
    -4, -4, -7, 6, -6, -12, -10, 1, -5,
    -- filter=53 channel=31
    5, -1, -4, 11, 2, 0, -6, 0, 5,
    -- filter=53 channel=32
    -7, -2, 8, 2, -11, -3, 8, 6, -4,
    -- filter=53 channel=33
    2, -7, 1, -1, 0, -3, -6, 1, -3,
    -- filter=53 channel=34
    -2, 0, -7, -3, 1, 9, -9, 3, -1,
    -- filter=53 channel=35
    -1, -14, -7, 0, -11, -16, -15, -3, -4,
    -- filter=53 channel=36
    -6, 7, -7, 8, 5, 2, 2, 7, 9,
    -- filter=53 channel=37
    -6, 11, 5, 12, 10, 3, 0, 4, 11,
    -- filter=53 channel=38
    -4, 1, -1, -2, -8, 0, 0, -10, -7,
    -- filter=53 channel=39
    4, -4, 9, 9, -6, -1, 6, 5, 1,
    -- filter=53 channel=40
    0, 0, 0, -8, -7, 0, 2, -11, -4,
    -- filter=53 channel=41
    2, -5, 8, 10, -2, -4, -1, 2, 3,
    -- filter=53 channel=42
    -9, 3, 0, -4, -7, -4, 2, -5, -1,
    -- filter=53 channel=43
    -12, -12, 1, -3, 0, -7, -8, -1, -9,
    -- filter=53 channel=44
    1, -1, -1, -3, -14, 5, 6, -10, 2,
    -- filter=53 channel=45
    -8, -2, -4, 1, -2, -4, -1, 9, -1,
    -- filter=53 channel=46
    -2, 4, -7, 6, 9, -3, 2, 8, 10,
    -- filter=53 channel=47
    6, -7, 0, 7, -1, 2, -5, -2, -7,
    -- filter=53 channel=48
    -8, 5, 5, 7, -2, -1, -7, 0, -3,
    -- filter=53 channel=49
    7, -8, 1, -7, -9, -7, 5, 7, -9,
    -- filter=53 channel=50
    -11, -1, 10, -6, 0, 5, 10, 4, -3,
    -- filter=53 channel=51
    -7, 0, 10, -5, -5, 1, 4, 0, 6,
    -- filter=53 channel=52
    -3, 5, -2, -3, -8, 4, 6, 9, 4,
    -- filter=53 channel=53
    -8, -2, 6, 4, 5, -10, -6, -3, 7,
    -- filter=53 channel=54
    0, 21, 21, 10, 10, 14, 15, 17, 17,
    -- filter=53 channel=55
    6, 7, -7, 4, 1, -2, 7, 5, 0,
    -- filter=53 channel=56
    -6, 5, 6, -1, 0, -3, 2, 0, 3,
    -- filter=53 channel=57
    0, 10, -5, 3, 0, -9, 2, -9, 2,
    -- filter=53 channel=58
    6, 6, 5, 8, -3, 7, -5, -6, 4,
    -- filter=53 channel=59
    7, -4, -5, 2, -5, 12, 3, -2, 0,
    -- filter=53 channel=60
    3, -8, 1, 7, 0, 16, 1, 3, 8,
    -- filter=53 channel=61
    0, -9, 4, -10, -4, 7, -7, 10, 4,
    -- filter=53 channel=62
    7, -6, 12, 5, -2, 9, -6, 7, 1,
    -- filter=53 channel=63
    -8, -6, -5, -9, 9, -8, 6, -1, 5,
    -- filter=54 channel=0
    0, 6, 7, 2, -6, -1, 3, 1, -3,
    -- filter=54 channel=1
    -1, 4, -4, 5, 10, -10, 3, 2, 4,
    -- filter=54 channel=2
    2, -5, 9, 0, -10, -2, 2, -8, 0,
    -- filter=54 channel=3
    5, 1, 9, 10, -8, 10, 9, -8, -6,
    -- filter=54 channel=4
    -1, -6, 7, -4, -6, 7, 1, -4, 4,
    -- filter=54 channel=5
    -5, 7, 8, 7, -3, 1, -10, 7, 8,
    -- filter=54 channel=6
    -6, 4, -8, -2, -7, -5, -6, -10, 5,
    -- filter=54 channel=7
    -6, 0, -8, 6, 8, 0, 6, 6, 4,
    -- filter=54 channel=8
    4, -8, 4, -8, -1, -5, 4, 3, -10,
    -- filter=54 channel=9
    -9, 2, 2, -2, 1, 6, 7, -3, 1,
    -- filter=54 channel=10
    0, 10, -9, 0, -3, -10, 2, -8, -6,
    -- filter=54 channel=11
    -10, 5, 3, -4, 4, 5, -8, 7, -7,
    -- filter=54 channel=12
    3, -5, 1, -1, 9, -6, -3, 4, 0,
    -- filter=54 channel=13
    3, 6, -9, -6, -4, -9, 0, 6, 1,
    -- filter=54 channel=14
    -4, 3, 2, 3, 0, 8, 0, -9, 2,
    -- filter=54 channel=15
    -8, 0, 0, 10, 8, -10, 7, 2, -9,
    -- filter=54 channel=16
    0, 7, -1, -1, 5, -6, 3, 2, 8,
    -- filter=54 channel=17
    3, -4, 0, 10, 2, 10, -10, 0, 10,
    -- filter=54 channel=18
    -8, 0, 4, 8, -5, 4, -1, 4, 6,
    -- filter=54 channel=19
    2, -4, -7, -5, -9, -2, 0, -5, -1,
    -- filter=54 channel=20
    -4, -5, -4, 6, 0, -6, 6, -10, 4,
    -- filter=54 channel=21
    -9, -5, 0, -6, -2, -1, -6, -1, 9,
    -- filter=54 channel=22
    -1, -4, -6, 10, 9, 10, 6, 3, 3,
    -- filter=54 channel=23
    3, -10, -2, -3, 0, -6, 8, -8, 0,
    -- filter=54 channel=24
    -5, -5, -1, 7, 9, -9, -7, 9, 2,
    -- filter=54 channel=25
    0, -7, 7, -4, 10, 1, -1, 0, 4,
    -- filter=54 channel=26
    -5, 7, 1, 4, -5, 2, -10, -3, 7,
    -- filter=54 channel=27
    5, -6, 5, -4, -6, 0, -2, -8, -1,
    -- filter=54 channel=28
    3, -2, 1, 1, 4, 9, -2, 3, -1,
    -- filter=54 channel=29
    0, 0, 4, -5, -3, 6, 1, 8, 8,
    -- filter=54 channel=30
    -2, 3, -1, -5, 8, -6, 0, 8, -1,
    -- filter=54 channel=31
    1, 0, 1, -9, 2, -1, 0, -8, 4,
    -- filter=54 channel=32
    -3, -6, -5, -7, 1, 10, 7, 3, 5,
    -- filter=54 channel=33
    7, 7, 10, 9, -10, -1, 2, 0, -8,
    -- filter=54 channel=34
    -7, -4, 6, 0, -1, -9, -5, 4, 0,
    -- filter=54 channel=35
    -2, 5, -8, 0, 0, 6, -10, 8, -2,
    -- filter=54 channel=36
    -4, 5, -4, -5, -8, 3, 10, -9, -3,
    -- filter=54 channel=37
    -4, 7, -3, 1, 9, -3, 5, -8, 2,
    -- filter=54 channel=38
    6, 1, -6, -9, 4, 0, -8, -9, 9,
    -- filter=54 channel=39
    -3, -6, 9, 0, 4, 2, 8, -8, 1,
    -- filter=54 channel=40
    4, -4, -1, -3, -2, 8, -6, 0, -2,
    -- filter=54 channel=41
    3, -9, 4, -4, -4, -8, -6, -4, -1,
    -- filter=54 channel=42
    3, -10, 10, 7, 4, -8, 9, 0, -6,
    -- filter=54 channel=43
    0, 2, 5, -6, -10, -3, -4, -4, 2,
    -- filter=54 channel=44
    -3, 0, -9, 10, -1, -7, -4, 4, -1,
    -- filter=54 channel=45
    8, -7, 3, 6, -4, -10, 1, 5, -1,
    -- filter=54 channel=46
    3, 7, -7, 9, 4, -9, -8, -10, -5,
    -- filter=54 channel=47
    8, 2, 0, -4, 9, 7, 5, -10, 7,
    -- filter=54 channel=48
    -1, -8, 1, -5, 4, 6, 2, 0, -8,
    -- filter=54 channel=49
    0, 4, 0, -5, 6, -1, -3, -1, -1,
    -- filter=54 channel=50
    -10, -2, 9, -9, 6, 0, -4, 7, 4,
    -- filter=54 channel=51
    -3, 6, 5, -4, -5, 8, 6, -5, -7,
    -- filter=54 channel=52
    5, 2, 10, 0, -8, -8, 7, -4, 2,
    -- filter=54 channel=53
    -4, -2, -9, -2, -4, 8, -4, 2, 0,
    -- filter=54 channel=54
    7, -1, -10, -5, 4, -8, 4, -6, -1,
    -- filter=54 channel=55
    8, 1, 5, 2, -5, 0, -7, 10, 4,
    -- filter=54 channel=56
    8, 1, 3, -1, -1, 2, 10, 6, 0,
    -- filter=54 channel=57
    3, 0, -8, 0, -1, 7, -7, 10, 8,
    -- filter=54 channel=58
    8, -3, 2, 1, -10, 9, 7, -5, 1,
    -- filter=54 channel=59
    -5, 6, 9, -5, 1, 9, 8, 0, 6,
    -- filter=54 channel=60
    -2, -3, 2, -9, 1, -8, 7, -7, -1,
    -- filter=54 channel=61
    -1, 6, -9, 3, -2, 0, -9, -4, -10,
    -- filter=54 channel=62
    0, 0, 6, 4, -4, 0, -2, -7, -8,
    -- filter=54 channel=63
    -7, 0, -8, 5, 8, 4, -5, 7, 7,
    -- filter=55 channel=0
    -2, 3, -9, -2, -5, 8, -11, -2, -7,
    -- filter=55 channel=1
    -4, -16, -3, -7, -10, -10, -16, -1, -7,
    -- filter=55 channel=2
    -13, 2, 5, -8, -2, -9, -20, -15, -16,
    -- filter=55 channel=3
    13, 11, 1, -1, 12, 3, -1, 0, 9,
    -- filter=55 channel=4
    11, 11, -6, 15, 12, 13, 0, 5, 11,
    -- filter=55 channel=5
    18, 4, 7, 17, 3, 2, 8, 10, -4,
    -- filter=55 channel=6
    -8, 3, 2, 4, -3, -4, -6, -14, 3,
    -- filter=55 channel=7
    1, -5, 6, 8, 4, 6, 9, 8, 12,
    -- filter=55 channel=8
    7, 14, 3, -1, 1, 0, 2, -2, 2,
    -- filter=55 channel=9
    20, 30, 31, 25, 37, 37, 29, 27, 26,
    -- filter=55 channel=10
    2, -4, 4, -18, -4, -15, -10, -16, -6,
    -- filter=55 channel=11
    -14, 6, 4, -11, 5, 1, 7, 3, -9,
    -- filter=55 channel=12
    7, 7, 9, -8, 0, 9, -3, 8, 5,
    -- filter=55 channel=13
    14, 11, 8, 6, 5, 6, 8, 7, -6,
    -- filter=55 channel=14
    2, 4, -8, -1, 9, 12, -1, 0, -5,
    -- filter=55 channel=15
    11, 19, 7, 8, 4, 1, 3, 7, -8,
    -- filter=55 channel=16
    6, 14, -7, 1, 19, 2, -6, 8, -12,
    -- filter=55 channel=17
    12, 4, 11, 8, 2, 7, 11, 7, -3,
    -- filter=55 channel=18
    15, 11, 4, 9, 16, -1, 10, 12, 3,
    -- filter=55 channel=19
    3, 9, 8, 7, 22, 5, -1, -1, 10,
    -- filter=55 channel=20
    6, 11, 3, 8, 15, 5, 7, 3, 13,
    -- filter=55 channel=21
    8, 7, -7, -1, -1, -7, 6, 8, -9,
    -- filter=55 channel=22
    7, 7, -8, 9, 4, -4, 8, -7, -2,
    -- filter=55 channel=23
    -17, -7, -5, -17, -9, -6, -14, -17, 1,
    -- filter=55 channel=24
    1, 13, 0, 0, 11, 6, 10, 1, -1,
    -- filter=55 channel=25
    -19, -14, 0, -15, -21, -8, -23, -13, -7,
    -- filter=55 channel=26
    -2, -2, -5, 2, 1, -5, 1, 13, -4,
    -- filter=55 channel=27
    -13, -5, -8, -2, -5, -6, -12, -5, -5,
    -- filter=55 channel=28
    -4, 9, 1, 18, 16, -3, 10, 17, 3,
    -- filter=55 channel=29
    18, 14, 9, 11, 28, 3, 0, 20, -2,
    -- filter=55 channel=30
    -8, 10, 0, -6, 11, 10, 11, 0, 13,
    -- filter=55 channel=31
    6, 1, 8, 2, -6, 1, 2, 3, -5,
    -- filter=55 channel=32
    -19, -2, 3, -3, -5, 7, -4, 0, 6,
    -- filter=55 channel=33
    -8, -3, 0, -7, -4, 3, 0, -1, -9,
    -- filter=55 channel=34
    -8, -3, -7, 9, -2, 7, 13, 1, -2,
    -- filter=55 channel=35
    -18, -25, -6, -39, -26, -15, -33, -31, -16,
    -- filter=55 channel=36
    0, -4, -8, -2, -13, 0, -4, 5, -1,
    -- filter=55 channel=37
    0, 21, 11, 19, 9, -1, 2, 13, 7,
    -- filter=55 channel=38
    -4, -12, 2, -2, 0, 4, 2, -2, 0,
    -- filter=55 channel=39
    -7, 0, 0, 10, -2, 10, 0, 7, 0,
    -- filter=55 channel=40
    -3, 0, 3, 5, -14, 4, 5, -4, 1,
    -- filter=55 channel=41
    13, 9, -6, 0, 8, -7, -9, 0, -10,
    -- filter=55 channel=42
    7, 9, 8, 0, -1, -8, 9, 0, 2,
    -- filter=55 channel=43
    -24, -16, -24, -12, -12, -22, -5, -13, -22,
    -- filter=55 channel=44
    -13, 3, 0, -11, -9, 7, -12, 3, -6,
    -- filter=55 channel=45
    -5, -1, 7, -5, -9, -2, 9, 5, 5,
    -- filter=55 channel=46
    2, 15, -3, 0, 17, -3, 11, 0, 8,
    -- filter=55 channel=47
    -9, -3, 0, -3, 5, 5, -9, -5, 7,
    -- filter=55 channel=48
    -4, 9, -3, 15, 5, 12, 9, 7, 10,
    -- filter=55 channel=49
    -12, -11, -5, 2, -9, 0, -5, -3, -10,
    -- filter=55 channel=50
    -3, 2, -2, 14, -3, 0, 6, 1, 10,
    -- filter=55 channel=51
    -4, -3, 9, -10, -17, 8, 4, 5, 3,
    -- filter=55 channel=52
    -7, 5, 1, 1, 9, 8, -6, 9, 3,
    -- filter=55 channel=53
    -9, -8, 2, -3, -8, -3, 3, -3, 12,
    -- filter=55 channel=54
    12, 18, 20, 32, 43, 32, 23, 24, 5,
    -- filter=55 channel=55
    5, 7, 0, -9, 5, -6, 7, -5, -10,
    -- filter=55 channel=56
    0, -2, -6, -1, 6, 0, 4, 5, -2,
    -- filter=55 channel=57
    -5, -1, -8, 1, 0, 3, 11, 6, 4,
    -- filter=55 channel=58
    6, -1, -3, -7, 4, 1, 12, -1, 5,
    -- filter=55 channel=59
    -7, 5, 11, -4, -5, -1, -8, 1, 0,
    -- filter=55 channel=60
    8, 3, 1, 13, 22, 3, 2, -1, 7,
    -- filter=55 channel=61
    2, 0, 12, 6, 3, 7, 0, 7, -3,
    -- filter=55 channel=62
    -2, 13, 5, 3, 8, -2, 10, 3, 2,
    -- filter=55 channel=63
    -3, -10, 10, -6, 10, -5, 0, 10, 4,
    -- filter=56 channel=0
    -10, -2, -5, 2, -9, 12, -15, -5, 4,
    -- filter=56 channel=1
    2, 4, -10, 0, -13, 10, 5, -7, 7,
    -- filter=56 channel=2
    8, -18, 13, -8, -18, 10, -1, -14, 12,
    -- filter=56 channel=3
    0, -1, 12, 3, 3, 1, -9, 4, 10,
    -- filter=56 channel=4
    1, 0, -6, -9, -3, 0, -8, 9, 2,
    -- filter=56 channel=5
    6, 3, -6, 11, 4, 2, 11, 4, 9,
    -- filter=56 channel=6
    1, -11, 10, -13, 5, 12, 0, 4, 14,
    -- filter=56 channel=7
    0, 15, 7, 11, 11, -5, 15, 11, 0,
    -- filter=56 channel=8
    7, -19, 11, 6, -4, 9, 0, -4, 11,
    -- filter=56 channel=9
    2, -2, 3, -4, -5, 6, 3, 3, -6,
    -- filter=56 channel=10
    0, -1, -4, 7, 10, -7, -7, 5, -5,
    -- filter=56 channel=11
    13, -8, 4, 16, -1, 0, -3, 1, 16,
    -- filter=56 channel=12
    -6, 2, 3, 5, -10, -4, 0, -5, 5,
    -- filter=56 channel=13
    6, 3, -2, -4, -3, 7, -14, -2, 1,
    -- filter=56 channel=14
    1, 1, 13, 1, 4, 10, 0, 12, -3,
    -- filter=56 channel=15
    -6, -18, 3, -7, -5, 26, -1, 1, 3,
    -- filter=56 channel=16
    8, -21, -2, -1, -8, 7, -3, -15, 17,
    -- filter=56 channel=17
    8, -15, -4, 6, -14, 9, 2, -11, 6,
    -- filter=56 channel=18
    -5, -1, -9, 2, 4, -2, -1, 4, -5,
    -- filter=56 channel=19
    3, -7, -8, 15, -4, 10, -1, 0, 10,
    -- filter=56 channel=20
    -1, 3, 17, -2, -2, 2, 0, -1, 0,
    -- filter=56 channel=21
    0, -9, -9, 3, -9, 3, 0, -8, -9,
    -- filter=56 channel=22
    0, 9, -10, -5, 8, 1, 4, 0, -5,
    -- filter=56 channel=23
    1, -3, 6, 9, 2, 7, -9, -7, 1,
    -- filter=56 channel=24
    5, 6, -5, 17, -6, 4, 1, -1, 3,
    -- filter=56 channel=25
    -6, -22, 4, -16, -21, 6, -11, -14, 16,
    -- filter=56 channel=26
    -1, 11, 15, 2, 0, 9, 10, 11, 19,
    -- filter=56 channel=27
    8, -19, 11, -2, -20, 11, -9, -11, 8,
    -- filter=56 channel=28
    18, -11, -4, 14, 3, 1, -3, 0, 5,
    -- filter=56 channel=29
    -4, -4, -3, -5, -4, 19, -10, -12, 6,
    -- filter=56 channel=30
    18, 18, 15, 19, 21, 28, 14, 0, 15,
    -- filter=56 channel=31
    5, 2, 6, 3, -1, -8, -2, -9, -9,
    -- filter=56 channel=32
    8, -6, 9, 1, 2, -5, 0, -11, 6,
    -- filter=56 channel=33
    -7, -9, 9, 1, -7, 8, 5, -5, 0,
    -- filter=56 channel=34
    12, 8, -4, -5, 12, 16, 12, 1, 7,
    -- filter=56 channel=35
    -12, -14, 13, -4, -12, 11, -14, -5, 19,
    -- filter=56 channel=36
    0, 9, -6, 7, -2, 4, 3, -1, -6,
    -- filter=56 channel=37
    7, -8, 2, 4, -11, 1, -5, -6, 9,
    -- filter=56 channel=38
    9, -20, -6, -12, -23, 17, -3, -11, 18,
    -- filter=56 channel=39
    -2, 8, 9, 0, 2, -2, -3, -6, 10,
    -- filter=56 channel=40
    -4, 8, -2, 7, -12, 0, 2, 9, 0,
    -- filter=56 channel=41
    10, -10, 7, -6, -8, 28, -2, -9, 21,
    -- filter=56 channel=42
    -6, -3, -5, 3, -7, -2, -6, -3, 9,
    -- filter=56 channel=43
    5, 6, -9, 3, -13, 1, -5, -6, 9,
    -- filter=56 channel=44
    6, 0, -2, -4, 1, -5, 0, 0, -4,
    -- filter=56 channel=45
    2, 9, -7, -1, 8, -5, -5, 7, 8,
    -- filter=56 channel=46
    -2, 2, 18, 3, 9, 8, -1, 0, 14,
    -- filter=56 channel=47
    -6, -6, 2, 10, -9, -8, 7, -7, 4,
    -- filter=56 channel=48
    -1, -12, 6, -12, 10, -1, -9, 1, 2,
    -- filter=56 channel=49
    2, 1, 10, -9, -10, 17, -4, 0, 5,
    -- filter=56 channel=50
    17, 19, 13, 21, 14, 10, 23, -3, 0,
    -- filter=56 channel=51
    1, -3, 0, 5, 3, -9, 5, 0, 0,
    -- filter=56 channel=52
    5, -2, -6, -9, 6, 9, -10, -9, 4,
    -- filter=56 channel=53
    9, 20, 15, 18, 1, 14, 22, -2, 6,
    -- filter=56 channel=54
    0, 0, 4, 10, 1, -5, 6, -3, -7,
    -- filter=56 channel=55
    -5, 2, 7, -7, 4, 6, 4, 2, -9,
    -- filter=56 channel=56
    -5, -1, -1, 6, 9, 9, -3, 0, 1,
    -- filter=56 channel=57
    -6, 4, -2, -6, 0, 3, 1, 7, 1,
    -- filter=56 channel=58
    -7, 9, -4, -13, 4, 1, -5, 1, -11,
    -- filter=56 channel=59
    -5, -15, 10, -5, -3, 16, -7, 5, 6,
    -- filter=56 channel=60
    -6, -8, 7, 6, -18, 25, -16, -13, 29,
    -- filter=56 channel=61
    16, -12, -10, 16, -20, 19, -1, -3, 16,
    -- filter=56 channel=62
    -4, 1, 0, 0, -18, 10, 4, -4, 9,
    -- filter=56 channel=63
    -8, 10, -1, 0, 0, 5, -4, 10, -7,
    -- filter=57 channel=0
    -2, -8, 13, -2, -13, -5, -1, 0, 1,
    -- filter=57 channel=1
    1, 2, 4, -3, -3, -2, -7, -2, -8,
    -- filter=57 channel=2
    -4, -5, -5, 5, -3, 0, 6, 3, -10,
    -- filter=57 channel=3
    0, 6, -3, 6, 1, 2, 0, 0, -12,
    -- filter=57 channel=4
    -2, -4, -11, 2, -9, 7, 7, 11, 8,
    -- filter=57 channel=5
    10, 8, -4, -1, 0, 3, 7, 2, 0,
    -- filter=57 channel=6
    -4, 0, 6, 1, -8, -1, 13, 1, 4,
    -- filter=57 channel=7
    0, -1, -8, -7, -4, 10, -1, 8, 10,
    -- filter=57 channel=8
    -4, -16, -12, 6, 6, -11, 19, 6, 2,
    -- filter=57 channel=9
    7, 1, -5, -8, -10, -5, 5, 0, 8,
    -- filter=57 channel=10
    -9, -6, -7, 0, 4, -4, 11, -8, -4,
    -- filter=57 channel=11
    2, -3, -9, 9, -10, -3, 6, -1, -3,
    -- filter=57 channel=12
    5, 2, 0, 5, -7, 1, -3, -8, -1,
    -- filter=57 channel=13
    -12, 3, 1, 5, -15, -6, 9, -4, -5,
    -- filter=57 channel=14
    9, 6, -2, 8, 12, -5, 3, -5, 0,
    -- filter=57 channel=15
    5, -13, 8, 0, -16, 1, 20, 0, -5,
    -- filter=57 channel=16
    -1, -20, -5, 0, -7, 1, 13, 9, -9,
    -- filter=57 channel=17
    0, -6, -11, 3, 8, -14, -4, 12, 2,
    -- filter=57 channel=18
    2, -4, 2, 11, -4, 7, 8, -9, -6,
    -- filter=57 channel=19
    11, -8, 0, 1, 3, 0, -5, 2, -1,
    -- filter=57 channel=20
    2, 12, 13, -5, 7, 6, 12, 5, 12,
    -- filter=57 channel=21
    -3, -5, -6, -1, 3, 2, 9, 0, 9,
    -- filter=57 channel=22
    10, -7, 0, 4, -4, 0, -2, 10, -5,
    -- filter=57 channel=23
    -2, 0, -12, 8, 11, -9, -3, 9, -7,
    -- filter=57 channel=24
    6, -8, -14, 7, 2, -6, -1, 7, -3,
    -- filter=57 channel=25
    6, -7, -8, -5, -5, -9, 2, 3, -1,
    -- filter=57 channel=26
    -6, 10, 13, 3, 7, 10, -2, -3, 10,
    -- filter=57 channel=27
    9, -5, 4, 16, -2, -6, 16, 10, 4,
    -- filter=57 channel=28
    -6, -7, -13, 8, 0, -2, -1, 11, 0,
    -- filter=57 channel=29
    6, -23, 7, 15, -16, -15, 11, 9, 4,
    -- filter=57 channel=30
    -1, 15, 0, -4, 17, -1, -10, 20, -2,
    -- filter=57 channel=31
    1, 10, 7, 7, -4, -7, 6, -3, 6,
    -- filter=57 channel=32
    4, 11, -11, 5, 0, -3, -4, 4, 6,
    -- filter=57 channel=33
    -4, 6, 0, -3, 10, 3, -5, -6, 3,
    -- filter=57 channel=34
    1, 6, 2, -7, -2, 12, 8, -9, -2,
    -- filter=57 channel=35
    9, 0, 8, 4, 0, -8, 0, 0, -4,
    -- filter=57 channel=36
    0, 4, -5, 4, -2, -5, 0, 3, 7,
    -- filter=57 channel=37
    10, -5, 9, 3, -10, 3, 6, -4, -5,
    -- filter=57 channel=38
    -5, 0, 9, 10, -14, 0, 13, 8, 4,
    -- filter=57 channel=39
    9, 0, -6, -8, -1, -6, 0, 9, -6,
    -- filter=57 channel=40
    2, -4, 7, 0, -6, 5, 5, -4, 11,
    -- filter=57 channel=41
    -3, -12, 1, 16, 4, -4, 2, 12, -6,
    -- filter=57 channel=42
    -8, 1, 5, 1, 3, 10, 3, 9, -6,
    -- filter=57 channel=43
    4, 14, 0, -4, -2, 16, -2, 10, 11,
    -- filter=57 channel=44
    -5, 7, 0, -9, 2, -8, 5, 3, 2,
    -- filter=57 channel=45
    -3, -1, -3, -10, 7, -5, 10, -1, 2,
    -- filter=57 channel=46
    4, -4, -2, 2, 5, -1, -5, 2, 12,
    -- filter=57 channel=47
    9, 3, 6, 1, 6, -9, 1, -1, -8,
    -- filter=57 channel=48
    -8, -13, 5, -5, 3, 7, 9, -6, -1,
    -- filter=57 channel=49
    4, 0, -7, 16, 6, 1, -3, 4, 5,
    -- filter=57 channel=50
    -2, 1, 9, -2, -1, -6, 1, 1, 0,
    -- filter=57 channel=51
    1, -2, 5, -6, -7, -10, 8, 0, -6,
    -- filter=57 channel=52
    2, 7, -9, 7, -9, 7, -6, -3, -7,
    -- filter=57 channel=53
    0, 10, 7, 13, 15, -12, 0, 2, 8,
    -- filter=57 channel=54
    -4, 3, 4, 0, 9, -7, 12, 3, -1,
    -- filter=57 channel=55
    0, 2, -5, -1, -9, 6, -2, -1, 4,
    -- filter=57 channel=56
    -7, 4, 11, -6, 1, 1, -2, 2, 8,
    -- filter=57 channel=57
    -7, -2, -3, 8, -5, -5, 4, 9, 3,
    -- filter=57 channel=58
    -3, -4, -2, 1, -2, 3, 5, -10, 3,
    -- filter=57 channel=59
    4, -16, -1, -2, -5, 4, 12, 3, -12,
    -- filter=57 channel=60
    -5, -18, 4, 20, -4, -8, 28, 7, -13,
    -- filter=57 channel=61
    -5, 4, 4, 3, -10, -5, 12, 0, 6,
    -- filter=57 channel=62
    0, 2, -4, -6, 6, -10, 0, -1, -4,
    -- filter=57 channel=63
    0, 0, -3, -1, -6, 5, -6, 1, 4,
    -- filter=58 channel=0
    -1, 12, -1, 16, -2, 1, -3, 8, 0,
    -- filter=58 channel=1
    9, 4, 8, 10, 5, 2, 4, 7, 5,
    -- filter=58 channel=2
    4, 8, 14, -2, 7, -1, 13, 11, -2,
    -- filter=58 channel=3
    10, 0, -8, -9, -5, 7, 0, -4, 6,
    -- filter=58 channel=4
    5, -2, 0, -3, -1, -4, 0, 0, -10,
    -- filter=58 channel=5
    -3, -10, 8, -14, 5, 0, -7, 0, -2,
    -- filter=58 channel=6
    0, 12, 5, 4, 13, -3, 1, 14, -3,
    -- filter=58 channel=7
    -1, -8, -7, -3, -6, -6, -5, -2, -8,
    -- filter=58 channel=8
    -12, -13, 1, -12, -1, -1, -5, -11, 4,
    -- filter=58 channel=9
    -7, -12, 3, -11, -5, 15, 0, -9, 14,
    -- filter=58 channel=10
    5, 8, 10, 24, 11, 18, 13, 25, 16,
    -- filter=58 channel=11
    -7, 0, -6, 7, 0, 10, -9, -5, -5,
    -- filter=58 channel=12
    9, 5, -9, -1, 0, -9, -3, 8, -2,
    -- filter=58 channel=13
    3, 0, -4, -17, -18, 0, -14, -13, 6,
    -- filter=58 channel=14
    -11, 0, -11, 0, 4, 4, -3, 1, 1,
    -- filter=58 channel=15
    -10, -6, -8, 0, -9, 0, -18, -13, 4,
    -- filter=58 channel=16
    0, -16, 1, -9, -17, -3, -17, -13, 3,
    -- filter=58 channel=17
    4, 4, -7, -4, 2, 3, 1, -9, 5,
    -- filter=58 channel=18
    -12, -10, -7, 0, -16, -1, -14, -12, 1,
    -- filter=58 channel=19
    -6, 10, 5, -3, -2, 9, -11, -5, -5,
    -- filter=58 channel=20
    9, -5, 0, -7, 3, 5, -6, -5, 9,
    -- filter=58 channel=21
    3, 0, 9, -8, -9, 0, -6, 8, 7,
    -- filter=58 channel=22
    -9, -10, -3, 0, 9, -7, 0, 0, -6,
    -- filter=58 channel=23
    10, 13, 2, 20, 19, 8, 6, 15, 10,
    -- filter=58 channel=24
    -6, 1, 4, -8, -4, 4, -1, -7, -7,
    -- filter=58 channel=25
    4, 17, 0, 16, 9, 1, 7, 15, 15,
    -- filter=58 channel=26
    -5, 7, 0, 5, 2, 6, 9, 12, 12,
    -- filter=58 channel=27
    8, 5, 9, 17, 19, 6, 9, 9, 3,
    -- filter=58 channel=28
    -1, -15, -6, -16, -12, -11, -16, -19, -4,
    -- filter=58 channel=29
    -19, -7, -11, -22, -10, 5, -10, -11, -13,
    -- filter=58 channel=30
    9, -2, -2, 1, 12, 3, 4, 2, 6,
    -- filter=58 channel=31
    5, 4, -1, -3, 4, 1, 5, 0, -4,
    -- filter=58 channel=32
    19, 24, 17, 21, 25, 22, 23, 25, 16,
    -- filter=58 channel=33
    3, 1, 2, 2, -9, -4, -3, 0, 0,
    -- filter=58 channel=34
    6, 6, 3, 5, -10, 0, 9, -4, 5,
    -- filter=58 channel=35
    26, 33, 12, 18, 33, 12, 22, 28, 13,
    -- filter=58 channel=36
    -2, 0, -1, 5, 11, 6, 4, 15, -2,
    -- filter=58 channel=37
    -5, 2, 7, -8, -10, 4, -1, -6, -3,
    -- filter=58 channel=38
    10, 4, 5, 10, 2, 5, 2, 0, 12,
    -- filter=58 channel=39
    7, 9, -6, -8, 7, -1, -10, -8, -4,
    -- filter=58 channel=40
    -7, 9, 7, 7, -1, 8, -4, -2, 1,
    -- filter=58 channel=41
    0, 5, -4, 0, -10, 7, -10, 3, 13,
    -- filter=58 channel=42
    0, -6, -8, -8, -5, 8, -5, 8, -8,
    -- filter=58 channel=43
    9, 12, 3, 15, 14, 17, -6, 16, 16,
    -- filter=58 channel=44
    14, 3, 3, 15, 2, 3, 7, 8, -4,
    -- filter=58 channel=45
    -9, 0, -3, 0, -4, -2, -4, -9, -6,
    -- filter=58 channel=46
    0, 8, 6, -4, -5, 0, -9, 2, -7,
    -- filter=58 channel=47
    -10, 0, -10, 2, -8, 1, 3, -2, 0,
    -- filter=58 channel=48
    -15, 1, -5, -14, -15, -11, 2, -10, 6,
    -- filter=58 channel=49
    7, 14, 9, 18, 2, 14, 9, 0, 9,
    -- filter=58 channel=50
    3, 9, -5, 3, 0, 5, 1, 6, -2,
    -- filter=58 channel=51
    5, 8, -2, 14, 18, -2, 11, -2, 0,
    -- filter=58 channel=52
    3, -6, 3, 3, -1, 1, -10, -3, 6,
    -- filter=58 channel=53
    -2, 10, 12, 15, 12, 2, 8, 16, 13,
    -- filter=58 channel=54
    -7, 0, -2, -11, 3, 7, -12, -6, 4,
    -- filter=58 channel=55
    -9, 4, 8, 2, -5, 7, 0, -10, -7,
    -- filter=58 channel=56
    4, -4, 5, 5, 3, 2, 9, 1, -3,
    -- filter=58 channel=57
    -7, 6, -3, -3, 0, 2, -7, -6, -6,
    -- filter=58 channel=58
    9, 3, 11, 2, 7, 10, 0, -6, 5,
    -- filter=58 channel=59
    6, 1, -2, 10, 2, 12, -8, -4, 1,
    -- filter=58 channel=60
    -6, -5, -10, -10, -2, -11, -13, -16, 7,
    -- filter=58 channel=61
    0, -11, -4, -1, -2, -5, -5, 3, 1,
    -- filter=58 channel=62
    1, 0, -4, -10, -7, -5, -11, -7, -11,
    -- filter=58 channel=63
    5, 9, 6, -4, -3, -8, -1, -8, -1,
    -- filter=59 channel=0
    -8, 10, -3, 6, -2, 5, 7, 5, 8,
    -- filter=59 channel=1
    -6, -10, -9, -16, -9, 2, -5, 10, -5,
    -- filter=59 channel=2
    1, 2, 1, 5, 0, -9, -1, 4, -1,
    -- filter=59 channel=3
    -5, -2, -1, 16, -5, -7, 8, 5, 7,
    -- filter=59 channel=4
    8, -5, -6, 2, 6, -5, 12, 2, -8,
    -- filter=59 channel=5
    0, 11, 3, -5, 7, -5, 9, 6, 7,
    -- filter=59 channel=6
    4, -9, -8, 6, -8, -4, 0, -7, 5,
    -- filter=59 channel=7
    -2, 0, -8, -7, -3, 8, -8, 5, 4,
    -- filter=59 channel=8
    13, 10, -1, 7, 17, -1, 16, 20, -9,
    -- filter=59 channel=9
    1, -18, -24, -4, -19, -28, 1, -4, -23,
    -- filter=59 channel=10
    -14, 1, 12, 0, 2, 6, -10, 3, -3,
    -- filter=59 channel=11
    -6, 6, -2, 2, 10, -9, 0, 5, 3,
    -- filter=59 channel=12
    -3, -9, -9, 9, -2, 0, -7, 8, 1,
    -- filter=59 channel=13
    13, -10, -7, 6, 9, -17, 7, 12, -13,
    -- filter=59 channel=14
    8, -8, -8, 0, 2, 11, 5, 6, 7,
    -- filter=59 channel=15
    -1, 4, -11, 13, 13, -7, 12, 12, 3,
    -- filter=59 channel=16
    17, 0, -11, 24, 11, -2, 0, 10, -7,
    -- filter=59 channel=17
    5, 2, -3, 12, 15, -2, 0, 6, 12,
    -- filter=59 channel=18
    -5, 0, 7, 11, 2, -2, 1, 1, -7,
    -- filter=59 channel=19
    -1, -3, -3, 1, -4, -1, 4, -11, -4,
    -- filter=59 channel=20
    -8, -4, 0, -2, -14, -1, -13, 0, 0,
    -- filter=59 channel=21
    1, 9, -5, 7, 10, 4, 10, 3, -1,
    -- filter=59 channel=22
    3, -7, -4, 6, 2, 4, -8, 7, 0,
    -- filter=59 channel=23
    -12, -2, 8, 0, 4, 0, 6, 3, 15,
    -- filter=59 channel=24
    9, -7, -13, 7, 13, 7, 0, 8, 5,
    -- filter=59 channel=25
    9, -5, 4, -10, -10, -4, -8, 9, -9,
    -- filter=59 channel=26
    -14, -4, -9, -1, -8, -11, -10, -2, 0,
    -- filter=59 channel=27
    10, 0, 1, -2, 2, 3, 0, 5, 3,
    -- filter=59 channel=28
    0, 9, -2, 5, 3, -4, 5, 4, -13,
    -- filter=59 channel=29
    18, -8, -12, 5, 5, -8, 7, -6, -22,
    -- filter=59 channel=30
    -13, -1, -4, -19, -8, 7, -10, 6, 10,
    -- filter=59 channel=31
    -7, 4, -1, -10, -2, 5, -10, 8, 5,
    -- filter=59 channel=32
    -13, 1, -3, -14, -7, 3, -10, -8, 11,
    -- filter=59 channel=33
    0, -9, 2, -2, -6, -4, -4, 3, -10,
    -- filter=59 channel=34
    1, -11, -1, 6, -8, -3, -5, -9, 8,
    -- filter=59 channel=35
    0, 13, 13, 0, 7, 2, -9, -1, 8,
    -- filter=59 channel=36
    -9, 0, 7, -5, -6, 0, -2, -10, -9,
    -- filter=59 channel=37
    4, -6, -4, 2, -3, -7, 8, -1, -10,
    -- filter=59 channel=38
    1, 5, -5, -3, 12, -6, 14, 13, -3,
    -- filter=59 channel=39
    8, 3, -7, 0, 5, 9, 9, -4, -5,
    -- filter=59 channel=40
    -10, 2, -7, -9, -6, 0, -1, -9, -1,
    -- filter=59 channel=41
    0, 5, -14, 12, 19, -9, 2, 12, 0,
    -- filter=59 channel=42
    2, 9, 1, 4, -5, -3, -3, 2, 9,
    -- filter=59 channel=43
    -22, -20, -11, -29, -31, -20, -16, -15, -7,
    -- filter=59 channel=44
    -5, -8, -8, -13, -6, 9, -7, 0, 6,
    -- filter=59 channel=45
    0, 1, -2, -3, -8, 3, 0, -5, 4,
    -- filter=59 channel=46
    1, -3, 1, -3, -7, 6, 6, -14, 4,
    -- filter=59 channel=47
    -10, 4, -5, -1, 7, 3, 3, 2, -1,
    -- filter=59 channel=48
    6, -11, -3, 0, -11, 3, 2, -3, -6,
    -- filter=59 channel=49
    2, 13, -3, 4, 9, -2, -10, 15, -1,
    -- filter=59 channel=50
    -5, -5, 0, -4, -13, -13, -5, -8, -5,
    -- filter=59 channel=51
    6, 3, 9, 5, 14, 10, -9, 17, 12,
    -- filter=59 channel=52
    -4, 4, -8, 1, 10, 10, -7, 10, 8,
    -- filter=59 channel=53
    0, -5, -4, -5, -5, -1, -15, 7, 10,
    -- filter=59 channel=54
    -14, -1, -16, 0, -18, -23, -11, -5, -21,
    -- filter=59 channel=55
    -7, 6, -2, -1, -4, 8, 4, 10, 3,
    -- filter=59 channel=56
    -10, -11, 0, -10, -9, -8, 6, -4, -3,
    -- filter=59 channel=57
    -6, 4, 0, -4, -10, 9, 5, 2, 2,
    -- filter=59 channel=58
    -6, -8, 5, -6, -2, 0, -7, -7, 7,
    -- filter=59 channel=59
    9, 10, 0, 9, 0, -3, 3, 4, -2,
    -- filter=59 channel=60
    15, 12, -17, 27, 25, 1, 9, 20, -5,
    -- filter=59 channel=61
    6, 2, -11, 12, 8, 0, 0, 16, 4,
    -- filter=59 channel=62
    0, 6, 6, 13, 2, -2, 11, -4, -4,
    -- filter=59 channel=63
    1, 5, 0, 5, -4, -9, 5, 0, -9,
    -- filter=60 channel=0
    10, -3, -1, -9, 6, 11, 8, -3, 2,
    -- filter=60 channel=1
    7, 7, -5, -6, 1, 3, -4, 0, 2,
    -- filter=60 channel=2
    2, 5, -5, 7, -7, 10, -5, 5, -7,
    -- filter=60 channel=3
    0, 3, 8, -4, -8, -9, 1, -5, 4,
    -- filter=60 channel=4
    -3, 8, -8, 0, 4, -3, 0, 0, 8,
    -- filter=60 channel=5
    4, 8, 7, -2, 2, 4, -1, -4, -7,
    -- filter=60 channel=6
    -5, 8, -7, -1, 9, 2, 8, 7, 11,
    -- filter=60 channel=7
    8, 4, 5, 0, -7, -8, 6, -4, 6,
    -- filter=60 channel=8
    -3, -1, 4, -1, 0, -10, -9, 0, 7,
    -- filter=60 channel=9
    -1, -2, -1, -5, -5, 0, -8, 9, 2,
    -- filter=60 channel=10
    11, -2, 0, -1, 5, -2, 2, 1, 4,
    -- filter=60 channel=11
    0, 5, 0, -2, 0, -10, -3, 3, 1,
    -- filter=60 channel=12
    6, -5, -7, -5, 3, -1, 2, 2, -10,
    -- filter=60 channel=13
    10, 10, -4, 10, 8, 7, -8, -8, 5,
    -- filter=60 channel=14
    1, -2, -6, 8, 2, -2, 8, 2, 6,
    -- filter=60 channel=15
    -10, -3, 2, 0, 0, -2, -8, 7, -5,
    -- filter=60 channel=16
    1, -9, -7, -2, 0, -7, -6, 8, 7,
    -- filter=60 channel=17
    -9, 0, 9, -2, -1, -4, -6, -3, 0,
    -- filter=60 channel=18
    0, -5, 9, -7, -3, 0, 9, -7, 8,
    -- filter=60 channel=19
    -4, 1, -5, 1, 0, -7, -4, 5, -4,
    -- filter=60 channel=20
    1, -6, -6, 1, 1, -3, 8, -5, -9,
    -- filter=60 channel=21
    0, -8, 8, -8, 9, 0, 5, 6, 8,
    -- filter=60 channel=22
    0, 0, -1, -2, 0, 10, 9, 0, 3,
    -- filter=60 channel=23
    6, 8, 1, -7, 4, 5, 1, 7, 0,
    -- filter=60 channel=24
    1, -6, 4, -5, 3, 10, 0, 3, -7,
    -- filter=60 channel=25
    7, -8, -7, -9, -8, -1, -2, 0, -6,
    -- filter=60 channel=26
    4, -7, 10, 7, -6, -6, -7, 6, 0,
    -- filter=60 channel=27
    -8, -5, 0, -1, 1, 6, -3, 10, 3,
    -- filter=60 channel=28
    5, 8, 10, 3, 0, 1, -8, 0, 4,
    -- filter=60 channel=29
    -3, -4, -8, -8, 8, -6, 9, 6, -7,
    -- filter=60 channel=30
    -2, -7, 9, 11, 0, -1, 0, -4, 3,
    -- filter=60 channel=31
    4, 1, -6, -7, 1, -8, -1, -9, 1,
    -- filter=60 channel=32
    8, 4, 0, 4, 4, 1, -8, 9, -8,
    -- filter=60 channel=33
    10, -9, 4, 0, 0, 8, 6, 0, -7,
    -- filter=60 channel=34
    2, -5, 5, -1, 10, 3, 0, -9, 2,
    -- filter=60 channel=35
    3, -3, 8, 0, -5, 9, 4, 5, 5,
    -- filter=60 channel=36
    -6, -5, -8, -4, -8, -3, 9, 0, 3,
    -- filter=60 channel=37
    -4, 7, 6, 0, 0, -4, -8, -6, 3,
    -- filter=60 channel=38
    -5, -6, -3, -6, 6, 8, -9, 4, -9,
    -- filter=60 channel=39
    8, 0, 5, -5, 3, 3, -1, -3, 1,
    -- filter=60 channel=40
    10, 0, 2, -6, 4, -8, 7, -9, 0,
    -- filter=60 channel=41
    -5, 2, -1, -10, 2, -8, 0, -6, 2,
    -- filter=60 channel=42
    1, -1, -9, -8, 3, 9, 0, 4, 3,
    -- filter=60 channel=43
    0, -1, -3, -6, 1, 9, -1, -5, -4,
    -- filter=60 channel=44
    7, -7, 3, 8, -8, 5, -8, -8, 4,
    -- filter=60 channel=45
    0, 6, -10, 3, -4, -1, 1, 10, 0,
    -- filter=60 channel=46
    8, 5, 10, -4, 8, 1, 10, -8, 8,
    -- filter=60 channel=47
    -8, 4, 1, -7, -3, 2, 6, 0, 1,
    -- filter=60 channel=48
    7, -4, -1, 2, -5, -2, 8, -2, -7,
    -- filter=60 channel=49
    4, -8, 0, 8, 6, -2, -8, -7, 4,
    -- filter=60 channel=50
    0, 7, 7, -8, -10, -5, -10, -4, 5,
    -- filter=60 channel=51
    -4, 2, -2, 12, 10, 10, 6, -1, 6,
    -- filter=60 channel=52
    -4, -2, -3, 0, -5, 8, 1, -4, 10,
    -- filter=60 channel=53
    -4, -8, -1, 11, 2, 10, 8, 10, 10,
    -- filter=60 channel=54
    -3, -10, -3, 7, -2, 8, 8, 6, 6,
    -- filter=60 channel=55
    3, -7, 10, 9, 8, 1, 0, 4, 1,
    -- filter=60 channel=56
    -4, 8, -10, 4, 9, -9, -4, 8, 7,
    -- filter=60 channel=57
    -10, 7, -2, -7, 8, 4, 1, 2, -8,
    -- filter=60 channel=58
    11, 10, 8, -7, 7, 7, 9, -6, 1,
    -- filter=60 channel=59
    2, -9, 1, 6, 8, 5, -4, 0, 9,
    -- filter=60 channel=60
    3, 0, -8, -3, -10, -7, 0, -2, 0,
    -- filter=60 channel=61
    -6, -9, -3, 9, 0, -5, 9, -6, 6,
    -- filter=60 channel=62
    8, 10, -10, 0, -5, -2, 1, 9, 5,
    -- filter=60 channel=63
    9, 6, 7, -9, 0, 7, 7, 2, 1,
    -- filter=61 channel=0
    -7, 2, -4, 1, 16, 13, -1, 7, 1,
    -- filter=61 channel=1
    -6, 2, -8, 0, -1, 5, -19, -4, 7,
    -- filter=61 channel=2
    -15, -11, -2, -5, -5, -5, -11, -7, -4,
    -- filter=61 channel=3
    -2, 3, -10, -14, -3, -5, -12, 5, -5,
    -- filter=61 channel=4
    10, 5, 12, -6, -4, 9, -5, 5, 9,
    -- filter=61 channel=5
    -7, 10, 5, 5, -5, 14, -7, 1, 3,
    -- filter=61 channel=6
    -6, -2, -7, -1, 2, -10, 1, 5, -10,
    -- filter=61 channel=7
    8, 0, -5, 12, 0, 3, 0, 13, 10,
    -- filter=61 channel=8
    0, 0, 8, -5, 16, 14, 8, 8, -4,
    -- filter=61 channel=9
    5, -8, -1, 10, 5, -5, 4, 12, 5,
    -- filter=61 channel=10
    9, -9, 7, 3, 2, 6, -7, -6, 5,
    -- filter=61 channel=11
    1, 0, -2, -12, 6, 12, -7, -3, -2,
    -- filter=61 channel=12
    -3, -2, 4, 1, -5, -9, -10, 7, -9,
    -- filter=61 channel=13
    -1, 1, -7, 4, 3, 1, -1, 12, 7,
    -- filter=61 channel=14
    11, 8, 14, 8, 13, 16, -2, 10, 12,
    -- filter=61 channel=15
    -8, 6, -2, -11, 12, 4, 1, 11, -9,
    -- filter=61 channel=16
    3, -2, -8, 1, -8, -10, 0, -4, 7,
    -- filter=61 channel=17
    -9, 3, -5, -1, -1, 2, -10, 12, 10,
    -- filter=61 channel=18
    12, 0, 7, 9, 3, 5, 5, 2, -2,
    -- filter=61 channel=19
    3, 3, 3, 4, -12, -6, -6, -8, -4,
    -- filter=61 channel=20
    -6, 12, 11, 13, 0, -2, -3, 1, 11,
    -- filter=61 channel=21
    0, 5, 7, -7, -7, 9, -8, 9, 6,
    -- filter=61 channel=22
    8, -5, 0, 4, 5, -2, 4, -8, 10,
    -- filter=61 channel=23
    0, -6, -3, -1, 4, -5, -7, 0, 8,
    -- filter=61 channel=24
    10, 3, 0, -6, 6, 2, 0, -4, -2,
    -- filter=61 channel=25
    -4, -18, -8, -22, -13, -4, -18, -14, -19,
    -- filter=61 channel=26
    -5, 5, 6, 10, 4, 1, -3, -1, 0,
    -- filter=61 channel=27
    -6, -6, -6, -16, -9, 3, -17, 3, 10,
    -- filter=61 channel=28
    8, 4, -6, 4, -7, -9, 0, 0, 10,
    -- filter=61 channel=29
    -12, -1, 2, -8, 13, -14, 1, 17, 3,
    -- filter=61 channel=30
    3, 8, 13, 4, 1, 28, 21, 11, 28,
    -- filter=61 channel=31
    0, 8, 10, -10, -9, 7, 7, 3, -4,
    -- filter=61 channel=32
    9, 1, 4, 1, -8, 0, 6, -2, -2,
    -- filter=61 channel=33
    -6, -4, -9, -8, 2, 5, -3, -8, -7,
    -- filter=61 channel=34
    -3, 14, 3, 4, -1, 5, 3, 11, 0,
    -- filter=61 channel=35
    -12, -4, -5, -11, 0, -6, -14, 0, -9,
    -- filter=61 channel=36
    -6, 7, 7, -7, -6, -5, 5, -6, -5,
    -- filter=61 channel=37
    1, -9, -11, -3, 0, 7, -3, -7, -7,
    -- filter=61 channel=38
    4, -2, -11, 0, 9, -4, -13, -3, 9,
    -- filter=61 channel=39
    -6, -4, -5, -9, 0, 3, -6, -10, 1,
    -- filter=61 channel=40
    -10, -1, 10, 3, 8, 6, 6, -8, 4,
    -- filter=61 channel=41
    -13, -4, 1, -8, 5, 6, -6, 8, 4,
    -- filter=61 channel=42
    0, 10, 2, -2, -8, -1, -1, 7, 0,
    -- filter=61 channel=43
    -8, -10, -5, -6, -12, -1, -4, -5, 1,
    -- filter=61 channel=44
    -8, -9, 8, 1, -2, 12, 10, 3, -3,
    -- filter=61 channel=45
    9, 7, 4, 9, 4, -3, -7, 0, 0,
    -- filter=61 channel=46
    -6, 2, 1, 4, 10, -1, 13, 6, 6,
    -- filter=61 channel=47
    -6, -3, 0, 2, 0, -2, 9, 0, 6,
    -- filter=61 channel=48
    -11, -3, -1, -6, -7, -11, 3, 12, -6,
    -- filter=61 channel=49
    0, 10, -5, 3, 1, -3, 6, 6, 2,
    -- filter=61 channel=50
    10, -2, -2, 1, 0, 12, 6, 8, 0,
    -- filter=61 channel=51
    -3, 11, 2, 9, 6, 0, 13, 4, 10,
    -- filter=61 channel=52
    6, -5, 3, 2, -2, -3, 0, -4, -3,
    -- filter=61 channel=53
    10, 7, 7, 10, -4, 20, 10, -6, 13,
    -- filter=61 channel=54
    4, -2, 5, -1, 9, 13, 3, 13, 14,
    -- filter=61 channel=55
    1, -2, 8, -8, -8, 4, -6, 3, -10,
    -- filter=61 channel=56
    11, 7, 2, 11, -1, 5, 10, 12, 13,
    -- filter=61 channel=57
    10, -5, 1, 7, 9, -1, -2, 6, 4,
    -- filter=61 channel=58
    6, -4, -10, 7, -1, -10, 1, 5, -11,
    -- filter=61 channel=59
    -11, 2, -11, -14, 10, 5, -13, -7, -6,
    -- filter=61 channel=60
    -3, 16, 3, -10, 18, 10, 0, 17, 0,
    -- filter=61 channel=61
    1, 13, 14, -4, 5, 12, -5, 17, 18,
    -- filter=61 channel=62
    -6, 2, 0, -5, -9, -10, -10, -8, 9,
    -- filter=61 channel=63
    1, -4, 4, 9, 5, -1, -9, 0, 2,
    -- filter=62 channel=0
    0, -3, -3, 10, -10, 0, 5, 2, 1,
    -- filter=62 channel=1
    -9, -7, -6, 5, -8, -5, 9, -5, -8,
    -- filter=62 channel=2
    1, -2, 3, -7, -6, 1, -2, 8, -3,
    -- filter=62 channel=3
    4, 9, 9, 2, -6, 2, 2, 9, 0,
    -- filter=62 channel=4
    5, -4, -1, 9, 8, -8, -1, -1, -6,
    -- filter=62 channel=5
    -5, 0, -4, -3, 2, 0, 7, -4, -5,
    -- filter=62 channel=6
    -1, 0, 5, -1, -4, 0, -9, -8, 9,
    -- filter=62 channel=7
    -1, 0, 0, -4, -5, -3, 6, 11, -8,
    -- filter=62 channel=8
    6, -1, 5, 2, -3, -10, 2, -12, -11,
    -- filter=62 channel=9
    -2, 11, 1, 7, 9, 4, -8, 3, 9,
    -- filter=62 channel=10
    0, -8, 0, -4, 8, 5, -8, 1, 7,
    -- filter=62 channel=11
    8, -5, 1, 2, -7, -3, 7, 1, -12,
    -- filter=62 channel=12
    0, -6, -3, -6, -9, -1, -9, -3, -8,
    -- filter=62 channel=13
    7, 3, 5, -6, 10, -9, -6, -9, 5,
    -- filter=62 channel=14
    -7, 8, -6, -6, 7, -8, -7, -7, -4,
    -- filter=62 channel=15
    4, 8, -4, 2, -3, 7, -8, -1, -7,
    -- filter=62 channel=16
    -7, -1, 11, 9, -2, -3, 0, 1, -8,
    -- filter=62 channel=17
    -2, -4, 0, 2, -3, -6, -9, 7, 5,
    -- filter=62 channel=18
    3, -8, 7, -4, 3, 3, -9, 7, -2,
    -- filter=62 channel=19
    -7, -1, 0, -10, -4, 9, -2, -10, 8,
    -- filter=62 channel=20
    -3, 7, 9, 6, 7, -8, -1, -8, 5,
    -- filter=62 channel=21
    -7, 9, -9, 4, 8, 10, -7, 6, 0,
    -- filter=62 channel=22
    -9, 8, -8, 1, 5, -3, 8, -10, 5,
    -- filter=62 channel=23
    1, -9, 1, -10, -4, -4, 2, 2, -7,
    -- filter=62 channel=24
    7, 6, -6, 7, 4, -7, 8, 7, -10,
    -- filter=62 channel=25
    10, 10, 4, 5, -2, -6, -7, 2, -1,
    -- filter=62 channel=26
    8, -9, 0, 4, 2, -1, 4, 0, -7,
    -- filter=62 channel=27
    -3, -7, 6, -6, -6, -10, 0, -11, 8,
    -- filter=62 channel=28
    -2, -6, -7, -8, -9, -8, 0, -5, 0,
    -- filter=62 channel=29
    14, 12, 7, 3, 1, -5, 8, -5, -2,
    -- filter=62 channel=30
    -2, 7, -7, -2, -5, -3, 0, 1, 3,
    -- filter=62 channel=31
    -3, 4, -8, -2, 4, -9, 7, 4, -2,
    -- filter=62 channel=32
    0, 8, -2, 7, 2, 3, -1, -8, 7,
    -- filter=62 channel=33
    1, 5, 4, -10, -9, -2, -7, 8, -2,
    -- filter=62 channel=34
    -7, 3, -9, 10, 1, -8, 2, -6, 7,
    -- filter=62 channel=35
    2, 0, 0, -5, -2, -11, -8, 7, 2,
    -- filter=62 channel=36
    -2, -8, -8, -6, -2, -1, 0, 5, -8,
    -- filter=62 channel=37
    -9, -3, 7, -9, 5, 7, 4, 8, -5,
    -- filter=62 channel=38
    -7, 11, 12, 9, -10, -1, 0, -9, -2,
    -- filter=62 channel=39
    -7, -1, 4, 1, -3, 1, 5, -2, 3,
    -- filter=62 channel=40
    -10, 0, 9, 6, 0, -3, 8, -2, 1,
    -- filter=62 channel=41
    -4, 0, -5, 5, -9, -11, -8, 0, -2,
    -- filter=62 channel=42
    -2, -2, 0, 4, -2, 6, 7, 3, -4,
    -- filter=62 channel=43
    4, -5, 10, -3, -3, 1, 5, 6, -7,
    -- filter=62 channel=44
    8, -7, 6, 1, 10, 3, 10, 8, 0,
    -- filter=62 channel=45
    -7, -4, 0, 3, -4, 7, 1, -3, 4,
    -- filter=62 channel=46
    12, 0, 6, 1, 9, -4, 3, 0, 12,
    -- filter=62 channel=47
    -8, -8, 1, -2, -9, -10, 4, 4, 7,
    -- filter=62 channel=48
    0, -6, 0, 0, -10, 8, -4, 2, 6,
    -- filter=62 channel=49
    -7, -8, -10, -8, -4, -3, 2, 6, 8,
    -- filter=62 channel=50
    -2, -3, 6, -8, 7, 8, 11, 8, -2,
    -- filter=62 channel=51
    9, 0, -10, -8, 5, 2, 4, 4, 4,
    -- filter=62 channel=52
    -2, 2, -6, 4, 4, 8, 10, 9, 1,
    -- filter=62 channel=53
    2, 2, 0, -6, 7, -7, -8, -4, 9,
    -- filter=62 channel=54
    8, 8, 0, -8, 1, 4, 7, 8, -7,
    -- filter=62 channel=55
    4, 3, -8, 6, -7, -7, 7, 4, 5,
    -- filter=62 channel=56
    -5, 7, 3, 0, -4, -6, 1, -1, 4,
    -- filter=62 channel=57
    -6, -2, -5, 6, -2, 5, -8, -10, -7,
    -- filter=62 channel=58
    8, 4, -4, 0, 9, 4, 0, -1, 3,
    -- filter=62 channel=59
    7, -7, -2, -8, 7, 3, 0, -6, 0,
    -- filter=62 channel=60
    12, 13, 13, 7, 6, 8, -8, 1, 4,
    -- filter=62 channel=61
    4, 3, -5, 3, -3, -7, 8, 1, -7,
    -- filter=62 channel=62
    6, 5, 4, 0, -4, 0, -4, 4, 5,
    -- filter=62 channel=63
    4, -6, 3, -8, -3, 8, -9, -7, -8,
    -- filter=63 channel=0
    1, 7, 13, 12, 11, 18, 13, 5, 15,
    -- filter=63 channel=1
    7, 11, 3, -4, -2, 7, 10, 6, 10,
    -- filter=63 channel=2
    -6, -4, 6, -5, 7, -4, 1, 6, -8,
    -- filter=63 channel=3
    -5, -2, -7, 7, -11, -7, -10, 4, -1,
    -- filter=63 channel=4
    10, 2, -8, 8, 9, -8, 8, -10, -3,
    -- filter=63 channel=5
    -1, -8, -10, 3, 0, -5, 4, -9, -5,
    -- filter=63 channel=6
    9, -6, 1, 3, 7, -8, 9, 5, -1,
    -- filter=63 channel=7
    -1, -3, 4, 2, -8, 7, 8, 2, -5,
    -- filter=63 channel=8
    -11, 7, 4, 7, 7, -1, -14, -5, -15,
    -- filter=63 channel=9
    5, 4, 9, -12, 0, 4, -12, 0, 3,
    -- filter=63 channel=10
    9, 24, 15, 23, 11, 12, 18, 17, 19,
    -- filter=63 channel=11
    -7, -2, 2, 6, 10, -2, 8, 0, -10,
    -- filter=63 channel=12
    5, 6, 5, 0, 2, 4, -9, -3, 8,
    -- filter=63 channel=13
    -2, -5, -4, -11, -2, -7, -12, 1, -1,
    -- filter=63 channel=14
    -1, 7, 9, 10, 0, 11, -8, 3, -5,
    -- filter=63 channel=15
    3, 0, -13, -4, -3, 0, 2, -8, -2,
    -- filter=63 channel=16
    -16, -16, 0, -20, -9, -15, -9, -18, -18,
    -- filter=63 channel=17
    -11, 8, 7, 3, 3, -2, 3, -11, -4,
    -- filter=63 channel=18
    11, 0, 2, -7, 7, 8, 0, -5, -3,
    -- filter=63 channel=19
    6, 1, 4, 3, 3, -4, -9, -11, -2,
    -- filter=63 channel=20
    -9, -3, -6, 0, 3, -3, 2, 7, 6,
    -- filter=63 channel=21
    8, 1, -9, -5, -8, 1, 0, -7, -1,
    -- filter=63 channel=22
    -10, 2, 9, 2, -1, -5, 0, 0, 3,
    -- filter=63 channel=23
    16, 27, 15, 24, 20, 14, 14, 21, 8,
    -- filter=63 channel=24
    0, -9, -3, 7, 5, -6, -3, -2, 6,
    -- filter=63 channel=25
    3, 0, 8, 4, -2, -2, 15, 11, 6,
    -- filter=63 channel=26
    2, -7, 4, 10, 3, -8, 3, -4, 4,
    -- filter=63 channel=27
    15, 1, 10, 0, 17, 1, 1, 8, -3,
    -- filter=63 channel=28
    -19, -16, -3, -19, -15, -20, -5, -16, -17,
    -- filter=63 channel=29
    -24, -6, -6, -24, -10, -23, -7, -23, -22,
    -- filter=63 channel=30
    8, 11, 11, 5, 9, 0, -5, 12, 2,
    -- filter=63 channel=31
    11, 2, 0, 12, 14, -3, 2, -3, 5,
    -- filter=63 channel=32
    10, 15, 7, 7, 15, 6, 16, 12, 20,
    -- filter=63 channel=33
    -1, 2, 4, 9, -2, -7, -9, -6, -4,
    -- filter=63 channel=34
    3, -1, -4, 0, 0, 8, -8, -3, 0,
    -- filter=63 channel=35
    15, 17, 24, 21, 38, 13, 11, 28, 27,
    -- filter=63 channel=36
    0, -2, -4, 3, 11, 6, 8, 0, 8,
    -- filter=63 channel=37
    -10, 8, 1, -5, 4, -11, -12, 0, 7,
    -- filter=63 channel=38
    -4, 14, -2, 7, 0, 4, 2, -1, -3,
    -- filter=63 channel=39
    -1, -5, -10, 3, 5, 3, 3, 10, 8,
    -- filter=63 channel=40
    -1, 11, 7, -3, 6, -5, 3, 9, 7,
    -- filter=63 channel=41
    -1, 0, -9, -1, 5, -5, 0, 7, 0,
    -- filter=63 channel=42
    10, -7, -7, 0, 0, 7, -7, 1, -8,
    -- filter=63 channel=43
    2, 5, 2, -11, -5, -10, -4, -9, -2,
    -- filter=63 channel=44
    13, 12, -1, 10, 0, -1, 5, 7, -3,
    -- filter=63 channel=45
    5, 9, 0, 4, -8, -8, 9, -3, 5,
    -- filter=63 channel=46
    6, -7, 4, 0, 1, 3, 1, 8, 6,
    -- filter=63 channel=47
    3, -3, -3, 2, -9, 9, -5, -3, -6,
    -- filter=63 channel=48
    -9, -7, -1, 0, -8, -13, -8, -14, 0,
    -- filter=63 channel=49
    14, 3, 12, 5, 17, 18, 11, 21, 4,
    -- filter=63 channel=50
    -8, -1, -6, 5, -7, -6, -8, -10, 9,
    -- filter=63 channel=51
    4, 13, 6, 11, 17, 20, 21, 23, 21,
    -- filter=63 channel=52
    -3, -3, 9, 3, 4, -2, 9, -4, 6,
    -- filter=63 channel=53
    12, -2, 14, 5, 3, 1, 0, 9, -1,
    -- filter=63 channel=54
    4, 5, 5, -7, -9, 3, -5, 8, 1,
    -- filter=63 channel=55
    0, -7, 3, -2, 10, 4, -1, -9, 8,
    -- filter=63 channel=56
    -5, -6, -6, -8, 3, 1, 10, -5, 10,
    -- filter=63 channel=57
    -4, 0, -4, 4, -7, -4, 6, 4, -3,
    -- filter=63 channel=58
    7, 8, 2, 1, 4, 7, 3, 3, -6,
    -- filter=63 channel=59
    -1, -8, -10, -9, -6, 9, -3, 3, -3,
    -- filter=63 channel=60
    4, -5, -9, -7, 4, -9, -10, -12, -2,
    -- filter=63 channel=61
    -1, -1, 10, 10, 10, 10, 9, 3, 9,
    -- filter=63 channel=62
    -3, -3, 4, -1, -3, -10, -7, -9, 7,
    -- filter=63 channel=63
    8, -1, 0, 4, 7, 2, 6, -5, 3,
    -- filter=64 channel=0
    -1, -5, 2, 2, -5, -3, -3, 7, 9,
    -- filter=64 channel=1
    -2, -11, -12, -4, -12, -11, -9, -3, -15,
    -- filter=64 channel=2
    -11, -12, -10, 7, -13, 2, 4, -13, -6,
    -- filter=64 channel=3
    -12, -7, -12, 2, -12, 4, -1, 1, -10,
    -- filter=64 channel=4
    10, 6, 4, 11, 5, 2, -2, 9, -2,
    -- filter=64 channel=5
    0, -4, 4, -5, 4, 0, 3, 8, 5,
    -- filter=64 channel=6
    -2, 10, 0, 11, -1, -7, 9, -8, 8,
    -- filter=64 channel=7
    11, -3, -6, -5, -4, 8, -6, 9, 10,
    -- filter=64 channel=8
    -6, 2, 10, 0, 0, 5, -4, 9, 13,
    -- filter=64 channel=9
    3, 9, 6, -1, 0, 9, 14, 21, 13,
    -- filter=64 channel=10
    12, 6, 11, 6, 6, 10, -6, -5, -2,
    -- filter=64 channel=11
    -4, 8, -8, 10, -4, 5, -6, -9, -1,
    -- filter=64 channel=12
    -2, -1, -7, 9, -1, -6, 7, -6, 10,
    -- filter=64 channel=13
    -7, 0, 13, 7, 13, 5, 3, 10, 2,
    -- filter=64 channel=14
    -8, -4, 7, 0, 9, -2, 10, 7, -4,
    -- filter=64 channel=15
    4, -6, 2, 9, 3, -1, 0, 1, 11,
    -- filter=64 channel=16
    0, -6, -9, 4, 0, 4, -11, -10, 0,
    -- filter=64 channel=17
    -1, 11, 0, 2, 4, -8, -4, -1, -6,
    -- filter=64 channel=18
    17, 7, 15, 13, 18, 20, 2, 21, 21,
    -- filter=64 channel=19
    -2, 0, -9, -2, 5, 4, -2, -1, -1,
    -- filter=64 channel=20
    -5, 1, -1, -6, -3, 4, 0, 14, -2,
    -- filter=64 channel=21
    -9, -7, 4, 0, 8, 7, -9, 10, 7,
    -- filter=64 channel=22
    -6, 9, 6, 5, 5, 4, -3, 0, 10,
    -- filter=64 channel=23
    9, 0, -5, 0, -7, 2, -6, -4, -8,
    -- filter=64 channel=24
    -7, -4, -9, -5, 6, -5, 9, 7, -1,
    -- filter=64 channel=25
    -13, -16, -12, -8, -19, -15, -16, -13, -11,
    -- filter=64 channel=26
    3, -7, -2, -5, -7, -1, -7, -3, -5,
    -- filter=64 channel=27
    7, -4, -11, -10, -15, 2, -10, -2, 5,
    -- filter=64 channel=28
    12, 0, 11, 0, 6, -4, 4, 6, 7,
    -- filter=64 channel=29
    6, 3, -1, -3, -8, 13, -4, 1, 10,
    -- filter=64 channel=30
    -6, 4, -3, 7, 12, -4, 9, 1, 13,
    -- filter=64 channel=31
    -8, -8, 10, -4, -7, 1, 5, 5, 2,
    -- filter=64 channel=32
    2, -11, -2, -13, -5, -2, 2, -5, -2,
    -- filter=64 channel=33
    8, -7, -3, -1, -9, 9, 0, 9, 4,
    -- filter=64 channel=34
    6, -6, -8, 0, -5, 13, 9, 6, 13,
    -- filter=64 channel=35
    -3, 0, -1, -4, -14, 3, 5, -13, 0,
    -- filter=64 channel=36
    -4, 7, 10, 4, -6, 3, 8, -1, 6,
    -- filter=64 channel=37
    0, -6, -3, -6, -7, -8, 4, -8, 5,
    -- filter=64 channel=38
    -5, -5, -8, 8, -5, -8, -1, -12, 2,
    -- filter=64 channel=39
    6, -4, -7, -8, 6, 1, 4, -1, 7,
    -- filter=64 channel=40
    8, -9, -7, 10, -11, -4, -9, 0, 0,
    -- filter=64 channel=41
    5, 7, 5, 3, -6, 8, 5, -2, 9,
    -- filter=64 channel=42
    7, 4, 0, 3, 5, 7, -5, -9, -8,
    -- filter=64 channel=43
    6, 0, -7, -4, -6, -1, 14, 9, -8,
    -- filter=64 channel=44
    0, 0, -10, 7, -9, -7, -3, -6, -7,
    -- filter=64 channel=45
    3, 9, 2, -9, -9, -1, 6, 2, 5,
    -- filter=64 channel=46
    -6, 1, 12, 8, -5, -5, -2, -5, 8,
    -- filter=64 channel=47
    5, 4, 4, -1, -4, -3, -7, 10, 0,
    -- filter=64 channel=48
    4, -9, -6, 3, 0, 4, 5, 8, 7,
    -- filter=64 channel=49
    1, 2, 7, 5, -3, -7, -4, -7, 0,
    -- filter=64 channel=50
    -2, 9, 1, 6, -3, 7, 13, -3, -4,
    -- filter=64 channel=51
    -1, 16, 14, 0, 6, 15, 9, 2, 3,
    -- filter=64 channel=52
    -5, -6, 4, -4, 5, 5, 2, -7, 1,
    -- filter=64 channel=53
    -7, 12, 5, 5, -3, -11, -2, 8, 5,
    -- filter=64 channel=54
    0, 8, -4, 11, 0, -6, 0, 2, -5,
    -- filter=64 channel=55
    -6, 3, 9, 8, -4, 7, 6, -2, 1,
    -- filter=64 channel=56
    10, 8, 8, -7, 2, 11, 9, -7, 2,
    -- filter=64 channel=57
    7, 0, -5, -5, 5, -3, -1, 6, 0,
    -- filter=64 channel=58
    0, 8, -1, 11, -1, 11, 7, 3, 9,
    -- filter=64 channel=59
    -8, -15, -8, -4, 2, 1, -10, -4, -5,
    -- filter=64 channel=60
    8, -5, 9, 2, 8, -5, 7, 5, -1,
    -- filter=64 channel=61
    -4, 10, -6, 7, 0, 9, -7, 9, 0,
    -- filter=64 channel=62
    -9, -4, -9, -7, 4, -8, -1, -11, -9,
    -- filter=64 channel=63
    0, 10, -5, -2, -1, 3, -2, 9, -7,
    -- filter=65 channel=0
    -6, -2, -4, 0, -1, -1, 6, -10, -1,
    -- filter=65 channel=1
    1, 0, 10, -1, -4, 1, -4, -1, -1,
    -- filter=65 channel=2
    -10, -2, 6, 3, -4, 5, -4, 0, -4,
    -- filter=65 channel=3
    -4, 5, 4, 7, 0, -7, -8, -1, -9,
    -- filter=65 channel=4
    -9, -9, 8, 3, -6, -10, -2, -6, -5,
    -- filter=65 channel=5
    0, 0, 6, -1, -7, 2, -6, 4, -10,
    -- filter=65 channel=6
    2, -1, -10, 6, -9, -4, 4, -7, 0,
    -- filter=65 channel=7
    -8, -7, 4, 2, 2, 1, 0, 7, -6,
    -- filter=65 channel=8
    -4, 4, 0, -5, 0, 3, -8, 2, -5,
    -- filter=65 channel=9
    9, 0, 9, 9, 4, -6, -8, -3, -8,
    -- filter=65 channel=10
    0, -2, -9, -4, -6, 2, -8, 8, -5,
    -- filter=65 channel=11
    4, -1, 6, 9, 6, 4, 1, -5, 1,
    -- filter=65 channel=12
    -1, -5, -2, -1, 6, 6, -9, 3, -1,
    -- filter=65 channel=13
    -8, 1, 5, -8, -6, -2, 7, 10, 5,
    -- filter=65 channel=14
    0, 6, 3, 4, 3, -7, 4, 3, 6,
    -- filter=65 channel=15
    6, -10, 6, 7, 4, 9, 0, 2, 7,
    -- filter=65 channel=16
    6, 8, -4, 0, -4, 3, -9, -7, 8,
    -- filter=65 channel=17
    -8, 8, -4, 5, -10, 0, 6, -6, 4,
    -- filter=65 channel=18
    5, 5, -9, -3, 2, 5, 9, 2, -8,
    -- filter=65 channel=19
    6, 8, 7, 6, 10, -5, 0, -4, 0,
    -- filter=65 channel=20
    -10, 5, -5, 5, 6, -10, 10, 3, -3,
    -- filter=65 channel=21
    1, 0, -10, 1, 0, -3, 1, 8, -2,
    -- filter=65 channel=22
    -7, 9, -10, 6, -9, -6, -4, 0, -3,
    -- filter=65 channel=23
    7, -7, -7, -2, -9, 4, -9, 9, -4,
    -- filter=65 channel=24
    3, 2, -4, 0, -4, -4, 1, -5, 0,
    -- filter=65 channel=25
    -1, -5, -3, -5, 2, 8, 3, 7, 6,
    -- filter=65 channel=26
    -3, 0, 1, -5, 0, -1, 1, 8, 4,
    -- filter=65 channel=27
    1, 2, -4, 0, 6, 3, -3, -9, -5,
    -- filter=65 channel=28
    -9, -3, 9, -3, -8, -8, -6, 0, 0,
    -- filter=65 channel=29
    -7, 6, 10, -7, 8, -9, -9, 3, 0,
    -- filter=65 channel=30
    -3, -1, -10, -4, 6, 8, -1, 2, 5,
    -- filter=65 channel=31
    -8, 5, -6, -10, 2, -7, 3, 7, 3,
    -- filter=65 channel=32
    -1, 1, 1, 4, 4, -9, 7, 7, -4,
    -- filter=65 channel=33
    -2, 8, -7, 6, 4, 5, -2, -2, 0,
    -- filter=65 channel=34
    -2, 5, -10, 7, 7, 3, -10, -10, -5,
    -- filter=65 channel=35
    -6, -5, 5, 0, -1, 4, -4, 6, 2,
    -- filter=65 channel=36
    2, -8, -8, 1, 0, -4, 9, 0, -7,
    -- filter=65 channel=37
    10, 2, 3, -9, -8, -8, 2, -3, 9,
    -- filter=65 channel=38
    10, -2, -9, -8, -5, 8, 2, -4, 4,
    -- filter=65 channel=39
    -10, -6, -4, 7, 3, -10, 5, -1, 9,
    -- filter=65 channel=40
    5, 0, -2, -2, 0, 3, -2, 0, 5,
    -- filter=65 channel=41
    -5, -2, -3, -9, -7, -6, 6, 0, 5,
    -- filter=65 channel=42
    8, -4, -1, -3, -8, 4, 0, 10, 1,
    -- filter=65 channel=43
    -8, -7, 1, -2, -5, 5, 0, 5, 1,
    -- filter=65 channel=44
    0, -7, -5, -3, -9, 0, 8, 3, 0,
    -- filter=65 channel=45
    6, -7, 3, 7, -5, 0, 0, 0, -5,
    -- filter=65 channel=46
    1, 3, 0, 7, -10, -3, -3, -5, -6,
    -- filter=65 channel=47
    8, -5, 6, -7, -7, 4, 0, 0, 9,
    -- filter=65 channel=48
    -9, 5, -2, 7, -1, -6, -1, -8, 7,
    -- filter=65 channel=49
    2, -9, 0, 0, 6, 6, 9, -9, 1,
    -- filter=65 channel=50
    2, 7, 8, 3, -1, 0, -7, 0, 1,
    -- filter=65 channel=51
    -7, 7, -3, 7, -6, 10, 5, -9, 9,
    -- filter=65 channel=52
    0, -7, -2, -1, 7, -5, 1, 3, -8,
    -- filter=65 channel=53
    0, -1, 9, -8, -2, -7, -9, -6, 10,
    -- filter=65 channel=54
    -7, -9, -10, -9, 3, 0, 5, -3, -4,
    -- filter=65 channel=55
    -9, 4, -2, -5, 8, 10, 7, 7, -4,
    -- filter=65 channel=56
    9, 0, 3, 3, -4, 5, -9, -2, -5,
    -- filter=65 channel=57
    3, 1, 0, -8, -3, 3, 9, -1, 5,
    -- filter=65 channel=58
    0, -9, 6, 6, -5, 8, -9, -10, -8,
    -- filter=65 channel=59
    -9, -8, 5, -7, -4, -2, 5, 2, -4,
    -- filter=65 channel=60
    7, -4, -9, -7, -9, -6, -4, 5, 6,
    -- filter=65 channel=61
    5, 3, 9, -6, 9, 4, 3, 0, -5,
    -- filter=65 channel=62
    7, -4, 0, -9, 5, -3, 1, -7, 0,
    -- filter=65 channel=63
    0, 7, 3, -2, -1, 9, 3, 0, -3,
    -- filter=66 channel=0
    15, 8, -16, 11, 13, -7, 0, 8, -12,
    -- filter=66 channel=1
    -12, 11, -2, -6, 17, -4, -12, 4, -11,
    -- filter=66 channel=2
    -7, 6, -15, -11, 13, -16, -8, 11, -7,
    -- filter=66 channel=3
    12, 6, -15, 5, 11, -2, 14, 0, -12,
    -- filter=66 channel=4
    0, 15, 4, -5, 8, 0, -3, 15, -14,
    -- filter=66 channel=5
    2, 10, 0, -10, 15, 3, 4, 6, 10,
    -- filter=66 channel=6
    -1, -4, -12, -1, 1, -15, -3, 2, -5,
    -- filter=66 channel=7
    13, 10, 4, 1, 6, 20, -4, 19, 2,
    -- filter=66 channel=8
    -8, 8, -22, -15, 31, -18, -5, 27, -11,
    -- filter=66 channel=9
    7, -5, -2, 8, -2, 2, 9, -7, 2,
    -- filter=66 channel=10
    -2, -4, -6, 6, -13, -5, 6, 1, -9,
    -- filter=66 channel=11
    -14, 16, 0, -4, 8, -1, -10, 16, -2,
    -- filter=66 channel=12
    7, 8, 7, 9, -5, 8, 7, 3, -4,
    -- filter=66 channel=13
    10, 6, -6, 2, 13, -5, 11, -2, -6,
    -- filter=66 channel=14
    5, 13, 6, 5, 16, 10, 14, 3, 12,
    -- filter=66 channel=15
    7, 7, -29, 5, 22, -34, -3, 18, -12,
    -- filter=66 channel=16
    -4, 19, -23, -1, 23, -18, 3, 23, -17,
    -- filter=66 channel=17
    -13, 18, -13, -11, 21, -17, -8, 26, 1,
    -- filter=66 channel=18
    11, 3, 4, 3, -3, -15, 14, 0, 1,
    -- filter=66 channel=19
    -11, 14, -3, -31, 2, 9, -22, 8, 10,
    -- filter=66 channel=20
    22, 14, 1, 11, -4, 15, 10, -3, 4,
    -- filter=66 channel=21
    5, 0, 6, -7, -10, -7, -11, -7, -4,
    -- filter=66 channel=22
    0, 3, -1, 6, -4, 7, 8, 8, 0,
    -- filter=66 channel=23
    -11, -3, 0, -3, 10, -2, 0, 1, 3,
    -- filter=66 channel=24
    -5, 18, 6, -13, 21, 0, -13, 22, -3,
    -- filter=66 channel=25
    1, 0, -12, -5, 6, -26, 8, 0, -6,
    -- filter=66 channel=26
    19, 18, 17, 32, 13, 5, 14, 18, 15,
    -- filter=66 channel=27
    -8, 8, -11, -12, 28, -24, -14, 23, -9,
    -- filter=66 channel=28
    -4, 15, -17, -23, 21, -16, -18, 12, -1,
    -- filter=66 channel=29
    12, 12, -19, 9, 7, -41, 9, 18, -25,
    -- filter=66 channel=30
    12, 52, 13, 5, 48, 39, 8, 49, 28,
    -- filter=66 channel=31
    7, 7, -6, 6, 2, -2, 2, -8, 0,
    -- filter=66 channel=32
    -12, 6, 3, 1, -4, 5, -10, 0, -7,
    -- filter=66 channel=33
    0, 6, 9, 0, -8, 0, 0, 8, 7,
    -- filter=66 channel=34
    3, 3, 13, 3, 8, -4, 0, 18, 12,
    -- filter=66 channel=35
    1, 16, -8, -7, 16, -14, 3, 6, -6,
    -- filter=66 channel=36
    -9, 4, 9, -9, 7, 9, 2, -7, 0,
    -- filter=66 channel=37
    -8, 6, -3, -3, 10, -2, -13, 0, 0,
    -- filter=66 channel=38
    -2, 8, -9, -2, 32, -14, -9, 15, -7,
    -- filter=66 channel=39
    -8, -4, -6, 4, -8, -5, 8, 7, 2,
    -- filter=66 channel=40
    -8, 7, -9, 5, 4, -7, 10, 12, 11,
    -- filter=66 channel=41
    -8, 29, -23, 10, 26, -27, 3, 11, -18,
    -- filter=66 channel=42
    -6, -7, 7, -7, -9, -4, 2, -1, -7,
    -- filter=66 channel=43
    -11, -6, 10, -8, 0, -8, 0, -1, -3,
    -- filter=66 channel=44
    -14, 4, 5, -7, 4, 3, -11, 9, 19,
    -- filter=66 channel=45
    8, -8, 6, 6, 5, 7, 10, -10, 0,
    -- filter=66 channel=46
    29, 19, 8, 28, 18, 19, 27, 12, 0,
    -- filter=66 channel=47
    0, 6, -6, -3, -4, 1, -10, -10, 6,
    -- filter=66 channel=48
    15, -2, -15, 17, -8, -16, 12, 13, 3,
    -- filter=66 channel=49
    10, 16, -18, 0, 0, -9, -3, -2, 3,
    -- filter=66 channel=50
    -4, 17, 21, -1, 18, 32, 9, 15, 6,
    -- filter=66 channel=51
    2, 4, -1, -6, -5, -7, -6, 10, 10,
    -- filter=66 channel=52
    -6, 7, 10, 0, -9, 5, 1, -7, -6,
    -- filter=66 channel=53
    14, 23, 8, 10, 31, 26, 8, 28, 32,
    -- filter=66 channel=54
    -11, 9, 4, -6, 16, -9, -14, 11, 2,
    -- filter=66 channel=55
    -3, 4, 10, 4, -10, -5, -8, -10, 6,
    -- filter=66 channel=56
    0, 5, 17, 11, 0, 9, 0, 8, 3,
    -- filter=66 channel=57
    -5, 2, 1, 6, 0, -4, -6, -1, -5,
    -- filter=66 channel=58
    -2, 1, -6, 10, -8, 1, 3, 4, 9,
    -- filter=66 channel=59
    15, 0, -16, 19, 7, -16, -3, 7, -4,
    -- filter=66 channel=60
    -1, 27, -14, 1, 36, -38, 2, 22, -30,
    -- filter=66 channel=61
    -17, 23, -3, -11, 35, -15, -20, 23, -2,
    -- filter=66 channel=62
    -14, 4, -10, -1, 23, -15, -7, 11, -14,
    -- filter=66 channel=63
    -9, -2, -7, -5, -9, -10, -1, -7, -3,
    -- filter=67 channel=0
    -4, 0, -1, -8, -4, -3, -2, -5, 8,
    -- filter=67 channel=1
    3, 1, -3, 8, 3, -10, 11, -3, -2,
    -- filter=67 channel=2
    -3, 3, -6, -3, -5, -7, 7, -1, -4,
    -- filter=67 channel=3
    -9, 0, -9, 7, -8, 0, -1, -10, -2,
    -- filter=67 channel=4
    -3, 2, -2, -4, -5, -7, -3, -4, 6,
    -- filter=67 channel=5
    -2, 9, -7, 6, -3, -9, -8, -2, -9,
    -- filter=67 channel=6
    -5, -4, -6, -7, 4, 0, 1, 7, 4,
    -- filter=67 channel=7
    -3, 8, -3, 0, -7, -1, -8, 1, -7,
    -- filter=67 channel=8
    15, -5, -4, 6, -13, 9, 11, -11, -3,
    -- filter=67 channel=9
    -4, -1, 10, 14, 7, -5, 0, 10, 7,
    -- filter=67 channel=10
    0, -2, 3, 8, 2, 6, -6, -8, 4,
    -- filter=67 channel=11
    1, -7, -1, 0, 2, -1, 6, -4, 4,
    -- filter=67 channel=12
    1, -7, 4, 8, 0, -4, 3, 0, 3,
    -- filter=67 channel=13
    1, 8, 0, 5, -8, 1, -9, -1, -3,
    -- filter=67 channel=14
    4, 2, -7, 10, 9, -7, -1, -4, -6,
    -- filter=67 channel=15
    -5, -4, 5, 10, 0, 9, -5, -5, 10,
    -- filter=67 channel=16
    6, 7, 5, 2, 0, -1, 1, -6, -1,
    -- filter=67 channel=17
    2, -4, 0, 11, -1, 1, -3, -11, 10,
    -- filter=67 channel=18
    2, -1, 13, 2, -6, 0, -3, -6, 14,
    -- filter=67 channel=19
    -1, 0, -5, 10, 9, 4, -6, 5, -9,
    -- filter=67 channel=20
    8, 0, -7, 11, 1, 10, 12, 1, 14,
    -- filter=67 channel=21
    -6, 1, 3, 8, 5, 0, 8, 1, 1,
    -- filter=67 channel=22
    -5, 7, 0, 5, -6, 5, 7, 7, -5,
    -- filter=67 channel=23
    9, 7, -5, -6, 2, 4, -2, 7, 6,
    -- filter=67 channel=24
    6, 10, 8, 2, 2, 8, -4, -2, 9,
    -- filter=67 channel=25
    1, -10, -9, -2, 4, -7, 10, 6, 10,
    -- filter=67 channel=26
    -9, -2, -7, -9, 3, 0, 3, 0, 6,
    -- filter=67 channel=27
    -8, -4, -7, -5, -11, -1, -9, 0, 7,
    -- filter=67 channel=28
    0, 5, 0, -6, 0, 2, 11, -1, 1,
    -- filter=67 channel=29
    -2, 1, -9, -5, -6, -11, -8, -2, -3,
    -- filter=67 channel=30
    1, -3, -9, 0, -2, -4, 10, 0, -8,
    -- filter=67 channel=31
    2, 4, 4, 8, 0, -8, 2, 0, -3,
    -- filter=67 channel=32
    5, -8, 0, -8, -1, 0, 2, 5, -8,
    -- filter=67 channel=33
    0, 0, -8, -1, 8, -5, 4, 10, -2,
    -- filter=67 channel=34
    7, -7, -9, -5, 5, -3, -4, -5, -9,
    -- filter=67 channel=35
    8, 5, 4, -6, -5, -3, -6, -3, -1,
    -- filter=67 channel=36
    -5, -8, 2, -10, 6, -9, -3, -9, -1,
    -- filter=67 channel=37
    8, 8, -3, 7, 3, -1, 1, -11, -2,
    -- filter=67 channel=38
    12, -8, -2, -1, -4, -1, 5, 4, 6,
    -- filter=67 channel=39
    -3, 7, 2, 10, -6, 1, -1, 0, 0,
    -- filter=67 channel=40
    6, 9, -1, 7, -7, -8, -2, -3, -6,
    -- filter=67 channel=41
    0, -1, 4, -6, -14, 6, 0, -8, -1,
    -- filter=67 channel=42
    -7, 8, 10, 0, -10, -9, 0, 8, 6,
    -- filter=67 channel=43
    11, 2, -4, 2, -1, -1, 6, 3, -11,
    -- filter=67 channel=44
    -3, 0, 6, -4, -5, 1, 0, -9, 3,
    -- filter=67 channel=45
    3, 1, 10, 6, 3, 0, -8, -3, 0,
    -- filter=67 channel=46
    10, 4, -1, -5, -4, -8, 1, -4, 9,
    -- filter=67 channel=47
    -6, -4, -6, 3, -1, 1, 6, 4, 9,
    -- filter=67 channel=48
    -2, -8, 8, 4, -10, 5, -6, 9, -3,
    -- filter=67 channel=49
    7, 0, 12, 5, 6, 2, 3, 7, 0,
    -- filter=67 channel=50
    3, 9, -8, 13, 10, -7, -7, 2, 7,
    -- filter=67 channel=51
    -5, -3, 1, -1, -8, 8, -6, -8, -2,
    -- filter=67 channel=52
    -1, -2, -3, -9, 10, 4, -3, -4, 5,
    -- filter=67 channel=53
    -1, -6, 1, 10, -4, -4, 0, 0, 5,
    -- filter=67 channel=54
    8, 0, 4, -8, 5, 0, -3, -3, 4,
    -- filter=67 channel=55
    -7, -9, -9, -4, 3, 9, -2, -3, 0,
    -- filter=67 channel=56
    0, 9, -3, 5, -6, 5, 9, 10, -10,
    -- filter=67 channel=57
    -2, 2, 4, 7, 1, 8, -10, -5, -4,
    -- filter=67 channel=58
    7, 9, 10, 10, -1, 9, 7, 1, 7,
    -- filter=67 channel=59
    1, 0, -11, 2, -5, 8, 6, 5, 11,
    -- filter=67 channel=60
    -4, -1, 8, 8, -11, -9, 0, 5, 11,
    -- filter=67 channel=61
    3, -4, 7, 1, -6, 1, 1, -12, -9,
    -- filter=67 channel=62
    0, -4, 3, 3, 4, 5, -3, 5, -5,
    -- filter=67 channel=63
    10, 7, -2, -4, 2, -7, 8, -5, 2,
    -- filter=68 channel=0
    7, 0, -9, 6, 7, 6, 2, -5, -10,
    -- filter=68 channel=1
    8, 3, 0, 7, -3, 8, -1, -1, 4,
    -- filter=68 channel=2
    0, -3, 3, 5, 0, 6, 1, 5, -6,
    -- filter=68 channel=3
    5, -2, 2, -10, 4, 0, 7, -3, -9,
    -- filter=68 channel=4
    -8, 0, 4, -7, 10, -1, 12, 11, 11,
    -- filter=68 channel=5
    -5, -6, 6, 0, 8, -9, 2, -4, -9,
    -- filter=68 channel=6
    -9, -7, 7, 1, -1, 8, 12, 4, -8,
    -- filter=68 channel=7
    -4, 6, 2, 5, 5, -7, 4, 0, -1,
    -- filter=68 channel=8
    4, 2, -13, 0, -1, -1, 5, 11, 8,
    -- filter=68 channel=9
    -5, -1, -3, -8, 0, 6, 6, 12, 8,
    -- filter=68 channel=10
    5, -8, 9, 2, 6, 8, -7, 1, 7,
    -- filter=68 channel=11
    2, -4, 6, 0, 7, -7, 0, 0, 12,
    -- filter=68 channel=12
    9, -7, -4, -5, 9, 8, 6, 7, -6,
    -- filter=68 channel=13
    2, 7, 3, 2, 7, -2, 5, 1, 7,
    -- filter=68 channel=14
    -10, -8, -2, 7, -8, 8, -9, -4, -6,
    -- filter=68 channel=15
    -5, -11, 4, 10, 5, -7, 0, 0, 2,
    -- filter=68 channel=16
    -15, -7, -4, 0, 3, 3, 15, 16, -3,
    -- filter=68 channel=17
    -7, -7, -3, 0, 3, -1, 16, -4, 1,
    -- filter=68 channel=18
    1, 15, -2, 7, 4, 14, 4, -3, 0,
    -- filter=68 channel=19
    9, 3, 1, 11, 11, -5, -1, -2, 10,
    -- filter=68 channel=20
    -9, 8, 8, 0, -3, -1, 2, -5, -10,
    -- filter=68 channel=21
    3, 6, 9, -8, 11, -8, 2, 9, 11,
    -- filter=68 channel=22
    -9, 10, 3, -1, 9, 3, -2, 9, -10,
    -- filter=68 channel=23
    -9, 0, -6, 4, 0, 9, 3, 1, 3,
    -- filter=68 channel=24
    3, -10, -1, 9, 1, 7, 13, -2, -4,
    -- filter=68 channel=25
    -8, -12, -18, 2, -11, -3, 4, 0, -7,
    -- filter=68 channel=26
    -6, -5, -7, -9, 2, -4, -3, 4, -3,
    -- filter=68 channel=27
    -15, -10, -19, 12, 5, -13, 10, 11, 2,
    -- filter=68 channel=28
    5, 1, -3, 4, 9, 5, 13, 2, 8,
    -- filter=68 channel=29
    -5, -15, -14, -2, 10, 0, 7, 14, 1,
    -- filter=68 channel=30
    0, -8, -11, 4, 4, 2, -5, -5, -9,
    -- filter=68 channel=31
    -9, 3, -8, -1, 7, -1, -10, 5, 9,
    -- filter=68 channel=32
    -4, -2, -12, 4, 4, -9, -1, 0, 0,
    -- filter=68 channel=33
    8, 7, 3, 0, 2, 3, 3, 0, -5,
    -- filter=68 channel=34
    5, -4, -6, -3, 2, 4, 9, -4, 5,
    -- filter=68 channel=35
    4, -12, 1, 8, 0, -8, -2, 0, -7,
    -- filter=68 channel=36
    3, 0, -1, -6, 7, -10, 8, 2, 1,
    -- filter=68 channel=37
    -6, -6, -10, 2, 6, -9, 2, 11, 1,
    -- filter=68 channel=38
    -13, 0, -17, -8, 0, -4, 5, 7, -6,
    -- filter=68 channel=39
    -5, 1, 0, -5, -8, 2, 6, -8, -4,
    -- filter=68 channel=40
    -7, 8, 4, 10, 1, 6, -1, -6, -5,
    -- filter=68 channel=41
    -14, -12, -2, 1, 5, 4, 18, 12, -9,
    -- filter=68 channel=42
    -3, 7, 7, 5, 6, 0, -9, 1, 0,
    -- filter=68 channel=43
    15, 4, 10, 8, -6, 2, 13, -1, 0,
    -- filter=68 channel=44
    0, -7, -3, -4, 0, -4, -5, -4, -7,
    -- filter=68 channel=45
    0, -2, -1, -2, -5, 3, -8, -5, -2,
    -- filter=68 channel=46
    0, 6, -4, 4, 3, -7, 3, 5, 4,
    -- filter=68 channel=47
    6, -8, -1, -10, -1, 9, 9, 9, -3,
    -- filter=68 channel=48
    0, 9, -12, 0, -7, 3, -6, -7, 0,
    -- filter=68 channel=49
    6, 2, -7, 6, 12, 5, 5, -6, 4,
    -- filter=68 channel=50
    -1, -10, 4, -7, -11, 8, 0, -3, 3,
    -- filter=68 channel=51
    -5, -6, 12, -1, -9, -7, 2, 4, 0,
    -- filter=68 channel=52
    8, -7, -5, 1, 5, -1, -1, -8, 10,
    -- filter=68 channel=53
    -6, 4, -9, 0, -12, -8, -10, -11, 4,
    -- filter=68 channel=54
    5, 0, 5, -1, 9, -3, 4, 7, 3,
    -- filter=68 channel=55
    -5, 0, -9, -9, -5, 0, -5, -7, -8,
    -- filter=68 channel=56
    3, 5, 5, 5, -10, -1, 1, -3, 8,
    -- filter=68 channel=57
    -9, 2, -5, 8, 1, -7, 2, -10, 2,
    -- filter=68 channel=58
    3, 1, 12, 0, 10, 8, 1, -8, 3,
    -- filter=68 channel=59
    -14, -14, -5, -8, -7, -14, -1, 7, 2,
    -- filter=68 channel=60
    -16, -1, -16, -1, -1, -1, 14, 3, -2,
    -- filter=68 channel=61
    2, -7, -12, -7, -7, -11, 10, 14, 10,
    -- filter=68 channel=62
    2, 2, -6, 9, 5, -9, 7, -8, 5,
    -- filter=68 channel=63
    6, 0, -8, 2, -4, -3, -10, 9, 0,
    -- filter=69 channel=0
    -1, 10, -10, -2, -3, -5, 11, -2, 3,
    -- filter=69 channel=1
    7, 1, 7, 4, 10, 5, 5, -9, 8,
    -- filter=69 channel=2
    -5, 6, -7, 0, 7, -14, 6, 0, 3,
    -- filter=69 channel=3
    6, 4, 1, 1, 10, -8, -9, 1, -6,
    -- filter=69 channel=4
    -5, -5, 5, -6, -1, -4, 3, 0, 5,
    -- filter=69 channel=5
    -4, -6, -4, -1, -10, -2, -3, -1, 6,
    -- filter=69 channel=6
    -5, 0, -6, 0, -3, -4, 0, 1, -8,
    -- filter=69 channel=7
    0, 3, 9, -3, -2, 3, 0, -7, -3,
    -- filter=69 channel=8
    0, -2, -13, 6, -4, 1, 10, -8, 2,
    -- filter=69 channel=9
    5, 11, 2, 2, 0, -6, 4, 8, 12,
    -- filter=69 channel=10
    -7, 1, 11, 7, 3, 3, 9, 0, -6,
    -- filter=69 channel=11
    -5, 10, 9, 8, 0, 8, -5, 11, -8,
    -- filter=69 channel=12
    -8, -4, 10, -1, -7, 5, -2, -6, 4,
    -- filter=69 channel=13
    -2, 0, -9, 6, 4, -3, -6, -4, -3,
    -- filter=69 channel=14
    -8, -7, -6, 5, -1, 8, -7, 4, -5,
    -- filter=69 channel=15
    -2, -4, -5, -8, -2, -12, -4, -2, 0,
    -- filter=69 channel=16
    -8, -4, -13, 9, 4, -5, 6, 6, -5,
    -- filter=69 channel=17
    8, 5, -1, -5, 7, -6, -2, 1, -9,
    -- filter=69 channel=18
    4, -7, -2, -6, 7, 6, -2, -4, 7,
    -- filter=69 channel=19
    -9, 2, 8, -9, -5, -7, -12, 0, 0,
    -- filter=69 channel=20
    -1, -2, -1, 1, -2, 4, 5, -7, -4,
    -- filter=69 channel=21
    7, 3, 7, 9, -10, 9, 9, -3, 9,
    -- filter=69 channel=22
    -1, -8, -4, 7, 7, 4, 0, 5, 9,
    -- filter=69 channel=23
    1, 7, 10, 6, 8, 5, 4, 0, 9,
    -- filter=69 channel=24
    6, -2, -4, -5, 6, 9, 7, 11, -6,
    -- filter=69 channel=25
    -7, 10, 0, -7, -9, -11, -6, 5, -6,
    -- filter=69 channel=26
    -1, -3, -4, 4, -3, 4, -6, -10, -8,
    -- filter=69 channel=27
    -5, 3, -9, 9, 3, -7, 0, 12, -13,
    -- filter=69 channel=28
    2, 7, -8, 4, 8, 7, -8, -9, -8,
    -- filter=69 channel=29
    1, -4, -17, 6, 3, -11, 0, -3, -13,
    -- filter=69 channel=30
    -5, 2, 16, -5, -4, 0, -1, 12, 11,
    -- filter=69 channel=31
    0, -7, -2, 0, -8, 9, 3, -4, 9,
    -- filter=69 channel=32
    8, -3, -6, 8, -3, 2, 8, 2, 1,
    -- filter=69 channel=33
    0, -2, 3, -1, -1, 2, -5, -9, -4,
    -- filter=69 channel=34
    -2, -4, -9, 6, 5, 9, 2, -2, 5,
    -- filter=69 channel=35
    14, 8, 0, 6, 16, 0, 4, 8, 0,
    -- filter=69 channel=36
    0, 6, 0, -10, 2, 4, 3, 8, -2,
    -- filter=69 channel=37
    -10, 6, -2, -2, -5, 5, -7, 8, -8,
    -- filter=69 channel=38
    -7, 9, 4, 5, 9, -9, -5, -1, 5,
    -- filter=69 channel=39
    -9, -2, 9, -9, 7, 8, -9, -3, -7,
    -- filter=69 channel=40
    2, -5, 0, -6, 1, 10, -4, 0, -9,
    -- filter=69 channel=41
    6, 6, -12, -6, 4, -16, 8, 0, -15,
    -- filter=69 channel=42
    -2, -7, 0, 7, -4, -3, -4, -7, 0,
    -- filter=69 channel=43
    -8, 5, 0, 0, 4, -8, -10, -7, -10,
    -- filter=69 channel=44
    10, -2, 3, 0, -6, 8, 6, 2, 3,
    -- filter=69 channel=45
    3, -10, -5, 9, -4, 9, 8, 4, -4,
    -- filter=69 channel=46
    -9, -10, 5, 9, -9, -5, 10, 9, -6,
    -- filter=69 channel=47
    -5, -5, -6, -9, 10, -8, 2, 6, 2,
    -- filter=69 channel=48
    5, -1, 2, -10, 1, -1, -9, -8, -10,
    -- filter=69 channel=49
    1, 11, -9, 10, 3, 0, 0, 8, -6,
    -- filter=69 channel=50
    -1, 0, 7, -7, 0, 0, 5, -3, -3,
    -- filter=69 channel=51
    -3, -2, 0, -3, 6, 0, -6, 1, 2,
    -- filter=69 channel=52
    7, 0, 0, 5, 7, 10, 0, -7, -7,
    -- filter=69 channel=53
    -6, 12, 15, -1, 13, 0, 3, 5, 10,
    -- filter=69 channel=54
    -4, 11, 0, -6, 6, -1, -8, 11, -4,
    -- filter=69 channel=55
    -9, -3, -1, 4, -8, 10, 3, 3, 9,
    -- filter=69 channel=56
    5, -4, 1, -2, -1, 6, -6, -7, 0,
    -- filter=69 channel=57
    4, -1, 7, 9, -6, -10, 9, 0, 7,
    -- filter=69 channel=58
    5, 0, 6, -4, 2, 3, -9, 9, 5,
    -- filter=69 channel=59
    11, 2, -12, -8, -6, 0, 3, 4, 4,
    -- filter=69 channel=60
    13, 7, -8, 13, 5, -2, -2, 3, -14,
    -- filter=69 channel=61
    9, 3, 6, 1, 13, 3, -2, 12, -3,
    -- filter=69 channel=62
    -2, -2, 0, -1, 0, 4, -2, 2, 2,
    -- filter=69 channel=63
    -8, 6, 9, 9, 0, -7, 8, -3, 3,
    -- filter=70 channel=0
    -10, 0, -13, -9, 4, -6, -14, -7, 11,
    -- filter=70 channel=1
    2, -6, 1, 9, -2, 21, 4, 0, 1,
    -- filter=70 channel=2
    6, 6, 12, 10, 11, 23, -2, 8, 16,
    -- filter=70 channel=3
    5, 6, 1, -4, 8, 17, -12, -2, 10,
    -- filter=70 channel=4
    -9, 7, 4, 0, 2, 5, -7, 1, 3,
    -- filter=70 channel=5
    5, 0, 17, 11, 1, 14, 4, 9, 4,
    -- filter=70 channel=6
    0, 12, 2, 0, 8, 5, 4, 4, 1,
    -- filter=70 channel=7
    -6, 0, 12, 2, 3, 10, 2, 6, -1,
    -- filter=70 channel=8
    2, -4, 17, -10, -6, 15, -20, 0, 16,
    -- filter=70 channel=9
    -5, -9, -7, -11, 3, 0, -19, -15, -15,
    -- filter=70 channel=10
    1, -7, -7, -10, 2, 0, 5, -7, 6,
    -- filter=70 channel=11
    -12, -12, 5, -12, 1, 14, -8, -6, 0,
    -- filter=70 channel=12
    8, -6, -1, 7, 0, 5, 0, -7, 7,
    -- filter=70 channel=13
    0, 6, 3, 10, 11, 17, 4, 4, 11,
    -- filter=70 channel=14
    0, 3, 4, -8, 10, 1, -2, -5, 0,
    -- filter=70 channel=15
    10, -3, 4, -7, 15, 6, -10, 6, 19,
    -- filter=70 channel=16
    10, 15, 30, -5, 22, 20, -3, 14, 23,
    -- filter=70 channel=17
    2, -8, 12, -12, -9, 9, -12, -3, -2,
    -- filter=70 channel=18
    -5, 0, -9, 10, 12, 7, -3, 2, 3,
    -- filter=70 channel=19
    9, 0, 6, 13, 6, 19, 9, 8, 16,
    -- filter=70 channel=20
    3, 1, 8, -3, 2, 13, 3, -3, 8,
    -- filter=70 channel=21
    3, -7, 1, 5, 6, -3, -1, 6, -11,
    -- filter=70 channel=22
    9, 9, 10, 5, 9, 5, 8, -2, 1,
    -- filter=70 channel=23
    -12, -14, -14, -10, -1, -13, -7, -14, 7,
    -- filter=70 channel=24
    6, -3, 11, 0, -10, -5, 0, 2, -2,
    -- filter=70 channel=25
    11, 16, 19, 0, 7, 8, -4, -2, 16,
    -- filter=70 channel=26
    3, 12, 14, 5, 14, 7, 0, 5, 16,
    -- filter=70 channel=27
    -10, -2, 13, -11, -9, 4, 0, -5, 14,
    -- filter=70 channel=28
    5, 6, 3, 9, 4, 23, -5, -5, 21,
    -- filter=70 channel=29
    -3, 7, 20, 11, 15, 32, -3, 0, 19,
    -- filter=70 channel=30
    7, 0, 4, 15, 15, 10, 2, 2, 13,
    -- filter=70 channel=31
    7, 2, -13, -8, -8, 0, -4, -13, -13,
    -- filter=70 channel=32
    -4, -2, -2, -12, -3, -1, 0, -2, -1,
    -- filter=70 channel=33
    8, 8, -6, 5, 4, 3, -10, 1, 0,
    -- filter=70 channel=34
    -2, -3, 0, 5, 0, 10, -4, -6, 7,
    -- filter=70 channel=35
    -15, -15, -11, 0, -18, 3, -9, -1, 0,
    -- filter=70 channel=36
    0, 6, -5, -12, -11, -9, -11, -10, -1,
    -- filter=70 channel=37
    6, 3, -3, 1, -6, 8, -12, -4, 7,
    -- filter=70 channel=38
    -9, 5, 14, -14, 0, 17, -10, -4, 16,
    -- filter=70 channel=39
    -7, 0, -8, -2, -1, 9, 9, 10, 1,
    -- filter=70 channel=40
    -6, -5, 7, 9, -6, 5, 5, 9, -10,
    -- filter=70 channel=41
    6, 6, 0, 1, -6, 7, -14, 5, 16,
    -- filter=70 channel=42
    -8, 0, -6, 7, 7, 3, 7, 0, -3,
    -- filter=70 channel=43
    27, 23, 19, 30, 19, 22, 34, 19, 12,
    -- filter=70 channel=44
    5, -7, 10, -10, -3, 11, 6, 3, -4,
    -- filter=70 channel=45
    -10, -5, 0, -9, -3, 5, 0, -4, 9,
    -- filter=70 channel=46
    13, 15, 6, 0, -1, 7, 0, 1, 5,
    -- filter=70 channel=47
    2, 8, -3, 1, 5, -5, 10, 0, 3,
    -- filter=70 channel=48
    2, 8, 14, 0, 10, 17, -5, 18, 13,
    -- filter=70 channel=49
    -5, -9, 4, 3, -5, -8, 3, 1, 3,
    -- filter=70 channel=50
    18, 11, 6, 0, 18, 0, -1, 17, -1,
    -- filter=70 channel=51
    -10, 0, -18, 1, -1, -17, 2, 0, -8,
    -- filter=70 channel=52
    8, 0, -3, -3, 8, 8, 2, 3, 6,
    -- filter=70 channel=53
    1, -7, -4, 0, 6, 0, 3, -3, 10,
    -- filter=70 channel=54
    -22, -15, -16, -22, -5, -9, -25, -18, -7,
    -- filter=70 channel=55
    4, 7, 3, 8, -9, -1, 0, -8, -3,
    -- filter=70 channel=56
    2, -1, 8, -3, -5, 8, 8, -2, 13,
    -- filter=70 channel=57
    5, -4, -5, -1, -9, -8, 10, -2, 8,
    -- filter=70 channel=58
    10, 7, 9, 10, 10, 11, -2, -2, 0,
    -- filter=70 channel=59
    3, 11, 4, 2, 10, 19, -12, -1, 11,
    -- filter=70 channel=60
    -7, -12, 14, -5, -1, 11, -22, -5, 14,
    -- filter=70 channel=61
    0, -20, 2, -2, -12, 9, -13, -21, 1,
    -- filter=70 channel=62
    -12, -1, -4, -10, 5, 8, -1, -5, 5,
    -- filter=70 channel=63
    -9, -4, -3, 0, 10, -5, 3, -2, 4,
    -- filter=71 channel=0
    10, -4, 8, -5, -7, 2, -5, -9, 3,
    -- filter=71 channel=1
    17, 11, 15, 4, 8, -5, 5, -9, -10,
    -- filter=71 channel=2
    14, 4, 13, -13, -8, -8, 1, -1, 4,
    -- filter=71 channel=3
    -3, 5, 4, 5, 1, -3, -3, 4, -5,
    -- filter=71 channel=4
    0, 15, 3, -9, 8, 3, -3, -2, 4,
    -- filter=71 channel=5
    -8, 7, 10, -2, -2, -6, -8, -3, -8,
    -- filter=71 channel=6
    1, 5, 9, 4, -1, 8, -2, 11, -10,
    -- filter=71 channel=7
    -5, -1, 0, -1, 6, -9, -4, -1, -8,
    -- filter=71 channel=8
    21, 19, 10, -7, 1, -12, -10, 0, -7,
    -- filter=71 channel=9
    -5, -8, -12, 10, -11, -9, -3, 3, -1,
    -- filter=71 channel=10
    2, 3, -4, 13, -1, 15, 10, 10, 0,
    -- filter=71 channel=11
    16, 9, 11, 6, -3, 5, -9, -13, -7,
    -- filter=71 channel=12
    11, -7, 8, 0, 0, -8, -1, 4, -8,
    -- filter=71 channel=13
    13, 8, -3, 16, 15, 5, -11, -4, -3,
    -- filter=71 channel=14
    7, -6, 7, -7, 9, 2, -1, -2, -8,
    -- filter=71 channel=15
    15, 8, 7, 0, 0, -13, -1, -10, -7,
    -- filter=71 channel=16
    15, 18, 7, -8, -4, 5, -1, -17, -15,
    -- filter=71 channel=17
    13, 17, 0, 1, -1, 3, 3, -4, -11,
    -- filter=71 channel=18
    5, -1, -2, 13, -5, 7, 13, 12, 13,
    -- filter=71 channel=19
    7, 6, 1, 0, 1, -4, -6, -2, -5,
    -- filter=71 channel=20
    -3, -6, -5, -6, 11, -2, 0, 7, 7,
    -- filter=71 channel=21
    -1, -2, 5, -2, -3, 8, 7, 11, 0,
    -- filter=71 channel=22
    1, -8, 7, 11, 1, 7, 2, -7, 1,
    -- filter=71 channel=23
    3, -6, 9, 0, 7, 8, 6, 9, -8,
    -- filter=71 channel=24
    1, 7, 12, 4, -4, -1, 0, -4, -2,
    -- filter=71 channel=25
    3, 5, -2, 0, -8, -10, -14, -4, -7,
    -- filter=71 channel=26
    -11, -2, 8, 4, -3, -9, -11, 3, 4,
    -- filter=71 channel=27
    2, 10, 15, 3, -8, -5, -8, -18, -19,
    -- filter=71 channel=28
    21, 7, 21, 5, -9, 3, 11, 3, -6,
    -- filter=71 channel=29
    13, 28, 16, -6, -10, 6, -7, -17, -4,
    -- filter=71 channel=30
    -2, -4, 4, 0, -7, -5, -12, 3, -3,
    -- filter=71 channel=31
    1, -6, -6, -1, 9, 0, 7, -8, -4,
    -- filter=71 channel=32
    -4, 2, -2, 9, 0, 2, -12, -13, 5,
    -- filter=71 channel=33
    8, 7, -8, 6, 0, -5, 0, -1, 4,
    -- filter=71 channel=34
    1, 0, -9, -2, -8, -7, 4, 3, 0,
    -- filter=71 channel=35
    10, -2, 0, -5, -6, -9, -1, -11, 0,
    -- filter=71 channel=36
    -7, 5, -8, -8, 11, 7, 0, 0, -4,
    -- filter=71 channel=37
    -3, 7, 9, 4, -8, 5, -3, -15, -9,
    -- filter=71 channel=38
    6, 8, 16, -9, 5, -2, -5, -7, -17,
    -- filter=71 channel=39
    4, -3, 8, 2, 3, 0, 1, -1, 4,
    -- filter=71 channel=40
    -3, -3, 7, 3, 5, -4, 8, -11, -2,
    -- filter=71 channel=41
    6, 5, 12, -8, -4, -12, -16, -6, -2,
    -- filter=71 channel=42
    0, -3, 10, 0, -8, 10, -4, -1, 1,
    -- filter=71 channel=43
    20, 14, 4, 12, 13, 23, 0, -3, 6,
    -- filter=71 channel=44
    -10, 4, -5, -10, -4, 0, -6, -13, -3,
    -- filter=71 channel=45
    8, 3, -6, -6, 8, -6, -7, 0, 2,
    -- filter=71 channel=46
    5, -8, -2, 4, -5, -11, -7, 7, 3,
    -- filter=71 channel=47
    -7, -2, -4, -2, -9, 3, -3, 10, 0,
    -- filter=71 channel=48
    10, 15, 5, -4, -5, 7, -10, 4, 5,
    -- filter=71 channel=49
    -6, 11, -5, -4, -12, 2, -2, 9, 2,
    -- filter=71 channel=50
    -9, 2, 13, 0, 10, 3, -4, 6, -2,
    -- filter=71 channel=51
    0, -3, 0, 8, 10, 14, -3, 11, -1,
    -- filter=71 channel=52
    3, -2, -8, -4, 4, 0, 10, 3, -6,
    -- filter=71 channel=53
    -10, 6, -4, 0, -4, -7, -11, -14, -10,
    -- filter=71 channel=54
    9, 4, 0, -14, -11, 1, -14, -11, -12,
    -- filter=71 channel=55
    5, -9, -2, -9, -5, -7, -2, 4, -2,
    -- filter=71 channel=56
    8, 8, -1, 0, 8, 9, -6, -9, 6,
    -- filter=71 channel=57
    9, 10, 2, 7, -7, -6, -5, 4, 1,
    -- filter=71 channel=58
    -3, 0, 0, 11, 1, 3, 11, 5, 4,
    -- filter=71 channel=59
    15, 11, 2, -1, -13, 3, -13, -8, -11,
    -- filter=71 channel=60
    16, 19, 11, -2, 0, -2, -24, -7, -17,
    -- filter=71 channel=61
    16, 12, 8, 2, 1, 6, -17, -14, -10,
    -- filter=71 channel=62
    -2, 10, -1, 0, -5, -4, -8, 0, 4,
    -- filter=71 channel=63
    -10, -7, 5, 3, -3, 10, -8, 3, 5,
    -- filter=72 channel=0
    3, 6, 6, 8, 11, 0, -6, 15, 9,
    -- filter=72 channel=1
    -2, -22, -9, 0, -14, -10, -10, -3, -10,
    -- filter=72 channel=2
    9, -14, -8, -5, 0, -16, -6, -3, -16,
    -- filter=72 channel=3
    1, -5, -12, -2, -11, -7, 5, 3, -18,
    -- filter=72 channel=4
    7, 12, 8, 11, 8, 9, -1, 3, 13,
    -- filter=72 channel=5
    9, 0, 9, 0, 0, 1, 4, -3, 0,
    -- filter=72 channel=6
    6, -5, 5, 13, 12, 0, -7, 4, 3,
    -- filter=72 channel=7
    2, -3, -8, -12, -13, 6, 4, -11, -7,
    -- filter=72 channel=8
    6, 11, 14, 16, 12, 19, 10, 13, -2,
    -- filter=72 channel=9
    -13, -7, -18, -12, -15, -17, -12, -5, -15,
    -- filter=72 channel=10
    -10, -5, 0, -3, -6, 1, -4, -3, 2,
    -- filter=72 channel=11
    7, 1, 11, -3, 11, 3, 11, 10, -7,
    -- filter=72 channel=12
    1, 7, -8, 6, 0, 9, 9, 11, 6,
    -- filter=72 channel=13
    4, 20, 0, 7, 19, 4, 9, 14, 12,
    -- filter=72 channel=14
    3, -10, 2, -9, 0, 6, -9, -13, 5,
    -- filter=72 channel=15
    -1, 21, 5, 23, 13, 10, 0, 17, -6,
    -- filter=72 channel=16
    15, 11, -6, 9, 6, -6, 16, -4, -5,
    -- filter=72 channel=17
    -1, 8, 7, 17, 19, 10, 11, 9, 13,
    -- filter=72 channel=18
    20, 30, 18, 20, 29, 6, 17, 24, 22,
    -- filter=72 channel=19
    -4, -4, -10, 0, -19, -13, -6, -6, -17,
    -- filter=72 channel=20
    1, -18, -2, -8, -10, -3, -6, -9, -9,
    -- filter=72 channel=21
    -7, 6, 4, 10, 8, -8, 0, 3, -3,
    -- filter=72 channel=22
    -6, 5, -4, -9, -7, 0, 8, 5, -5,
    -- filter=72 channel=23
    4, 4, 8, 0, 2, 12, -3, 6, 4,
    -- filter=72 channel=24
    -3, 11, 0, 9, 11, 4, 6, 10, 16,
    -- filter=72 channel=25
    -15, -9, -27, -17, -23, -32, -10, -10, -32,
    -- filter=72 channel=26
    -2, -16, -7, -11, -9, -5, -2, -17, -10,
    -- filter=72 channel=27
    -9, 3, -11, -13, -9, -15, -6, -8, -9,
    -- filter=72 channel=28
    0, 12, 8, 7, 11, 1, 9, 6, 10,
    -- filter=72 channel=29
    0, 1, 1, 19, 19, -3, 0, 8, -4,
    -- filter=72 channel=30
    -25, -20, -10, -32, -16, -23, -21, -18, -1,
    -- filter=72 channel=31
    1, 5, -9, 2, -8, -10, -2, 0, -9,
    -- filter=72 channel=32
    -23, -18, -20, -20, -28, -9, -12, -11, -13,
    -- filter=72 channel=33
    -8, 4, 7, -3, -2, 6, 0, -2, 6,
    -- filter=72 channel=34
    1, -9, -14, -12, -1, 5, 0, 0, 4,
    -- filter=72 channel=35
    -1, -7, -14, -20, -13, -4, -22, -16, -9,
    -- filter=72 channel=36
    -1, 1, 11, -7, 2, 9, -1, 3, 2,
    -- filter=72 channel=37
    3, -13, 2, 6, -7, 0, -7, -3, -5,
    -- filter=72 channel=38
    8, -7, -12, 11, -4, -8, -9, 7, -7,
    -- filter=72 channel=39
    -5, 6, 6, -3, 8, -9, 5, 5, 5,
    -- filter=72 channel=40
    -2, -1, -10, -4, 0, -5, -7, -16, 3,
    -- filter=72 channel=41
    10, 12, -12, 15, 18, -4, -1, 5, -13,
    -- filter=72 channel=42
    -7, 0, -7, -6, 9, 5, 4, 7, -9,
    -- filter=72 channel=43
    -21, -25, -26, -30, -39, -36, -16, -27, -31,
    -- filter=72 channel=44
    -10, -25, 0, -7, -12, -10, -13, -17, -15,
    -- filter=72 channel=45
    8, -3, 1, -2, 6, -3, -9, -7, 8,
    -- filter=72 channel=46
    -12, -6, -9, 3, -14, -8, 4, -14, -5,
    -- filter=72 channel=47
    1, -8, 9, 7, 6, -9, 10, 9, 7,
    -- filter=72 channel=48
    2, 3, -9, -4, -5, 5, -8, 1, 4,
    -- filter=72 channel=49
    12, 20, 6, 11, 15, 2, -3, 2, 3,
    -- filter=72 channel=50
    -13, -25, -18, -6, -14, -13, 0, -3, -7,
    -- filter=72 channel=51
    9, 12, 3, 5, 16, 20, 9, 14, 6,
    -- filter=72 channel=52
    5, -7, 10, 8, -3, 5, 9, 1, -2,
    -- filter=72 channel=53
    -17, -26, -21, -15, -19, -21, -20, -25, -1,
    -- filter=72 channel=54
    5, 0, -13, 2, 1, -8, -10, -17, 0,
    -- filter=72 channel=55
    10, -7, 0, -2, 9, 10, -3, 7, -4,
    -- filter=72 channel=56
    -8, -14, -8, 1, -6, 9, 7, 8, 3,
    -- filter=72 channel=57
    -3, 6, -8, -6, 5, 0, -5, 5, -9,
    -- filter=72 channel=58
    4, -8, -9, 3, 7, 0, -3, 7, 6,
    -- filter=72 channel=59
    8, 6, -18, -3, -10, -13, -2, -19, -14,
    -- filter=72 channel=60
    16, 25, 10, 11, 33, 18, 6, 22, 0,
    -- filter=72 channel=61
    0, 1, 14, -2, 8, 4, 2, 9, 6,
    -- filter=72 channel=62
    0, 5, -1, 0, -9, -13, -2, -4, -8,
    -- filter=72 channel=63
    -7, 0, 8, 2, -3, 5, -3, 2, 6,
    -- filter=73 channel=0
    4, -4, 9, -6, -6, -9, -9, 1, 2,
    -- filter=73 channel=1
    2, -6, -7, -2, 0, 3, -8, -2, -5,
    -- filter=73 channel=2
    -5, -10, -3, -1, -2, -2, 0, -3, -7,
    -- filter=73 channel=3
    9, 4, 5, 14, 11, 21, 20, 18, 5,
    -- filter=73 channel=4
    0, -4, -10, 8, 10, -2, -5, -2, -9,
    -- filter=73 channel=5
    5, 8, 2, 17, 15, 0, 13, 9, 11,
    -- filter=73 channel=6
    -2, 8, -8, -10, -1, -5, 7, 0, 7,
    -- filter=73 channel=7
    0, 8, -1, 2, -3, -9, -8, 0, -1,
    -- filter=73 channel=8
    -22, -8, -1, -4, -2, 15, 5, 17, -2,
    -- filter=73 channel=9
    -4, 2, 7, 7, 27, 8, 1, 12, 7,
    -- filter=73 channel=10
    -3, 3, -6, -10, -3, -8, -8, -6, -11,
    -- filter=73 channel=11
    -16, -7, -1, 1, -8, 1, 0, 14, -5,
    -- filter=73 channel=12
    -3, 7, 9, -7, -6, 0, -9, 0, -1,
    -- filter=73 channel=13
    -9, -12, 3, -6, -7, 0, 15, 5, 0,
    -- filter=73 channel=14
    8, 9, 9, 9, 2, 5, 2, -1, -4,
    -- filter=73 channel=15
    -6, -8, 5, 8, 1, 3, 2, 6, 9,
    -- filter=73 channel=16
    -26, -14, -1, 5, 10, 1, 17, 14, 0,
    -- filter=73 channel=17
    -7, -15, 0, 0, -1, 6, 16, 1, 15,
    -- filter=73 channel=18
    1, 2, -3, -2, 13, -3, 1, -6, -2,
    -- filter=73 channel=19
    -6, -1, -1, 10, 12, 1, 0, 9, -6,
    -- filter=73 channel=20
    -5, -2, 6, -6, 0, -2, 8, 13, 4,
    -- filter=73 channel=21
    0, -3, 10, 9, 7, -3, -2, -2, 3,
    -- filter=73 channel=22
    4, 9, -8, -5, -4, 0, 8, -8, 2,
    -- filter=73 channel=23
    -4, 4, 8, -2, -6, -9, -9, -12, -2,
    -- filter=73 channel=24
    -2, -5, 6, -7, -2, 4, -6, 11, 11,
    -- filter=73 channel=25
    -18, -2, 0, -12, 4, 6, 9, 13, -5,
    -- filter=73 channel=26
    -9, 2, 3, 0, 11, -3, 5, 10, 0,
    -- filter=73 channel=27
    -10, -14, 0, -14, -11, -7, 1, 8, 5,
    -- filter=73 channel=28
    -12, -2, 1, 4, 5, 6, -2, 4, 11,
    -- filter=73 channel=29
    -14, 1, 0, 1, 18, 4, 14, 18, -4,
    -- filter=73 channel=30
    -3, -13, 4, -8, 8, 11, 9, -2, 0,
    -- filter=73 channel=31
    4, -5, -7, -7, -1, -7, 6, -8, 10,
    -- filter=73 channel=32
    3, 8, -2, 0, -5, -2, -3, 6, 4,
    -- filter=73 channel=33
    7, 3, 5, 1, -8, 10, -6, 9, -5,
    -- filter=73 channel=34
    2, 5, 2, 3, 0, -4, -3, 12, 7,
    -- filter=73 channel=35
    -18, 2, 3, -6, -15, 6, -4, -6, -4,
    -- filter=73 channel=36
    -2, 5, -7, 11, 0, 0, 8, -3, -9,
    -- filter=73 channel=37
    0, -1, 9, 0, 12, 11, 8, 0, 7,
    -- filter=73 channel=38
    -16, -14, -1, 0, 1, -8, -2, 7, 10,
    -- filter=73 channel=39
    -8, -10, 3, -1, 0, 0, -2, -8, 10,
    -- filter=73 channel=40
    7, 7, 0, 0, -2, 4, -4, -2, 6,
    -- filter=73 channel=41
    -3, -12, 2, 1, 4, 3, 17, 19, 7,
    -- filter=73 channel=42
    -4, 4, 6, -5, 4, -10, -10, -9, 7,
    -- filter=73 channel=43
    -8, -12, -2, 0, -4, 0, -2, -7, 6,
    -- filter=73 channel=44
    9, 4, 4, -1, 12, 9, -9, 10, -1,
    -- filter=73 channel=45
    -5, -4, -9, 4, -3, 7, -9, -2, 5,
    -- filter=73 channel=46
    -7, -4, 5, 1, 10, 1, 6, 7, 2,
    -- filter=73 channel=47
    -3, 5, -1, -1, -5, -6, -1, 0, 5,
    -- filter=73 channel=48
    -8, 6, -4, 5, 5, 0, 10, 14, 10,
    -- filter=73 channel=49
    -8, 3, 6, 2, -4, 9, 5, -1, 4,
    -- filter=73 channel=50
    -1, 0, -1, -10, -9, 8, -5, 8, -7,
    -- filter=73 channel=51
    8, 5, 1, -5, -16, 5, 1, 2, -4,
    -- filter=73 channel=52
    7, 2, 3, 8, -5, -4, -1, -4, -1,
    -- filter=73 channel=53
    10, -10, 7, -3, -3, 1, -11, 1, 3,
    -- filter=73 channel=54
    7, 0, 17, 5, 18, 12, 15, 17, 16,
    -- filter=73 channel=55
    5, 4, 5, 0, 8, -3, -7, -3, 3,
    -- filter=73 channel=56
    -10, -8, 5, -2, 10, 6, 0, 4, 0,
    -- filter=73 channel=57
    -8, 7, -3, 6, 4, -6, 6, 9, 0,
    -- filter=73 channel=58
    5, 14, 3, 1, -7, -2, 3, -4, 2,
    -- filter=73 channel=59
    -9, 0, 13, 9, 13, 12, 18, 15, -4,
    -- filter=73 channel=60
    -19, -12, -4, -2, -2, 11, 18, 5, 1,
    -- filter=73 channel=61
    -16, -18, 4, 0, -2, 8, 14, 12, 0,
    -- filter=73 channel=62
    7, -3, -1, 13, 2, 5, 12, 2, 11,
    -- filter=73 channel=63
    -9, 4, 4, -6, -3, 9, 2, -7, -3,
    -- filter=74 channel=0
    1, -2, 12, -9, 7, 11, -14, 7, 11,
    -- filter=74 channel=1
    -10, -13, -2, -7, -3, 7, -7, 1, 0,
    -- filter=74 channel=2
    -10, 5, 6, -9, -2, 15, -15, 5, 8,
    -- filter=74 channel=3
    -13, 0, -1, -3, 4, 11, -15, -5, 5,
    -- filter=74 channel=4
    -5, 0, 7, -2, 7, 18, -16, 5, 5,
    -- filter=74 channel=5
    -10, 6, -4, -3, -7, 8, -1, 7, 0,
    -- filter=74 channel=6
    4, 0, 7, 2, -3, 16, -16, 9, 8,
    -- filter=74 channel=7
    15, -4, 12, 1, 2, 5, 7, 0, 3,
    -- filter=74 channel=8
    -12, 9, 11, -11, -4, 27, -22, 9, 25,
    -- filter=74 channel=9
    -10, -13, -5, 3, -3, 0, 3, 0, -9,
    -- filter=74 channel=10
    7, 0, -3, -1, 0, 0, -1, 8, -3,
    -- filter=74 channel=11
    -12, -2, 11, -21, -3, 6, -10, 0, 8,
    -- filter=74 channel=12
    -6, -3, -5, 1, -6, 5, 7, 10, 0,
    -- filter=74 channel=13
    -9, 7, 11, -6, 2, 14, -3, 1, 1,
    -- filter=74 channel=14
    12, 0, 0, 2, 12, 13, -7, -1, 10,
    -- filter=74 channel=15
    -10, 5, 16, -20, 0, 17, -16, 14, 19,
    -- filter=74 channel=16
    -15, 4, 5, -21, 12, 21, -31, 7, 32,
    -- filter=74 channel=17
    -14, 6, 17, -9, 1, 4, -25, -8, 23,
    -- filter=74 channel=18
    1, 0, 0, -10, 1, 9, 10, 5, -2,
    -- filter=74 channel=19
    -10, 0, 1, -3, 0, 5, -1, -6, 8,
    -- filter=74 channel=20
    3, 8, 4, 0, 12, 6, 2, 9, 8,
    -- filter=74 channel=21
    -9, 5, 0, 0, 3, 6, 1, 9, 6,
    -- filter=74 channel=22
    0, 8, 3, -5, 9, 7, 0, -2, -3,
    -- filter=74 channel=23
    -4, 2, 6, -13, -11, 10, -8, -2, -4,
    -- filter=74 channel=24
    -15, -14, 13, -13, -14, 5, -13, 0, 1,
    -- filter=74 channel=25
    -1, -10, 13, -8, -3, 7, -13, -5, 4,
    -- filter=74 channel=26
    15, -1, 4, 5, 21, 18, 4, 3, 10,
    -- filter=74 channel=27
    -17, -4, 13, -20, 5, 25, -22, 8, 25,
    -- filter=74 channel=28
    -12, -13, -2, -3, 2, 13, -17, -2, 15,
    -- filter=74 channel=29
    -8, 7, 7, -14, 11, 28, -18, 16, 32,
    -- filter=74 channel=30
    18, 14, 13, 8, 13, 15, 21, 0, 26,
    -- filter=74 channel=31
    7, 1, -6, -8, 8, -3, 4, -7, 6,
    -- filter=74 channel=32
    4, -8, 11, -12, -11, -4, -3, -10, -4,
    -- filter=74 channel=33
    -10, -7, -6, 1, 0, -10, 9, 2, -1,
    -- filter=74 channel=34
    6, 13, -2, -1, -2, 2, 0, 4, 16,
    -- filter=74 channel=35
    -10, 6, 22, -5, 11, 5, -2, 7, 5,
    -- filter=74 channel=36
    11, 2, -10, 4, -9, 0, -4, -3, 8,
    -- filter=74 channel=37
    -6, -9, 6, -15, 7, 0, 1, 6, -7,
    -- filter=74 channel=38
    -21, -3, 8, -14, 5, 11, -17, 9, 30,
    -- filter=74 channel=39
    -5, 10, -3, 0, 10, 8, -10, -5, 5,
    -- filter=74 channel=40
    1, -5, -4, -11, 6, 4, -12, 1, 6,
    -- filter=74 channel=41
    -13, 8, 17, -18, 15, 25, -29, 19, 20,
    -- filter=74 channel=42
    9, 0, 2, 6, 3, 9, 0, -9, 8,
    -- filter=74 channel=43
    11, 2, -5, 8, -17, -12, -2, -12, 5,
    -- filter=74 channel=44
    -7, -11, 2, 6, 4, 7, 2, -4, 2,
    -- filter=74 channel=45
    2, -9, -5, -3, -8, -1, 9, -5, 9,
    -- filter=74 channel=46
    2, 9, 21, 11, 23, 8, 6, 10, 14,
    -- filter=74 channel=47
    -2, 6, 9, 5, 4, -3, -7, -5, -6,
    -- filter=74 channel=48
    -9, 0, 3, 5, 0, 12, -3, 12, 1,
    -- filter=74 channel=49
    -6, 5, 10, -15, 12, 11, -15, 0, 14,
    -- filter=74 channel=50
    11, 5, 6, 10, -5, 15, -1, 0, 11,
    -- filter=74 channel=51
    -4, -6, 3, -10, 10, -2, -10, -2, -7,
    -- filter=74 channel=52
    -8, 9, -7, -4, -1, 1, 9, 0, 1,
    -- filter=74 channel=53
    5, 0, 12, 16, -5, 18, 12, -11, 22,
    -- filter=74 channel=54
    -11, -14, 0, -13, -1, -8, -4, 0, 0,
    -- filter=74 channel=55
    -7, 2, 2, 8, 0, -8, -7, 0, 2,
    -- filter=74 channel=56
    4, 0, -3, 7, 0, 4, 9, 2, -2,
    -- filter=74 channel=57
    8, -3, 1, -4, 9, 8, 8, 4, -9,
    -- filter=74 channel=58
    10, -3, 3, -3, 8, -2, 1, 12, 5,
    -- filter=74 channel=59
    -9, -5, 12, -19, 3, 6, -20, 7, 24,
    -- filter=74 channel=60
    -23, -4, 27, -26, 12, 22, -24, 23, 26,
    -- filter=74 channel=61
    -5, 5, 19, -31, 0, 22, -32, 9, 17,
    -- filter=74 channel=62
    -20, -9, 13, -13, -9, 13, -18, 9, 14,
    -- filter=74 channel=63
    -9, 2, 7, 4, -9, -6, -10, 10, 2,
    -- filter=75 channel=0
    1, 9, 9, 13, 6, 0, -9, -4, 6,
    -- filter=75 channel=1
    16, 31, 16, 14, 39, 21, 22, 12, 12,
    -- filter=75 channel=2
    14, 38, 17, 18, 28, 19, 10, 3, 11,
    -- filter=75 channel=3
    23, 20, 12, 15, 2, -2, -6, 1, 7,
    -- filter=75 channel=4
    -2, -9, -11, -6, -12, -12, -2, -19, -17,
    -- filter=75 channel=5
    0, -5, -8, -16, -9, -11, 0, 5, -2,
    -- filter=75 channel=6
    6, 4, -4, 4, 8, 0, -9, 0, -1,
    -- filter=75 channel=7
    -3, -6, -6, -2, 4, 3, 5, 3, -8,
    -- filter=75 channel=8
    3, 17, -3, 4, -10, -8, -13, -16, -25,
    -- filter=75 channel=9
    -5, -14, -1, -9, -31, -7, -32, -26, -11,
    -- filter=75 channel=10
    12, 6, 13, 18, 7, 23, 0, 23, 13,
    -- filter=75 channel=11
    0, 13, -5, 14, 21, 0, 2, -10, -16,
    -- filter=75 channel=12
    -5, 7, 10, 2, 1, -2, -6, -10, -7,
    -- filter=75 channel=13
    6, -14, -3, -1, -1, 0, -3, -8, -19,
    -- filter=75 channel=14
    -1, 1, -6, 3, 5, -8, -5, 8, -6,
    -- filter=75 channel=15
    15, 6, 5, 0, -6, -16, -23, -24, -23,
    -- filter=75 channel=16
    15, 11, 9, 0, -3, 0, -23, -19, -19,
    -- filter=75 channel=17
    0, 14, -11, -10, 4, -5, -2, -5, -9,
    -- filter=75 channel=18
    -9, -18, -5, -4, -15, -20, -22, -15, -23,
    -- filter=75 channel=19
    -3, 11, 16, -7, 14, 10, -2, 0, -4,
    -- filter=75 channel=20
    8, -2, 5, -7, -1, 2, -1, -5, 9,
    -- filter=75 channel=21
    1, 3, -6, -2, -6, 4, 0, 2, 1,
    -- filter=75 channel=22
    0, 6, -9, 10, 10, -4, 5, 9, -5,
    -- filter=75 channel=23
    3, 24, 3, 11, 33, 16, 20, 11, 9,
    -- filter=75 channel=24
    -8, -7, 7, 4, -3, -3, -14, -10, -17,
    -- filter=75 channel=25
    31, 44, 20, 26, 43, 24, 8, 29, 15,
    -- filter=75 channel=26
    9, 14, 6, 18, 9, 8, 0, 13, -1,
    -- filter=75 channel=27
    25, 32, 3, 15, 38, 18, 10, 23, 0,
    -- filter=75 channel=28
    -4, 4, -13, -11, -24, -9, -17, -15, -9,
    -- filter=75 channel=29
    20, 8, -4, -12, -18, -15, -28, -34, -7,
    -- filter=75 channel=30
    14, 30, 16, 8, 35, 2, 4, 31, 2,
    -- filter=75 channel=31
    9, 8, -9, -3, 4, 8, 13, 6, 5,
    -- filter=75 channel=32
    12, 27, 10, 29, 36, 15, 23, 37, 11,
    -- filter=75 channel=33
    0, 8, 0, 0, -7, 3, -9, 5, -1,
    -- filter=75 channel=34
    0, 0, 0, -2, 11, 1, -3, 9, 7,
    -- filter=75 channel=35
    18, 48, 8, 29, 36, 32, 29, 33, 21,
    -- filter=75 channel=36
    -3, 5, 7, 8, -2, 14, 6, -2, 2,
    -- filter=75 channel=37
    -1, 5, 5, 2, 10, 6, -16, -13, 5,
    -- filter=75 channel=38
    16, 27, 11, 22, 22, 19, 8, 4, 5,
    -- filter=75 channel=39
    -3, 5, -5, -10, 4, -10, 3, 10, -9,
    -- filter=75 channel=40
    9, 18, 2, 1, 11, 9, 8, 13, 12,
    -- filter=75 channel=41
    7, 27, 14, 1, 4, 9, -19, -9, -17,
    -- filter=75 channel=42
    -5, 8, 7, 5, -6, 7, 7, -4, 2,
    -- filter=75 channel=43
    8, 23, 13, 30, 40, 32, 13, 29, 15,
    -- filter=75 channel=44
    14, 29, 15, 21, 26, 11, 17, 31, 12,
    -- filter=75 channel=45
    -1, -1, 3, 3, -7, -5, -5, -4, -2,
    -- filter=75 channel=46
    -1, -8, 7, 5, 0, 4, 3, -1, -8,
    -- filter=75 channel=47
    10, 3, 2, 7, -9, 0, -3, 8, 0,
    -- filter=75 channel=48
    9, -4, -12, 1, 0, -8, -15, -19, 0,
    -- filter=75 channel=49
    10, 11, 1, 8, 4, 0, 1, -2, 0,
    -- filter=75 channel=50
    -8, 13, 15, 13, 23, 1, 3, 6, 12,
    -- filter=75 channel=51
    -4, -4, 3, 0, 5, 6, 1, 13, 6,
    -- filter=75 channel=52
    -9, 2, 10, 9, -5, -9, 10, 0, 0,
    -- filter=75 channel=53
    4, 19, 20, 7, 36, 12, 21, 26, 6,
    -- filter=75 channel=54
    1, -6, 9, -16, -18, -6, -18, -17, 3,
    -- filter=75 channel=55
    -8, 4, 5, -2, 4, -2, -5, 5, -4,
    -- filter=75 channel=56
    2, 8, 9, 12, 8, 3, 12, 8, -3,
    -- filter=75 channel=57
    9, 0, 4, -8, 0, -10, 1, -1, 7,
    -- filter=75 channel=58
    -8, -7, 1, -6, 7, 0, -3, 4, 6,
    -- filter=75 channel=59
    21, 11, 16, 13, 16, -1, -9, -4, 11,
    -- filter=75 channel=60
    17, -2, -3, -9, -1, 1, -9, -16, -13,
    -- filter=75 channel=61
    6, 13, -1, 12, -2, 0, -16, -11, -16,
    -- filter=75 channel=62
    14, 3, 3, 14, 9, 3, 4, -5, -11,
    -- filter=75 channel=63
    -6, -7, 10, -3, 3, -5, 9, 1, 9,
    -- filter=76 channel=0
    -5, -11, -11, -4, -5, -10, 9, 0, -6,
    -- filter=76 channel=1
    -11, 5, 8, 1, 9, -3, 8, 3, -7,
    -- filter=76 channel=2
    -7, -6, -9, -12, -9, 0, -4, -5, -1,
    -- filter=76 channel=3
    4, 7, 1, -2, -4, -13, -11, -2, -10,
    -- filter=76 channel=4
    0, 10, -3, 13, 11, 7, 0, 4, 5,
    -- filter=76 channel=5
    7, 11, -9, 12, 13, 4, -6, -3, -2,
    -- filter=76 channel=6
    13, -4, -5, 3, 5, -1, -1, -1, -5,
    -- filter=76 channel=7
    -1, -4, 4, 8, 6, 5, -6, 2, 1,
    -- filter=76 channel=8
    5, 10, 0, -2, 15, 11, 1, 2, -8,
    -- filter=76 channel=9
    22, 45, 43, 41, 57, 46, 30, 61, 38,
    -- filter=76 channel=10
    11, 0, 0, -6, -8, -13, 0, 6, -6,
    -- filter=76 channel=11
    2, 6, -1, 2, -4, 4, -5, 5, 3,
    -- filter=76 channel=12
    -4, -5, 3, 0, 1, -1, -3, 9, -4,
    -- filter=76 channel=13
    2, 11, 7, 11, 15, 2, -1, 3, -7,
    -- filter=76 channel=14
    -2, -9, -11, 10, -6, -8, -3, -4, 4,
    -- filter=76 channel=15
    14, 6, -5, 0, -1, -12, 11, 0, -15,
    -- filter=76 channel=16
    5, 10, 4, -1, 14, 3, -4, 5, -1,
    -- filter=76 channel=17
    7, 11, -10, -4, -3, 0, 2, -7, -15,
    -- filter=76 channel=18
    25, 14, 19, 25, 28, 24, 27, 27, 20,
    -- filter=76 channel=19
    9, 17, 15, 11, 24, 19, 13, 7, 13,
    -- filter=76 channel=20
    15, 11, 10, 3, 12, 12, 13, 11, 12,
    -- filter=76 channel=21
    8, 0, 8, 9, -1, 11, 2, -6, -6,
    -- filter=76 channel=22
    -3, 7, 0, 0, -8, 10, -2, -4, -2,
    -- filter=76 channel=23
    -6, 0, -11, 5, -17, -4, -5, 4, 0,
    -- filter=76 channel=24
    -9, -4, -2, -1, -1, -2, 10, -8, -7,
    -- filter=76 channel=25
    -3, 0, -10, -12, -11, 0, -17, -22, -1,
    -- filter=76 channel=26
    -7, -4, 6, -10, 7, 6, -3, 6, -9,
    -- filter=76 channel=27
    -12, -8, -5, -12, -18, -3, -17, -21, -9,
    -- filter=76 channel=28
    0, 23, 9, 18, 24, 12, 2, 15, 3,
    -- filter=76 channel=29
    -9, 5, 4, 16, 9, 0, -3, 0, -4,
    -- filter=76 channel=30
    9, 2, -4, -3, -3, 2, 0, 3, 4,
    -- filter=76 channel=31
    -8, -6, 7, -9, -10, 10, 5, -7, -7,
    -- filter=76 channel=32
    -4, -13, 2, -4, 0, 4, -5, 6, 2,
    -- filter=76 channel=33
    -8, 10, 8, 10, 4, -4, 0, 1, -5,
    -- filter=76 channel=34
    -2, 8, 3, 1, 1, 9, 1, 3, -9,
    -- filter=76 channel=35
    -9, -10, 0, -15, -13, -21, -12, -16, -17,
    -- filter=76 channel=36
    -1, -6, 10, -8, -10, -9, -1, -6, 3,
    -- filter=76 channel=37
    8, 4, 8, 9, 13, 0, 4, 4, -3,
    -- filter=76 channel=38
    -1, -10, -14, 1, -17, -15, 0, -2, -6,
    -- filter=76 channel=39
    4, 5, -2, 9, 6, 9, -8, 8, -4,
    -- filter=76 channel=40
    -9, -11, 7, -5, -13, -4, -5, -11, -3,
    -- filter=76 channel=41
    3, -8, 3, -1, -3, -14, -9, -11, -21,
    -- filter=76 channel=42
    8, -1, 7, 3, 2, -7, -7, 10, -9,
    -- filter=76 channel=43
    -9, -16, -18, -14, -3, -14, 4, -14, 3,
    -- filter=76 channel=44
    -5, -1, 6, -7, -2, -3, -12, -5, 5,
    -- filter=76 channel=45
    6, 1, 10, 0, -6, 7, 4, -4, 0,
    -- filter=76 channel=46
    11, 3, -2, -3, -1, -4, -2, -3, -2,
    -- filter=76 channel=47
    7, -3, 9, 5, -7, -6, -5, -7, -7,
    -- filter=76 channel=48
    -4, 9, 4, -3, 6, -7, -8, -7, 0,
    -- filter=76 channel=49
    10, -5, -5, -5, 0, 7, 0, -11, 9,
    -- filter=76 channel=50
    4, 12, 4, 14, 8, -2, 11, 13, -4,
    -- filter=76 channel=51
    2, 4, 13, 6, -8, -9, 6, 3, 9,
    -- filter=76 channel=52
    -8, -5, 8, 0, -2, -9, 7, 4, 4,
    -- filter=76 channel=53
    6, -12, 0, 4, -1, 2, -5, 1, -3,
    -- filter=76 channel=54
    14, 34, 29, 20, 50, 41, 26, 37, 28,
    -- filter=76 channel=55
    0, 6, -8, 1, -7, 7, -10, 0, -8,
    -- filter=76 channel=56
    -10, -2, 6, -7, 3, -5, 8, 1, 9,
    -- filter=76 channel=57
    0, -5, 2, 3, -9, 4, -9, -6, -7,
    -- filter=76 channel=58
    21, 16, 6, 9, 4, 11, 12, 8, 12,
    -- filter=76 channel=59
    -11, -7, -1, -15, -15, -4, -15, -13, -13,
    -- filter=76 channel=60
    -6, 7, -4, 5, 11, -11, -5, 0, -17,
    -- filter=76 channel=61
    -4, -9, -5, 5, 3, -7, 5, 0, -19,
    -- filter=76 channel=62
    2, 3, -1, -3, 7, -9, -3, -6, -11,
    -- filter=76 channel=63
    9, 6, -4, 2, 7, -5, -9, 4, -9,
    -- filter=77 channel=0
    3, -3, 10, -2, 9, -2, 11, 5, 8,
    -- filter=77 channel=1
    -7, -8, 2, 7, 1, -6, -4, -2, -8,
    -- filter=77 channel=2
    2, -6, 3, -5, 3, -4, 9, -2, 1,
    -- filter=77 channel=3
    -2, 0, 2, -9, -6, -5, 5, -9, -3,
    -- filter=77 channel=4
    -10, 7, 0, -7, -6, -6, 3, 10, -2,
    -- filter=77 channel=5
    -10, 0, 7, 0, 9, -3, 0, -1, -3,
    -- filter=77 channel=6
    -5, 5, -8, -3, 11, 5, -5, -9, 0,
    -- filter=77 channel=7
    5, 1, 10, 7, 3, -8, -2, -6, 7,
    -- filter=77 channel=8
    5, -10, -4, 3, 0, -7, -7, 6, -4,
    -- filter=77 channel=9
    -4, 0, -1, -9, 2, 10, -11, 0, 4,
    -- filter=77 channel=10
    1, -9, -7, 6, 11, -8, 4, 6, 7,
    -- filter=77 channel=11
    3, 7, -3, -7, -9, -6, 8, -8, 3,
    -- filter=77 channel=12
    -2, -4, 0, -9, -2, 9, -1, -4, -9,
    -- filter=77 channel=13
    6, 9, 3, -4, -5, 3, 8, -3, -8,
    -- filter=77 channel=14
    -6, -9, 9, -4, 6, 3, 8, 0, 1,
    -- filter=77 channel=15
    -3, 7, -11, -2, 3, -11, 1, -4, -10,
    -- filter=77 channel=16
    2, -7, -2, 8, 2, -11, 4, -8, -13,
    -- filter=77 channel=17
    -10, -1, 8, -9, 6, -3, 9, -2, -6,
    -- filter=77 channel=18
    9, 1, -5, -6, 0, -4, 5, 11, 5,
    -- filter=77 channel=19
    -7, -5, 3, -3, 6, 5, 11, 9, 0,
    -- filter=77 channel=20
    6, 0, 7, -8, -8, -5, -7, 2, -7,
    -- filter=77 channel=21
    -6, 0, 9, 8, -5, 5, 6, -2, -3,
    -- filter=77 channel=22
    -1, 1, -7, 4, 0, -1, 0, -2, 0,
    -- filter=77 channel=23
    -5, 4, -8, 8, -4, -4, 5, -6, 0,
    -- filter=77 channel=24
    -1, 4, 0, 0, 5, 6, 5, 0, -10,
    -- filter=77 channel=25
    -5, -3, -7, 6, 9, 3, -6, -4, -10,
    -- filter=77 channel=26
    -4, 0, 0, 8, 1, 9, -8, -2, -5,
    -- filter=77 channel=27
    -11, -9, 2, 2, -7, 7, -3, -7, -8,
    -- filter=77 channel=28
    8, -1, 8, 8, -1, -9, 8, 6, -9,
    -- filter=77 channel=29
    -12, -10, -10, 6, 6, -3, 6, 8, 5,
    -- filter=77 channel=30
    4, 3, 10, -9, 0, 0, 0, -6, 3,
    -- filter=77 channel=31
    1, -2, -8, -9, 0, -5, -6, 1, -3,
    -- filter=77 channel=32
    0, 5, -10, -9, 1, 8, 5, -6, 11,
    -- filter=77 channel=33
    6, -9, 2, 2, -6, -9, 6, 9, -7,
    -- filter=77 channel=34
    -2, -2, -5, 4, -5, -4, -8, -7, 7,
    -- filter=77 channel=35
    -10, -3, 6, -8, -5, 7, 8, 11, -2,
    -- filter=77 channel=36
    3, 3, 0, 8, 10, 5, 2, -6, 0,
    -- filter=77 channel=37
    9, 4, 7, -3, 6, -6, -7, -10, 3,
    -- filter=77 channel=38
    -2, 4, 3, 10, 10, -1, -5, -8, -11,
    -- filter=77 channel=39
    -10, 6, 5, 3, -7, -7, -7, -6, 9,
    -- filter=77 channel=40
    -1, 2, 7, -4, 8, -8, 6, 8, -4,
    -- filter=77 channel=41
    -12, 8, 1, -2, -9, -2, -3, -4, -5,
    -- filter=77 channel=42
    -10, -9, 2, -10, -8, -4, 3, 6, 3,
    -- filter=77 channel=43
    -6, -7, 1, 5, 2, 8, -8, 7, 4,
    -- filter=77 channel=44
    9, 5, -2, 5, 0, -4, -3, 0, 5,
    -- filter=77 channel=45
    -9, 9, 7, 9, -5, 9, 7, 3, -10,
    -- filter=77 channel=46
    -3, 1, 11, 3, -9, 0, 9, 5, -3,
    -- filter=77 channel=47
    10, -4, -9, 0, -8, 4, 1, 6, -3,
    -- filter=77 channel=48
    4, 8, -10, -5, 0, -9, -8, 0, -6,
    -- filter=77 channel=49
    6, 9, 0, 11, 6, 8, 9, 7, -7,
    -- filter=77 channel=50
    8, -1, -6, 4, 2, -6, 4, 2, 3,
    -- filter=77 channel=51
    10, -2, 8, -7, 7, 1, -2, 7, 0,
    -- filter=77 channel=52
    8, 8, 0, 5, 0, -10, 7, -1, 6,
    -- filter=77 channel=53
    4, -3, -4, 8, 6, 3, 4, 1, 0,
    -- filter=77 channel=54
    0, 9, -4, 7, -9, 6, 8, 4, 2,
    -- filter=77 channel=55
    -5, -2, -2, -1, -7, 8, -3, -2, 6,
    -- filter=77 channel=56
    9, 6, -3, 5, -9, -5, -3, 8, 2,
    -- filter=77 channel=57
    -9, -9, 6, -3, -2, -7, 0, 3, 6,
    -- filter=77 channel=58
    2, 7, 8, -3, -8, 2, 5, -7, 8,
    -- filter=77 channel=59
    0, 8, 7, 7, 1, -5, 2, -3, 4,
    -- filter=77 channel=60
    -9, 3, 3, -7, 9, -9, 12, 4, -3,
    -- filter=77 channel=61
    -1, -10, 4, 3, -2, -1, -1, 11, -7,
    -- filter=77 channel=62
    5, -10, 9, -9, 7, 10, 3, 9, 0,
    -- filter=77 channel=63
    1, 6, 2, 0, -9, 3, -1, -7, -6,
    -- filter=78 channel=0
    -2, 4, 3, 0, 0, 8, 10, 2, 3,
    -- filter=78 channel=1
    3, 5, -12, -1, -2, -11, 2, 5, -3,
    -- filter=78 channel=2
    -4, -3, -8, -14, -13, 7, -2, -3, 1,
    -- filter=78 channel=3
    3, 2, 3, -4, 5, 2, 0, 5, 8,
    -- filter=78 channel=4
    4, -3, 7, 5, 2, 9, -11, 3, 5,
    -- filter=78 channel=5
    -10, 4, 2, -4, 6, 6, -1, -4, -1,
    -- filter=78 channel=6
    -5, 3, 1, -1, 0, -1, 0, 1, -6,
    -- filter=78 channel=7
    -5, 0, 7, -7, 7, 0, 1, -3, 5,
    -- filter=78 channel=8
    1, -12, -1, 0, -10, -5, 4, 3, -2,
    -- filter=78 channel=9
    -2, -1, 14, 0, 1, 5, -12, -8, -1,
    -- filter=78 channel=10
    -3, 11, 5, 6, 9, 1, 5, 6, 10,
    -- filter=78 channel=11
    4, -3, -3, 0, 0, -6, 3, -6, 7,
    -- filter=78 channel=12
    10, 2, 0, -1, 1, -2, -8, 1, 8,
    -- filter=78 channel=13
    -6, -6, 12, 3, -6, -2, -6, -5, -8,
    -- filter=78 channel=14
    6, -1, -5, 4, -7, -3, 1, 5, 7,
    -- filter=78 channel=15
    -2, 2, 5, -6, 1, 2, 3, -5, -3,
    -- filter=78 channel=16
    -16, -13, 10, -15, -18, -1, -17, -12, -10,
    -- filter=78 channel=17
    0, -12, 8, -11, 0, 2, 5, 0, 3,
    -- filter=78 channel=18
    -6, -3, 7, -1, -2, 10, -2, 3, 9,
    -- filter=78 channel=19
    -13, -15, -4, -17, -1, -8, 0, -14, -12,
    -- filter=78 channel=20
    -9, 5, 8, 5, 0, -2, 3, -1, -9,
    -- filter=78 channel=21
    -2, 1, -1, 8, 1, 5, 1, -1, -7,
    -- filter=78 channel=22
    5, -8, -10, -3, 1, 9, 1, -4, -2,
    -- filter=78 channel=23
    4, 10, -5, -1, 12, 15, 13, 12, 7,
    -- filter=78 channel=24
    -7, -8, 10, 6, -7, -6, -5, -11, 0,
    -- filter=78 channel=25
    4, -8, 4, 3, 4, 0, -5, 7, 5,
    -- filter=78 channel=26
    2, -7, 10, 3, -8, -4, 1, -7, 0,
    -- filter=78 channel=27
    -9, 13, 2, 1, 12, 7, -2, 11, 13,
    -- filter=78 channel=28
    -8, -9, 0, -21, -17, -11, -6, -3, -9,
    -- filter=78 channel=29
    -13, -1, 7, -16, -21, 10, -17, -18, -13,
    -- filter=78 channel=30
    -13, -12, -3, 3, 2, 2, -4, 0, 0,
    -- filter=78 channel=31
    -1, -1, 1, 0, -7, 5, 13, 12, 6,
    -- filter=78 channel=32
    10, 14, 0, 12, 15, 3, 14, 13, 3,
    -- filter=78 channel=33
    -7, -1, 6, -6, -2, -8, -10, -10, 9,
    -- filter=78 channel=34
    2, -6, -1, -2, 0, 6, 6, -11, 1,
    -- filter=78 channel=35
    0, 20, 6, 4, 17, 5, 18, 17, 8,
    -- filter=78 channel=36
    11, -4, -1, 1, 10, 9, 8, 12, -3,
    -- filter=78 channel=37
    -7, -8, -8, 7, -11, -8, 7, -2, -1,
    -- filter=78 channel=38
    4, 5, 8, 2, 8, 15, 3, -1, 7,
    -- filter=78 channel=39
    1, -9, 9, -5, -9, -3, 2, 4, -7,
    -- filter=78 channel=40
    1, 10, 12, 7, 5, 12, -6, -5, 12,
    -- filter=78 channel=41
    7, -9, 20, 5, 6, 0, -3, -5, 8,
    -- filter=78 channel=42
    9, 8, -2, 6, -9, 10, -2, 9, -8,
    -- filter=78 channel=43
    -11, 4, 1, -10, 0, -10, 3, -10, 7,
    -- filter=78 channel=44
    -7, 1, 7, 4, -1, -2, -2, 5, 0,
    -- filter=78 channel=45
    -8, -2, 2, 5, -3, -10, -1, 6, 0,
    -- filter=78 channel=46
    2, 9, 11, 0, 3, -7, 9, 7, -9,
    -- filter=78 channel=47
    -1, -8, -10, 9, -6, -7, 2, 0, 9,
    -- filter=78 channel=48
    3, 1, 7, -12, -11, 4, -11, -10, -2,
    -- filter=78 channel=49
    12, 8, -1, 15, 12, 3, 14, 0, 2,
    -- filter=78 channel=50
    0, -1, -14, 2, 4, -5, 0, 0, -9,
    -- filter=78 channel=51
    9, 16, 2, 7, 11, 3, 5, 11, 13,
    -- filter=78 channel=52
    -9, -5, -1, -2, -9, 6, -7, 6, -5,
    -- filter=78 channel=53
    -8, 8, -12, 4, -5, -1, -5, 4, -7,
    -- filter=78 channel=54
    -2, 9, 0, 8, -2, 11, 8, -8, 0,
    -- filter=78 channel=55
    2, 4, -8, -6, 3, 9, -2, -8, 0,
    -- filter=78 channel=56
    -7, -1, -9, -3, -7, -5, -6, 8, 4,
    -- filter=78 channel=57
    3, 4, 0, 8, -8, 2, -10, 8, -6,
    -- filter=78 channel=58
    9, 3, 7, -9, -10, 3, 8, -6, -4,
    -- filter=78 channel=59
    0, -9, 16, 7, 5, 13, 2, -9, 0,
    -- filter=78 channel=60
    -8, -1, 21, -5, 10, 12, 0, -1, 5,
    -- filter=78 channel=61
    -10, 12, 12, 6, 3, 13, 0, 0, -5,
    -- filter=78 channel=62
    -6, 7, 9, 0, 0, 9, -1, -5, -4,
    -- filter=78 channel=63
    4, -10, -5, 7, -1, 0, 3, 1, 4,
    -- filter=79 channel=0
    -2, -19, -7, 0, -7, -11, 0, -13, -22,
    -- filter=79 channel=1
    -1, 22, 24, 10, 31, 23, 11, 27, 24,
    -- filter=79 channel=2
    14, 23, 27, 10, 31, 34, -11, 18, 13,
    -- filter=79 channel=3
    23, 39, 24, 28, 37, 26, 21, 26, 0,
    -- filter=79 channel=4
    -9, -15, -14, -6, -9, -14, -7, -11, -13,
    -- filter=79 channel=5
    18, 14, 0, 11, 27, 4, 2, 1, 5,
    -- filter=79 channel=6
    8, 7, 0, 11, 1, -9, -5, 3, 3,
    -- filter=79 channel=7
    -2, 8, 3, 3, 1, 4, 0, 2, 4,
    -- filter=79 channel=8
    8, 10, -16, 0, 1, -2, -13, -24, -15,
    -- filter=79 channel=9
    -9, 17, 2, 7, 27, 12, 7, 19, 13,
    -- filter=79 channel=10
    -15, -21, -3, 0, -13, -5, 2, 0, -2,
    -- filter=79 channel=11
    -8, 3, 5, 5, 0, 2, -3, -7, 1,
    -- filter=79 channel=12
    8, 6, 0, -8, -4, 0, 9, 4, 7,
    -- filter=79 channel=13
    0, 3, -7, 12, 19, 1, 6, 14, -4,
    -- filter=79 channel=14
    4, -5, -7, 9, -1, 1, 7, 10, -1,
    -- filter=79 channel=15
    7, 1, -17, 10, 7, -6, -17, -1, -31,
    -- filter=79 channel=16
    7, 18, 16, 25, 26, 12, -3, 5, -4,
    -- filter=79 channel=17
    -11, 9, -11, 8, 9, 4, -2, -9, -7,
    -- filter=79 channel=18
    -2, -5, -26, -9, -13, -11, -9, -17, -16,
    -- filter=79 channel=19
    16, 28, 7, 5, 36, 29, 16, 20, 23,
    -- filter=79 channel=20
    3, 2, 6, 9, 7, -4, 8, 9, 9,
    -- filter=79 channel=21
    2, 9, 1, -6, -8, -4, 6, -7, 1,
    -- filter=79 channel=22
    0, -5, -5, -8, 0, 9, 5, 1, -7,
    -- filter=79 channel=23
    -22, -5, -3, -9, -7, -10, -14, 0, -10,
    -- filter=79 channel=24
    -11, 3, 1, 0, 9, 3, -14, -3, -4,
    -- filter=79 channel=25
    5, 33, 17, 20, 43, 31, 1, 10, 29,
    -- filter=79 channel=26
    13, 11, -9, 4, 9, -7, 6, 7, 13,
    -- filter=79 channel=27
    4, 20, 5, 3, 8, 13, -9, -1, 8,
    -- filter=79 channel=28
    0, 23, -6, 1, 10, 8, -3, -3, -6,
    -- filter=79 channel=29
    18, 30, 0, 18, 41, -3, 9, 9, -21,
    -- filter=79 channel=30
    14, 13, 6, 4, 24, 4, 17, 28, 0,
    -- filter=79 channel=31
    -8, -4, 5, 5, -8, 2, 4, -5, -3,
    -- filter=79 channel=32
    1, 3, 1, 0, 1, 19, -12, -1, 14,
    -- filter=79 channel=33
    -5, 5, 3, -7, 9, 8, 4, 9, -6,
    -- filter=79 channel=34
    8, 13, 0, -4, -1, 9, -2, 1, 0,
    -- filter=79 channel=35
    -8, 12, 8, -11, -2, -3, -26, -3, -8,
    -- filter=79 channel=36
    -2, 0, 10, -10, -2, 8, 1, -4, 0,
    -- filter=79 channel=37
    18, 17, 5, 4, 23, 12, 0, 20, 8,
    -- filter=79 channel=38
    2, 15, -10, 4, 16, 1, 1, 3, -5,
    -- filter=79 channel=39
    -7, -5, 3, 0, -1, -4, -2, -7, -7,
    -- filter=79 channel=40
    9, 0, 9, -2, 10, -3, 3, 1, 0,
    -- filter=79 channel=41
    17, 7, -12, 16, 28, 0, -18, -3, -12,
    -- filter=79 channel=42
    -1, 10, 0, -4, 4, 8, -6, 6, -1,
    -- filter=79 channel=43
    -14, -21, -6, 0, 19, 8, -2, 3, 17,
    -- filter=79 channel=44
    9, 11, 12, 8, 11, 28, 6, 12, 9,
    -- filter=79 channel=45
    -3, 0, 7, 8, 4, 5, 6, -5, -4,
    -- filter=79 channel=46
    15, 0, -11, 5, 13, -7, 12, 16, 6,
    -- filter=79 channel=47
    -8, 0, 5, 6, 5, 1, 6, -4, 5,
    -- filter=79 channel=48
    15, 2, 9, 12, 15, 10, -5, 9, -8,
    -- filter=79 channel=49
    2, 3, -3, -3, -11, -4, -19, -15, -21,
    -- filter=79 channel=50
    1, 11, 6, 13, 11, 7, 0, 3, 7,
    -- filter=79 channel=51
    -2, -29, -9, -5, -24, -28, 1, -18, -9,
    -- filter=79 channel=52
    -8, 5, -9, -2, -2, -6, 1, -9, 2,
    -- filter=79 channel=53
    -1, 14, 9, 4, 5, 18, 4, 12, 18,
    -- filter=79 channel=54
    0, 23, 18, 14, 34, 18, 3, 3, 7,
    -- filter=79 channel=55
    -7, 6, 3, -7, 5, 9, -5, 0, 9,
    -- filter=79 channel=56
    10, 4, 3, -5, 2, 7, -3, -1, 6,
    -- filter=79 channel=57
    -1, 0, -1, 2, 10, 2, 0, 7, 7,
    -- filter=79 channel=58
    18, 0, 10, 18, 5, 2, 11, 16, 14,
    -- filter=79 channel=59
    17, 29, 7, 16, 17, 15, -6, 11, -2,
    -- filter=79 channel=60
    7, -3, -34, 4, 6, -22, -18, -2, -28,
    -- filter=79 channel=61
    -9, -6, -20, -16, 1, -8, -19, -21, -8,
    -- filter=79 channel=62
    1, 22, 19, 2, 15, 24, -5, 19, 11,
    -- filter=79 channel=63
    -9, 0, 10, 9, -4, 4, 0, 5, -6,
    -- filter=80 channel=0
    1, 3, 2, 9, 31, 18, 3, 10, 5,
    -- filter=80 channel=1
    0, -7, -18, -1, -1, -4, 2, -16, -10,
    -- filter=80 channel=2
    0, -12, -20, 0, -12, -22, -10, -16, -30,
    -- filter=80 channel=3
    6, 5, -10, -6, -2, -2, -9, -13, -8,
    -- filter=80 channel=4
    0, 18, 8, 18, 21, 3, -8, 14, 3,
    -- filter=80 channel=5
    9, -5, -6, 7, -12, 1, -5, -7, -9,
    -- filter=80 channel=6
    -5, 5, -7, 4, -1, 1, -4, 5, -6,
    -- filter=80 channel=7
    -6, -18, 1, 2, -3, -5, -16, -13, -1,
    -- filter=80 channel=8
    3, 19, -3, 29, 39, 7, 8, 13, -1,
    -- filter=80 channel=9
    -1, -16, -13, -12, -26, -31, 7, -13, -24,
    -- filter=80 channel=10
    -3, 11, 1, 8, 0, 18, 8, 0, 6,
    -- filter=80 channel=11
    -4, -3, 4, 6, 22, 10, 3, 2, 10,
    -- filter=80 channel=12
    11, 1, 7, 5, 5, 10, -3, -6, 9,
    -- filter=80 channel=13
    -5, 11, -11, 11, 15, -1, 5, 5, 3,
    -- filter=80 channel=14
    -9, -7, -7, -12, -5, 0, -11, -1, 4,
    -- filter=80 channel=15
    9, 5, -13, 20, 18, 12, 2, 8, -11,
    -- filter=80 channel=16
    19, -6, -17, 21, 1, -14, 0, -10, -24,
    -- filter=80 channel=17
    0, 7, -2, -1, 14, 22, 0, 7, 5,
    -- filter=80 channel=18
    11, 19, -2, 10, 28, 8, 10, 10, -4,
    -- filter=80 channel=19
    -14, -25, -14, -3, -11, -13, 1, -5, -6,
    -- filter=80 channel=20
    -10, -21, -23, -9, -7, -10, -6, -5, -11,
    -- filter=80 channel=21
    8, -1, 9, -2, 6, 10, 7, 2, 10,
    -- filter=80 channel=22
    -11, 4, 0, -9, 9, -3, 6, 8, -6,
    -- filter=80 channel=23
    -7, 10, 15, -5, 22, 25, -4, 7, 12,
    -- filter=80 channel=24
    13, 12, 0, 1, 18, 17, -1, 11, 18,
    -- filter=80 channel=25
    3, -18, -23, -10, -5, -16, -14, -15, -32,
    -- filter=80 channel=26
    -17, -26, -16, -16, -28, -7, -19, -11, -20,
    -- filter=80 channel=27
    9, 16, -8, 11, 22, 3, -7, 4, 5,
    -- filter=80 channel=28
    13, 10, -13, 2, 3, 6, -10, 4, 1,
    -- filter=80 channel=29
    3, 4, -15, 14, 9, -19, 5, -8, -15,
    -- filter=80 channel=30
    -33, -38, -13, -23, -30, -12, -32, -27, -11,
    -- filter=80 channel=31
    0, -5, 3, 0, -9, -6, 1, 11, -5,
    -- filter=80 channel=32
    -11, 0, -11, -13, -15, -13, -7, 1, 0,
    -- filter=80 channel=33
    7, 5, 6, 9, 10, 9, -4, 1, 1,
    -- filter=80 channel=34
    2, -3, -1, 0, -11, 0, -12, -15, -5,
    -- filter=80 channel=35
    -3, 21, -3, 9, 8, 13, -14, 1, -6,
    -- filter=80 channel=36
    -1, -8, 0, 4, 4, -6, 9, 11, 11,
    -- filter=80 channel=37
    -7, -18, -18, -1, 1, 0, -13, -12, -7,
    -- filter=80 channel=38
    0, 14, -11, 10, 12, 2, 10, 9, -3,
    -- filter=80 channel=39
    3, -8, 9, -6, 1, 10, -2, 5, 0,
    -- filter=80 channel=40
    4, 3, -3, -8, -1, 0, -14, -7, -12,
    -- filter=80 channel=41
    6, 18, 6, 25, 20, 13, -4, 18, -10,
    -- filter=80 channel=42
    9, 1, 0, -1, 10, 10, 0, -1, -3,
    -- filter=80 channel=43
    -43, -46, -26, -40, -43, -28, -19, -22, -11,
    -- filter=80 channel=44
    -15, -10, -2, -7, -13, -17, -22, -17, -8,
    -- filter=80 channel=45
    2, 8, 9, -10, -2, 3, -10, 0, 3,
    -- filter=80 channel=46
    -10, -8, -8, 0, -5, -15, -15, -9, -4,
    -- filter=80 channel=47
    -10, -7, 1, 0, -3, -5, 5, 9, -2,
    -- filter=80 channel=48
    8, 1, -19, 6, -9, -14, -10, 5, -10,
    -- filter=80 channel=49
    4, 17, 17, 20, 28, 23, 3, 12, 15,
    -- filter=80 channel=50
    -18, -19, -16, -32, -33, -8, -3, -20, -8,
    -- filter=80 channel=51
    0, 26, 24, 19, 29, 20, 11, 28, 22,
    -- filter=80 channel=52
    -7, 5, 8, 7, 8, 8, -2, 2, -8,
    -- filter=80 channel=53
    -6, -26, -12, -27, -29, -2, -29, -20, -4,
    -- filter=80 channel=54
    0, -24, -7, -17, -13, -13, -13, -21, -17,
    -- filter=80 channel=55
    -1, 10, -1, -8, -9, -10, -6, 0, -6,
    -- filter=80 channel=56
    -10, 2, -1, -12, 0, -11, 6, -11, -6,
    -- filter=80 channel=57
    -8, -10, 5, -1, 6, -1, 0, 10, 3,
    -- filter=80 channel=58
    -9, -8, 3, -11, -14, 2, -10, -4, 2,
    -- filter=80 channel=59
    -3, -2, -18, 9, 5, 3, 4, -5, 0,
    -- filter=80 channel=60
    6, 23, 0, 21, 50, 3, 5, 24, -7,
    -- filter=80 channel=61
    14, 17, 17, 24, 44, 29, 7, 30, 23,
    -- filter=80 channel=62
    12, 8, -5, 3, 8, 0, 4, 3, -4,
    -- filter=80 channel=63
    -6, -3, -1, 2, -1, 7, 7, -7, -7,
    -- filter=81 channel=0
    -8, 10, 1, 1, 7, -1, 6, 6, 2,
    -- filter=81 channel=1
    -10, -9, 0, 8, 10, -3, 6, 9, 9,
    -- filter=81 channel=2
    3, -9, -8, 4, 0, 2, 6, -4, 7,
    -- filter=81 channel=3
    -4, 1, 0, 7, -7, 5, 7, 5, -9,
    -- filter=81 channel=4
    -6, 0, 2, 7, -3, -8, -9, 4, 9,
    -- filter=81 channel=5
    -5, 3, -7, 5, -4, 3, -8, -3, -9,
    -- filter=81 channel=6
    9, -4, -3, -4, -7, 1, 0, -9, 1,
    -- filter=81 channel=7
    -1, -3, -4, 0, 0, 6, -3, -6, 8,
    -- filter=81 channel=8
    4, 0, -10, -1, 5, 0, -4, -9, 0,
    -- filter=81 channel=9
    -6, 1, 1, -8, -9, -3, 0, -10, 9,
    -- filter=81 channel=10
    4, -8, -8, 1, 1, 8, 4, 7, 0,
    -- filter=81 channel=11
    0, 0, 5, -4, -10, -7, 2, -5, 7,
    -- filter=81 channel=12
    7, 8, 10, 8, -5, 10, 9, -9, 0,
    -- filter=81 channel=13
    6, -5, 5, 4, -6, -1, -10, -9, 9,
    -- filter=81 channel=14
    -3, 8, 7, -4, -6, 0, 1, -1, 0,
    -- filter=81 channel=15
    2, -10, -5, -3, 7, 8, -8, 9, -10,
    -- filter=81 channel=16
    -1, 2, 0, -2, -4, -5, -3, -4, -9,
    -- filter=81 channel=17
    8, -9, 0, -3, 9, -3, -1, 6, 0,
    -- filter=81 channel=18
    -3, -2, -10, 10, -6, 5, -5, 8, -8,
    -- filter=81 channel=19
    -5, 1, 5, -8, -10, -7, -9, 3, -10,
    -- filter=81 channel=20
    1, -7, -9, -1, 0, -6, -2, 4, 0,
    -- filter=81 channel=21
    -5, 7, -8, 3, 4, 6, -2, -2, 0,
    -- filter=81 channel=22
    -1, 4, 1, 0, -6, -2, 1, 0, -9,
    -- filter=81 channel=23
    -5, -10, -10, 2, -10, 9, 7, -11, 3,
    -- filter=81 channel=24
    5, 5, -1, 6, -10, 7, 9, 5, -1,
    -- filter=81 channel=25
    5, 0, 6, 0, 2, 10, -10, 1, 7,
    -- filter=81 channel=26
    -6, -3, -1, 3, -7, 5, -6, -5, -8,
    -- filter=81 channel=27
    -7, -3, -7, -1, 5, -8, -5, -2, -7,
    -- filter=81 channel=28
    2, 0, -7, 7, 8, 6, 2, -6, -10,
    -- filter=81 channel=29
    9, -2, 4, 0, -6, 4, 2, -7, -10,
    -- filter=81 channel=30
    -7, 10, 0, 1, -2, 6, -3, 1, 3,
    -- filter=81 channel=31
    -6, -3, -10, 2, -3, -6, -4, 0, 8,
    -- filter=81 channel=32
    -2, 4, 0, -3, -9, -4, -10, 10, -4,
    -- filter=81 channel=33
    -4, -4, 2, 7, 0, 2, -4, 2, -8,
    -- filter=81 channel=34
    -8, 10, -1, -1, -9, -2, 1, -10, -1,
    -- filter=81 channel=35
    -9, -5, 3, 6, 0, 0, 6, -5, 2,
    -- filter=81 channel=36
    0, -8, 0, -8, 5, -3, 7, 10, 8,
    -- filter=81 channel=37
    0, 6, 0, -10, 4, -3, 0, 3, -9,
    -- filter=81 channel=38
    0, -3, -2, -8, -7, 5, 0, -5, 7,
    -- filter=81 channel=39
    3, 2, -10, -9, 4, -10, -8, 9, 8,
    -- filter=81 channel=40
    -1, 7, 5, 2, 10, 8, -1, 5, 6,
    -- filter=81 channel=41
    -3, 4, -7, -6, -8, -10, -5, -6, 1,
    -- filter=81 channel=42
    0, -5, 10, -4, 6, -4, -3, 0, 1,
    -- filter=81 channel=43
    -4, 10, 1, 8, -5, -3, -3, 5, -9,
    -- filter=81 channel=44
    -6, 8, 8, -5, -4, 2, -8, 10, -7,
    -- filter=81 channel=45
    -3, 9, -7, -3, 7, -3, -5, 4, 6,
    -- filter=81 channel=46
    -5, 4, -5, 4, 6, 8, -6, -5, 0,
    -- filter=81 channel=47
    4, -8, 8, 0, -2, -5, 4, 9, 5,
    -- filter=81 channel=48
    3, 4, -8, -7, 6, -6, 6, -1, 10,
    -- filter=81 channel=49
    0, -2, 9, 9, 0, -1, -2, -6, 0,
    -- filter=81 channel=50
    -2, -1, 0, 6, 1, -8, 0, -2, 3,
    -- filter=81 channel=51
    -2, 3, -1, 8, 1, 8, 4, 4, 9,
    -- filter=81 channel=52
    4, -10, -8, 7, 2, -9, -7, -5, 4,
    -- filter=81 channel=53
    -5, 6, -9, 5, 5, 6, 1, -5, 2,
    -- filter=81 channel=54
    10, -3, -4, -10, -2, 1, 9, -8, -6,
    -- filter=81 channel=55
    2, 7, -4, -6, 5, -1, 4, -9, -4,
    -- filter=81 channel=56
    10, -3, 1, -9, 0, -10, -9, -7, 8,
    -- filter=81 channel=57
    -4, 0, 2, 6, 5, 8, -1, 0, 4,
    -- filter=81 channel=58
    0, 9, 5, 6, 0, -6, -4, -8, -3,
    -- filter=81 channel=59
    6, -8, 7, -6, -1, 4, 0, -4, 9,
    -- filter=81 channel=60
    -5, 6, 3, 4, 2, 1, 0, -4, 7,
    -- filter=81 channel=61
    8, -8, -10, -6, -3, 0, 1, -4, 6,
    -- filter=81 channel=62
    -10, -6, 2, -2, 10, -8, 1, 1, -7,
    -- filter=81 channel=63
    0, 1, 3, -9, 6, 8, -1, -4, 4,
    -- filter=82 channel=0
    0, -5, 2, 4, -5, 0, 9, -11, 6,
    -- filter=82 channel=1
    0, 5, -4, 6, 0, -5, 0, 7, 1,
    -- filter=82 channel=2
    5, -1, -5, -9, 1, 0, -2, -4, -10,
    -- filter=82 channel=3
    -8, -6, 3, 7, -11, -4, -4, 8, -3,
    -- filter=82 channel=4
    1, 1, 10, 1, 0, -3, -6, 4, 3,
    -- filter=82 channel=5
    8, 1, -10, -2, -12, 8, 2, -9, 0,
    -- filter=82 channel=6
    0, -9, 9, 5, -7, -7, -6, 0, 4,
    -- filter=82 channel=7
    -5, -9, -8, -9, 1, 0, -8, -5, 5,
    -- filter=82 channel=8
    10, 3, 7, -5, 0, -8, -2, -10, -9,
    -- filter=82 channel=9
    -4, 4, 9, 7, -5, 3, 0, 7, 1,
    -- filter=82 channel=10
    9, 4, 8, 9, 0, 8, -2, 7, -6,
    -- filter=82 channel=11
    10, 0, 8, 4, 0, 3, -6, 7, -1,
    -- filter=82 channel=12
    -8, 7, -9, -5, 0, -5, -5, 4, -7,
    -- filter=82 channel=13
    8, -4, 5, 8, 2, 6, 6, 6, 4,
    -- filter=82 channel=14
    -9, 5, 4, 1, 3, -5, 7, 8, -7,
    -- filter=82 channel=15
    -2, 4, -1, -11, 4, -3, -3, 3, 8,
    -- filter=82 channel=16
    7, -2, 10, -3, -11, 0, -1, -6, -13,
    -- filter=82 channel=17
    -3, 0, 9, 5, 2, 5, 4, -11, -5,
    -- filter=82 channel=18
    3, -5, -5, 4, 0, 4, 12, 4, 8,
    -- filter=82 channel=19
    3, 2, 2, 6, 7, -1, -2, 0, 4,
    -- filter=82 channel=20
    0, 6, -6, -8, -4, 3, -2, -2, 0,
    -- filter=82 channel=21
    2, 9, -3, 8, -9, -3, 6, 8, -2,
    -- filter=82 channel=22
    -3, -2, 0, 0, -8, -1, -5, -6, -8,
    -- filter=82 channel=23
    1, -5, 5, 10, 8, -5, 2, 1, 2,
    -- filter=82 channel=24
    12, 5, -5, -3, 0, -3, 0, -2, -7,
    -- filter=82 channel=25
    -4, 8, 11, -7, 7, 1, -9, 7, 9,
    -- filter=82 channel=26
    -2, 4, -7, 9, 5, 4, 6, -2, 0,
    -- filter=82 channel=27
    12, 8, -1, -4, 6, 9, -11, 2, 0,
    -- filter=82 channel=28
    9, -5, 0, 3, 3, 5, -10, -8, -4,
    -- filter=82 channel=29
    8, 12, 16, -10, -2, 2, 3, -17, -2,
    -- filter=82 channel=30
    -6, 0, -8, -10, 4, -8, -12, -2, 8,
    -- filter=82 channel=31
    -3, 3, -10, 10, 0, 6, -3, 2, -4,
    -- filter=82 channel=32
    0, 10, 1, -6, 4, 0, -4, -3, 10,
    -- filter=82 channel=33
    6, -1, 2, -9, -10, -6, 3, -4, 8,
    -- filter=82 channel=34
    9, 4, -3, 9, 1, 5, 4, -3, 3,
    -- filter=82 channel=35
    1, -2, 1, 3, -4, -6, 10, 7, -8,
    -- filter=82 channel=36
    -3, -1, -10, 0, -6, 0, 0, 5, 11,
    -- filter=82 channel=37
    11, -1, 7, 8, -7, -7, -2, -1, -3,
    -- filter=82 channel=38
    -4, 5, 13, -3, 1, 3, -1, -11, -11,
    -- filter=82 channel=39
    2, 2, 9, 5, 2, 5, 2, -2, 9,
    -- filter=82 channel=40
    4, 8, 0, -10, 5, -3, 9, -5, 3,
    -- filter=82 channel=41
    1, -5, 15, -11, -8, -2, -5, -11, -10,
    -- filter=82 channel=42
    -6, 4, -7, 0, 0, 2, 1, -5, -4,
    -- filter=82 channel=43
    13, 3, -3, -1, 6, 0, 0, 5, -7,
    -- filter=82 channel=44
    -9, 0, 2, 5, 6, 5, -9, 8, -1,
    -- filter=82 channel=45
    -4, -9, 5, -2, 3, -8, 1, -1, 7,
    -- filter=82 channel=46
    -2, 4, -3, -2, -1, 11, -2, 3, 0,
    -- filter=82 channel=47
    5, 4, -5, -4, 4, -9, -10, 9, 10,
    -- filter=82 channel=48
    -4, 10, -5, -8, 6, 10, 3, -11, 5,
    -- filter=82 channel=49
    -6, -3, -7, -4, 0, 5, 9, -2, 0,
    -- filter=82 channel=50
    -6, -2, -7, 8, 1, 0, 8, 6, 0,
    -- filter=82 channel=51
    -1, 6, -7, 3, -2, 1, -2, 0, 0,
    -- filter=82 channel=52
    -1, 9, 7, -3, -3, 0, -5, 6, 3,
    -- filter=82 channel=53
    -1, 0, -12, 0, -4, 5, -4, 3, 6,
    -- filter=82 channel=54
    6, 2, 7, -9, 2, 5, -4, 7, -2,
    -- filter=82 channel=55
    7, 4, 0, -3, 4, 1, -10, -6, -6,
    -- filter=82 channel=56
    -7, 3, 0, 8, 5, -7, 9, -5, 8,
    -- filter=82 channel=57
    8, 4, 3, 9, 3, -7, -2, -8, 4,
    -- filter=82 channel=58
    6, 10, 3, 8, -2, -3, -6, 9, 9,
    -- filter=82 channel=59
    -2, -8, 7, 6, -2, 4, 2, -3, -5,
    -- filter=82 channel=60
    8, 2, 20, -10, -8, 6, -12, -13, 6,
    -- filter=82 channel=61
    8, 9, -2, 9, -4, -8, 1, 4, -11,
    -- filter=82 channel=62
    -4, 1, -3, 2, -9, -1, 3, 0, 5,
    -- filter=82 channel=63
    -3, -8, -3, 1, 1, 7, -6, -9, -5,
    -- filter=83 channel=0
    2, 3, -6, -6, 3, -5, 3, 13, 3,
    -- filter=83 channel=1
    -1, 7, -10, -7, -13, 0, -5, -5, -8,
    -- filter=83 channel=2
    -5, 4, 5, 0, 0, 10, 11, 3, 14,
    -- filter=83 channel=3
    -12, 4, -2, -9, 0, 4, -8, -9, 0,
    -- filter=83 channel=4
    4, 5, -1, 9, -2, -8, 0, 13, -3,
    -- filter=83 channel=5
    5, -12, 6, 7, -12, -2, 4, -8, 0,
    -- filter=83 channel=6
    1, 6, 8, -6, -3, 8, 1, 13, 5,
    -- filter=83 channel=7
    3, 3, -7, 6, -13, -13, 2, 2, -8,
    -- filter=83 channel=8
    8, 1, -6, 6, -8, 2, 16, 15, 14,
    -- filter=83 channel=9
    -9, -12, 1, 0, -2, -9, 11, -7, 4,
    -- filter=83 channel=10
    -5, 6, 10, -5, 6, 13, 7, 0, -5,
    -- filter=83 channel=11
    6, -3, 2, 0, -2, -4, 2, 3, 6,
    -- filter=83 channel=12
    3, -6, -2, -4, -2, -1, 10, -1, -10,
    -- filter=83 channel=13
    6, -3, -14, 4, 6, -12, 13, 8, 12,
    -- filter=83 channel=14
    -8, -7, 0, 2, -7, -1, -4, 2, -4,
    -- filter=83 channel=15
    -1, -14, -13, 6, -1, -1, 15, 8, 2,
    -- filter=83 channel=16
    2, 0, -15, -2, -3, -3, 13, 8, 13,
    -- filter=83 channel=17
    8, -4, -6, 9, -6, 0, -1, 11, 9,
    -- filter=83 channel=18
    4, 7, -4, -3, 4, 13, 0, 11, 0,
    -- filter=83 channel=19
    3, -7, 0, 3, 5, 1, 4, -4, -8,
    -- filter=83 channel=20
    -14, 1, -9, 4, -4, -16, -12, -8, -3,
    -- filter=83 channel=21
    6, -5, 1, -7, -3, -4, 2, -6, -1,
    -- filter=83 channel=22
    10, 0, 7, -7, 0, 2, -10, 10, -9,
    -- filter=83 channel=23
    -5, 8, 2, 4, -6, 9, 3, 5, -6,
    -- filter=83 channel=24
    -1, -6, -12, 3, 0, -3, -1, 1, 0,
    -- filter=83 channel=25
    -10, 7, 2, 0, 4, -8, 11, 6, 3,
    -- filter=83 channel=26
    -12, 2, 4, -11, -13, 0, -2, -15, -15,
    -- filter=83 channel=27
    7, -3, -4, -3, -10, 3, 3, 14, 17,
    -- filter=83 channel=28
    1, 3, -7, 5, 9, 3, 10, 5, 1,
    -- filter=83 channel=29
    -7, -14, -6, -10, -9, -11, 13, 2, 16,
    -- filter=83 channel=30
    -12, -10, -18, -3, -23, -22, -15, -19, -8,
    -- filter=83 channel=31
    -1, 7, 1, 8, 8, 0, -2, -10, 7,
    -- filter=83 channel=32
    -8, 2, 10, 1, -1, -5, 4, -3, 1,
    -- filter=83 channel=33
    3, 8, 0, 6, 9, 9, 10, 1, 5,
    -- filter=83 channel=34
    4, 4, 6, -10, -12, 0, 2, 4, -1,
    -- filter=83 channel=35
    -1, -4, 12, -9, -5, 5, 4, 12, 12,
    -- filter=83 channel=36
    10, 9, -8, 4, 2, 0, -3, 0, -5,
    -- filter=83 channel=37
    -11, -12, 0, 0, 5, 4, -6, -11, -3,
    -- filter=83 channel=38
    -6, 5, -4, -10, -11, -2, 0, 5, 3,
    -- filter=83 channel=39
    0, 8, 4, 1, 2, -1, 1, 1, 1,
    -- filter=83 channel=40
    6, -9, -7, -7, 7, 6, 7, -10, -9,
    -- filter=83 channel=41
    3, -9, -10, -8, -8, 10, 9, 16, 14,
    -- filter=83 channel=42
    -10, 0, -8, 0, -1, 4, 4, 2, -5,
    -- filter=83 channel=43
    -7, -7, 0, -18, -9, -12, -9, -21, -7,
    -- filter=83 channel=44
    10, -12, -11, -1, 2, -3, -4, -6, -5,
    -- filter=83 channel=45
    -1, -2, -9, -2, -4, 0, 2, 9, -9,
    -- filter=83 channel=46
    -10, 0, -4, -5, -12, -16, -8, -12, -2,
    -- filter=83 channel=47
    7, 3, 2, -2, -8, 7, -9, -8, -6,
    -- filter=83 channel=48
    2, -11, -11, 3, -10, 0, 7, -1, 9,
    -- filter=83 channel=49
    -10, 0, -5, -5, 8, 11, -3, 1, 6,
    -- filter=83 channel=50
    -15, -11, -13, -10, -20, -21, 1, -2, -13,
    -- filter=83 channel=51
    -1, 5, 0, -2, 3, 10, 5, 11, 11,
    -- filter=83 channel=52
    9, 1, -10, 5, 6, 8, -3, 0, -5,
    -- filter=83 channel=53
    0, -2, -9, -5, -16, -5, -7, -14, -6,
    -- filter=83 channel=54
    -4, -15, 0, -1, -3, -9, -3, 7, -6,
    -- filter=83 channel=55
    -9, -9, -6, 7, 1, -5, -4, -6, -5,
    -- filter=83 channel=56
    1, 4, 6, -2, 5, -8, -8, -8, -9,
    -- filter=83 channel=57
    5, -4, 8, -1, -10, -5, -10, -7, 7,
    -- filter=83 channel=58
    0, 0, 10, 6, -7, -9, 9, -4, -9,
    -- filter=83 channel=59
    -4, -2, -4, -10, -4, -8, 4, 12, 8,
    -- filter=83 channel=60
    -9, -12, -8, 6, 6, 5, 20, 17, 24,
    -- filter=83 channel=61
    10, 6, -9, -7, 3, 3, 0, 3, 18,
    -- filter=83 channel=62
    6, -8, -2, 8, -1, 0, 8, 1, 1,
    -- filter=83 channel=63
    -7, -1, -2, 8, 0, -3, -1, -2, 4,
    -- filter=84 channel=0
    2, -3, -7, -5, -4, -10, -6, -6, -7,
    -- filter=84 channel=1
    0, -2, -7, -5, 0, -2, -2, 0, 14,
    -- filter=84 channel=2
    1, 3, -3, -1, 1, 10, 7, 2, 15,
    -- filter=84 channel=3
    2, 17, 14, 5, 6, 16, 10, 15, 15,
    -- filter=84 channel=4
    -13, -5, -3, -2, 0, -5, 6, 6, 5,
    -- filter=84 channel=5
    10, -1, 8, -5, 7, 3, -7, 12, 10,
    -- filter=84 channel=6
    -14, -4, -2, 8, -6, 0, -5, 7, 7,
    -- filter=84 channel=7
    0, 5, -4, 11, -4, -2, -1, 0, 10,
    -- filter=84 channel=8
    -3, -4, -20, -12, 2, 11, 2, 18, 4,
    -- filter=84 channel=9
    9, 17, 7, 8, 24, 20, 8, 10, 21,
    -- filter=84 channel=10
    -1, -7, 3, -10, -3, 5, -8, 5, 0,
    -- filter=84 channel=11
    -12, -5, -9, -13, -3, 5, -6, -3, 14,
    -- filter=84 channel=12
    10, 4, 1, 10, 9, 8, -1, 5, 4,
    -- filter=84 channel=13
    -10, -13, -2, -10, 3, -9, -5, 8, -4,
    -- filter=84 channel=14
    6, 5, -3, -3, 12, 3, 6, -1, 12,
    -- filter=84 channel=15
    -13, -10, 0, 9, 15, 13, -7, 18, 11,
    -- filter=84 channel=16
    -12, -4, -17, 2, -3, 16, 10, 13, 21,
    -- filter=84 channel=17
    -10, -9, -13, 2, 0, -4, -2, 15, 7,
    -- filter=84 channel=18
    -6, -6, -2, -12, -10, 0, -10, 4, -1,
    -- filter=84 channel=19
    5, 0, 1, 2, 15, 11, -4, 15, -1,
    -- filter=84 channel=20
    11, 10, -4, 6, 9, 0, -1, 5, 4,
    -- filter=84 channel=21
    8, 1, 3, 2, -10, 9, 2, -5, 5,
    -- filter=84 channel=22
    8, 0, 0, -5, 3, -7, 9, 5, 1,
    -- filter=84 channel=23
    -4, 1, -9, 0, -3, -5, 0, -8, 0,
    -- filter=84 channel=24
    -14, -8, -4, -8, -11, -8, -8, 3, -1,
    -- filter=84 channel=25
    0, -8, 6, -10, 11, 16, 3, 7, 11,
    -- filter=84 channel=26
    12, 2, 3, 14, 8, -3, 11, 9, 1,
    -- filter=84 channel=27
    -1, -5, -3, 3, 3, 6, -9, 6, 6,
    -- filter=84 channel=28
    -8, 0, -20, -7, 11, 6, 3, -2, 13,
    -- filter=84 channel=29
    0, -7, -18, 0, 10, -2, 0, 10, 15,
    -- filter=84 channel=30
    10, 25, -1, 11, 28, 19, 4, 21, 17,
    -- filter=84 channel=31
    -6, 6, -8, -5, -6, -2, 4, 3, -4,
    -- filter=84 channel=32
    2, 10, 14, 5, -3, 10, 10, 6, 14,
    -- filter=84 channel=33
    -8, -4, -8, -2, 7, 3, 8, 7, -7,
    -- filter=84 channel=34
    0, 6, 10, 4, -2, 12, 9, 13, 3,
    -- filter=84 channel=35
    0, -6, 10, 0, -1, 6, -1, 0, -1,
    -- filter=84 channel=36
    -2, 2, -7, -1, 2, -5, -6, 7, 0,
    -- filter=84 channel=37
    6, 11, 1, 10, 3, 9, 11, 18, 2,
    -- filter=84 channel=38
    -18, 1, -7, -13, -6, -7, 1, 19, 3,
    -- filter=84 channel=39
    -4, -1, -6, -4, -9, -2, 3, 4, 2,
    -- filter=84 channel=40
    -8, -1, 7, -3, 1, -5, 4, 3, -5,
    -- filter=84 channel=41
    0, -7, -15, -10, 17, 0, 14, 22, 18,
    -- filter=84 channel=42
    6, 0, -10, -4, 0, 2, 0, -4, 0,
    -- filter=84 channel=43
    -8, -5, -8, -9, -8, -13, -3, -1, -7,
    -- filter=84 channel=44
    7, 13, 17, -3, 16, 8, -3, 9, 18,
    -- filter=84 channel=45
    8, 5, 6, 8, -8, 9, -6, 9, 9,
    -- filter=84 channel=46
    1, -1, 4, 16, 12, 0, -1, 7, 7,
    -- filter=84 channel=47
    3, -3, 1, 2, 1, 0, 7, 5, -4,
    -- filter=84 channel=48
    -7, 3, -2, 5, 4, 2, 13, 0, 11,
    -- filter=84 channel=49
    6, 5, 4, 0, 9, 0, 6, 5, -1,
    -- filter=84 channel=50
    14, 7, -6, 0, 0, 9, -5, 5, 3,
    -- filter=84 channel=51
    -9, -15, -5, -9, -7, -4, -1, -7, -4,
    -- filter=84 channel=52
    10, -3, 7, 1, 6, -2, 7, 10, -2,
    -- filter=84 channel=53
    1, 11, 20, 11, 14, 12, 0, 16, 17,
    -- filter=84 channel=54
    10, 3, -4, 13, 11, 8, 3, 20, 21,
    -- filter=84 channel=55
    -3, -3, 2, 6, -6, 5, -5, -4, 9,
    -- filter=84 channel=56
    3, 11, 7, 6, 3, 4, 1, 13, 0,
    -- filter=84 channel=57
    -4, -9, 2, 9, -4, -9, 6, -1, -1,
    -- filter=84 channel=58
    9, 0, 6, 5, 6, 2, -2, -1, -4,
    -- filter=84 channel=59
    -5, 0, 8, 11, 6, 6, 3, 5, 5,
    -- filter=84 channel=60
    -6, -12, -14, -7, 8, -5, 1, 9, 13,
    -- filter=84 channel=61
    -7, -3, -18, -3, -11, -8, -3, 0, 9,
    -- filter=84 channel=62
    -12, -8, -3, -4, 9, 2, 0, 14, 2,
    -- filter=84 channel=63
    1, -5, 0, 8, 2, -4, -1, 10, -10,
    -- filter=85 channel=0
    -2, -8, -4, 2, 5, -9, -3, -4, -10,
    -- filter=85 channel=1
    5, 8, -9, 9, 8, 5, 9, 0, -8,
    -- filter=85 channel=2
    -5, 4, 5, -5, 6, 5, -5, -2, 4,
    -- filter=85 channel=3
    8, -9, -5, -9, 4, 0, -8, 6, -5,
    -- filter=85 channel=4
    9, 1, 4, 3, -7, -7, 8, 0, -8,
    -- filter=85 channel=5
    -9, 5, 10, 9, 0, -1, 2, 9, 1,
    -- filter=85 channel=6
    -8, 0, 0, -10, -5, -9, 4, -5, -1,
    -- filter=85 channel=7
    7, 8, 9, -9, -9, 5, 0, -4, 10,
    -- filter=85 channel=8
    -3, -5, -2, 0, 6, -3, -10, -4, -6,
    -- filter=85 channel=9
    0, 1, 6, -10, 6, -8, 4, 7, 3,
    -- filter=85 channel=10
    -3, 0, -4, 5, 8, 8, -5, -7, -1,
    -- filter=85 channel=11
    -5, 9, -2, -1, -9, 8, -3, -6, 6,
    -- filter=85 channel=12
    8, -2, -6, 4, 4, 10, 6, 9, -2,
    -- filter=85 channel=13
    6, 9, 6, 8, 5, 5, 3, -6, 2,
    -- filter=85 channel=14
    0, -6, -6, -7, 0, 10, -4, 0, 6,
    -- filter=85 channel=15
    4, 3, 2, -9, -1, 8, 0, 3, 0,
    -- filter=85 channel=16
    -3, 4, 6, -10, 0, 1, -10, -4, -6,
    -- filter=85 channel=17
    -1, 9, 5, -1, -8, -10, 7, -9, 0,
    -- filter=85 channel=18
    -10, -3, 0, -5, 5, 7, 9, 7, -2,
    -- filter=85 channel=19
    0, -3, 10, -5, -7, -7, -4, 4, 8,
    -- filter=85 channel=20
    -3, -3, -6, -10, 5, 7, 6, -9, 5,
    -- filter=85 channel=21
    -7, 4, -8, 0, -3, -4, 9, -2, -2,
    -- filter=85 channel=22
    -4, 5, -5, -7, 2, 5, 3, -6, 8,
    -- filter=85 channel=23
    7, 5, 9, 4, -1, -9, 4, -7, -1,
    -- filter=85 channel=24
    -2, 0, -10, -8, 9, -10, 9, -4, -4,
    -- filter=85 channel=25
    -4, -9, -8, -2, 5, -6, -7, -9, 0,
    -- filter=85 channel=26
    1, -10, 9, 0, -4, 0, 5, 1, -2,
    -- filter=85 channel=27
    -3, -7, -1, 4, -10, 9, 8, -2, 2,
    -- filter=85 channel=28
    7, 5, -5, 6, -1, -8, -5, -4, 0,
    -- filter=85 channel=29
    0, -1, -1, -7, 7, 5, 10, 7, -5,
    -- filter=85 channel=30
    -1, 9, 5, -3, 4, 7, 0, 7, -10,
    -- filter=85 channel=31
    4, -2, 7, 7, -3, -1, -3, -7, -6,
    -- filter=85 channel=32
    0, 9, -3, -3, 8, 0, -10, 6, 2,
    -- filter=85 channel=33
    -1, 7, 3, 0, 7, 4, 5, 6, 3,
    -- filter=85 channel=34
    0, -4, 7, -1, -5, 0, 0, 9, 0,
    -- filter=85 channel=35
    4, 2, -6, -8, 4, 4, 5, 5, -8,
    -- filter=85 channel=36
    4, -2, 0, -4, -2, -9, 6, -1, -5,
    -- filter=85 channel=37
    4, -1, 0, 2, -9, -4, -6, -7, -6,
    -- filter=85 channel=38
    6, -9, 0, -7, 0, 6, 9, 9, 4,
    -- filter=85 channel=39
    -1, 0, 5, 6, 2, -8, -5, -6, 1,
    -- filter=85 channel=40
    -3, 8, 6, 0, -2, 3, -1, 3, -8,
    -- filter=85 channel=41
    -10, 5, -6, -1, 8, -4, -9, -1, 5,
    -- filter=85 channel=42
    -9, -2, -5, 7, -6, 0, -9, -1, -7,
    -- filter=85 channel=43
    8, 5, 1, -3, -6, -10, -3, 1, -9,
    -- filter=85 channel=44
    -10, 8, -7, -1, 2, -1, -8, -2, 9,
    -- filter=85 channel=45
    3, -5, 6, -5, -4, 6, -3, 10, -3,
    -- filter=85 channel=46
    0, -10, -3, 2, -8, 5, -2, 7, 2,
    -- filter=85 channel=47
    0, 1, 1, 2, -7, 4, 3, 0, 8,
    -- filter=85 channel=48
    -7, 10, -1, -3, -9, -5, 10, -9, -7,
    -- filter=85 channel=49
    0, 3, -10, 3, 3, 2, -10, 7, 0,
    -- filter=85 channel=50
    -5, 7, 0, 4, -6, 2, -8, -4, -2,
    -- filter=85 channel=51
    0, 9, -5, -8, 9, -4, 2, -5, 3,
    -- filter=85 channel=52
    10, 8, 6, 0, -8, -8, -6, 3, 5,
    -- filter=85 channel=53
    -6, 9, 5, 1, 2, -4, -10, -4, 0,
    -- filter=85 channel=54
    0, -4, 3, 8, -7, -6, -7, 3, -7,
    -- filter=85 channel=55
    -4, -7, 0, -2, -7, 6, 2, 4, 2,
    -- filter=85 channel=56
    -4, 8, 2, 0, 8, 0, -7, 9, 9,
    -- filter=85 channel=57
    5, 3, -1, -6, -4, 8, -4, -7, -7,
    -- filter=85 channel=58
    3, -1, 6, -9, -7, 5, 1, -3, -4,
    -- filter=85 channel=59
    -10, -3, -10, 7, 7, -3, -1, -3, 6,
    -- filter=85 channel=60
    -1, -4, 0, 0, 3, 8, 1, 9, -3,
    -- filter=85 channel=61
    -6, -5, -1, 4, 1, -9, 8, -1, 1,
    -- filter=85 channel=62
    0, 10, -4, -6, -5, -5, -4, 0, 7,
    -- filter=85 channel=63
    1, 0, -6, 6, -6, -1, 1, -3, 3,
    -- filter=86 channel=0
    12, 7, -7, 6, 17, -8, 7, 4, 9,
    -- filter=86 channel=1
    -8, 9, 7, -7, 5, 2, -5, 9, 14,
    -- filter=86 channel=2
    -8, -3, -8, -20, 15, 4, -6, -6, 10,
    -- filter=86 channel=3
    -9, 0, 7, -2, 10, 0, -11, 3, 10,
    -- filter=86 channel=4
    -2, -2, 12, -12, -3, -8, -1, 8, 2,
    -- filter=86 channel=5
    0, 8, 5, 6, -7, 13, 0, 7, -2,
    -- filter=86 channel=6
    -9, 7, -2, -10, 11, -2, -8, -1, -11,
    -- filter=86 channel=7
    10, 9, 10, 10, 2, 15, 10, 9, 2,
    -- filter=86 channel=8
    -10, 9, -5, -23, 17, 5, -13, -3, -3,
    -- filter=86 channel=9
    0, 0, 17, -11, 4, 1, 5, 9, 9,
    -- filter=86 channel=10
    4, 1, -6, 9, 8, 4, 9, 0, 0,
    -- filter=86 channel=11
    -6, 10, 5, -16, 9, 0, -1, 4, 10,
    -- filter=86 channel=12
    0, 8, -5, -2, 2, 0, 2, 3, 3,
    -- filter=86 channel=13
    -4, 9, 0, -6, 5, -1, -14, -5, -8,
    -- filter=86 channel=14
    12, 6, 9, 0, 5, 16, -1, 16, 13,
    -- filter=86 channel=15
    0, 21, 1, -3, 18, -1, -5, 17, 2,
    -- filter=86 channel=16
    -8, -7, -8, -25, 14, 4, -24, 12, 0,
    -- filter=86 channel=17
    -4, 1, 10, 0, 7, 7, -10, 0, 9,
    -- filter=86 channel=18
    5, 6, 3, 2, -2, -13, 5, -8, -9,
    -- filter=86 channel=19
    -7, -3, 6, -5, -11, 18, -1, -12, 12,
    -- filter=86 channel=20
    10, 7, 0, 11, 6, -5, 14, -2, 5,
    -- filter=86 channel=21
    -3, 0, -9, -5, 4, -4, 8, -4, -1,
    -- filter=86 channel=22
    3, 4, 9, -2, 1, 0, 10, 0, 1,
    -- filter=86 channel=23
    6, -4, 3, 0, 7, -1, 10, -4, 2,
    -- filter=86 channel=24
    -12, 6, 0, -15, 2, 2, -9, 8, -4,
    -- filter=86 channel=25
    0, 10, -6, -1, 17, 14, -8, 4, 11,
    -- filter=86 channel=26
    2, 7, 16, 19, 18, 7, 4, 16, 11,
    -- filter=86 channel=27
    -3, 2, 0, 0, 3, 0, -5, 0, 11,
    -- filter=86 channel=28
    -10, 0, -10, -14, -14, 8, -13, 1, -6,
    -- filter=86 channel=29
    -20, 3, -12, -27, 7, 8, -18, 15, -1,
    -- filter=86 channel=30
    10, 20, 28, 29, 29, 35, 11, 27, 30,
    -- filter=86 channel=31
    1, -11, 8, -8, -5, 3, -6, -10, -5,
    -- filter=86 channel=32
    -3, 14, 13, 5, 18, 15, -5, 6, 14,
    -- filter=86 channel=33
    -5, 0, -8, -7, 4, 4, -2, -3, -1,
    -- filter=86 channel=34
    0, -1, 9, 13, 0, 3, 13, 10, -6,
    -- filter=86 channel=35
    -6, 14, -1, -2, 15, 0, 2, 22, -4,
    -- filter=86 channel=36
    9, 0, 4, 2, 7, -3, -7, -8, 3,
    -- filter=86 channel=37
    6, 8, 8, -12, 5, 4, -6, -7, -2,
    -- filter=86 channel=38
    -2, 16, 5, -11, 24, -5, -9, 2, 9,
    -- filter=86 channel=39
    -5, -4, 5, 7, 5, 4, 6, -10, 5,
    -- filter=86 channel=40
    4, 0, 9, 7, 5, -2, 5, 0, -4,
    -- filter=86 channel=41
    -13, 12, 0, -10, 16, 0, -16, 18, 0,
    -- filter=86 channel=42
    -4, 1, 1, -4, 3, 3, -7, -10, 0,
    -- filter=86 channel=43
    0, -8, 10, 2, 8, 14, 8, 9, 0,
    -- filter=86 channel=44
    10, 8, 4, 2, -4, 21, -1, 13, 12,
    -- filter=86 channel=45
    5, 6, -1, 3, 6, -7, -1, -3, 6,
    -- filter=86 channel=46
    0, 6, 11, 7, 20, 11, 0, 12, 8,
    -- filter=86 channel=47
    -7, 2, 3, 2, -1, -3, 4, 9, -7,
    -- filter=86 channel=48
    -1, 5, -9, -9, 4, -7, 0, 10, -10,
    -- filter=86 channel=49
    2, 18, -1, -13, -1, 5, -3, 8, -7,
    -- filter=86 channel=50
    5, 7, 8, 18, 0, 23, 15, 13, 24,
    -- filter=86 channel=51
    14, 3, -10, -5, 9, -11, 6, -8, -9,
    -- filter=86 channel=52
    -2, 8, 9, -9, 8, -6, -3, 1, 10,
    -- filter=86 channel=53
    3, 11, 8, 8, 12, 13, 1, 5, 19,
    -- filter=86 channel=54
    -8, -1, 14, -10, 8, 8, 0, 14, 16,
    -- filter=86 channel=55
    3, -9, -7, -4, 0, -8, -1, 8, 0,
    -- filter=86 channel=56
    10, 13, 8, 0, 10, 8, 7, 10, 9,
    -- filter=86 channel=57
    -2, 10, -4, -10, 1, -9, -10, -10, -9,
    -- filter=86 channel=58
    6, -3, -1, 6, 6, -8, -8, -7, -11,
    -- filter=86 channel=59
    -12, -1, -6, -15, 8, 0, 2, 11, -5,
    -- filter=86 channel=60
    -6, 12, 2, -11, 10, 10, -20, 9, -9,
    -- filter=86 channel=61
    -10, -5, 2, -14, 19, -3, -8, 10, 1,
    -- filter=86 channel=62
    -15, -9, 7, -15, 4, 5, -9, -1, 6,
    -- filter=86 channel=63
    8, 0, 6, 8, -4, -8, -5, 5, 9,
    -- filter=87 channel=0
    2, 1, 11, -9, 1, 14, -2, -6, 9,
    -- filter=87 channel=1
    -11, 3, -12, -18, 3, -3, -10, -10, 2,
    -- filter=87 channel=2
    -15, -10, -7, -8, -13, 4, -18, -12, 3,
    -- filter=87 channel=3
    -9, 5, 4, 3, 8, 15, -9, -5, 11,
    -- filter=87 channel=4
    10, 2, -1, -10, 5, 10, -1, -4, 9,
    -- filter=87 channel=5
    13, 9, 14, 14, 0, 16, -1, 14, 13,
    -- filter=87 channel=6
    -10, -4, -7, -10, -2, 0, 7, -4, 5,
    -- filter=87 channel=7
    -1, -1, 0, 1, 13, 7, 8, 6, 15,
    -- filter=87 channel=8
    2, 2, 1, 0, 10, 7, 2, 0, 12,
    -- filter=87 channel=9
    12, 20, 29, 17, 32, 24, -3, 21, 19,
    -- filter=87 channel=10
    8, -12, 0, -5, 3, -9, -5, 1, 1,
    -- filter=87 channel=11
    -12, -9, -8, -1, 2, 0, -8, 0, -6,
    -- filter=87 channel=12
    9, 1, 5, 5, 0, -2, 7, 2, 5,
    -- filter=87 channel=13
    -2, 1, 8, 8, 17, 5, -13, -2, 3,
    -- filter=87 channel=14
    11, 9, 15, 16, 7, 11, 2, 15, 3,
    -- filter=87 channel=15
    -5, -5, 1, -3, 16, 16, -4, 8, -3,
    -- filter=87 channel=16
    1, -8, -3, -9, 7, 10, -3, -10, -5,
    -- filter=87 channel=17
    -1, 5, -3, -9, -1, 0, -12, -3, -3,
    -- filter=87 channel=18
    9, -4, 3, 4, 14, 7, -3, 10, 3,
    -- filter=87 channel=19
    0, 10, 8, -11, -5, 5, 1, 0, -11,
    -- filter=87 channel=20
    11, 4, 17, 17, 25, 17, 7, 24, 14,
    -- filter=87 channel=21
    -8, 1, -7, -9, -8, 6, 7, 0, 6,
    -- filter=87 channel=22
    5, 9, -6, 9, 1, -5, 8, -2, -8,
    -- filter=87 channel=23
    -2, -12, -6, 3, -9, 10, -10, 4, 11,
    -- filter=87 channel=24
    6, 5, -9, -10, -6, 13, -3, 11, 0,
    -- filter=87 channel=25
    -19, -5, 0, -19, 0, 0, -17, -13, -9,
    -- filter=87 channel=26
    17, 18, 1, 1, 4, 13, 10, 19, 5,
    -- filter=87 channel=27
    -12, -11, -3, -11, -5, 5, -12, -5, 12,
    -- filter=87 channel=28
    0, 9, 4, -11, 14, 7, -12, 5, 7,
    -- filter=87 channel=29
    -11, 2, -8, -17, 6, 0, -5, -6, -8,
    -- filter=87 channel=30
    27, 38, 27, 32, 26, 25, 27, 28, 26,
    -- filter=87 channel=31
    -2, 1, -4, 8, -3, -9, 3, 4, 1,
    -- filter=87 channel=32
    11, 11, 14, 0, -7, 13, -3, 9, 19,
    -- filter=87 channel=33
    -1, 3, 4, -8, 6, 9, 10, 7, 3,
    -- filter=87 channel=34
    12, 17, 1, 1, 7, -1, 10, 9, 3,
    -- filter=87 channel=35
    -5, 0, 8, -13, -7, -7, -16, 1, 2,
    -- filter=87 channel=36
    7, -7, 4, -7, -11, -4, -6, 0, 2,
    -- filter=87 channel=37
    -3, 10, 1, 0, 3, 0, -8, 9, 0,
    -- filter=87 channel=38
    -1, -12, -5, -13, -12, -2, -12, -7, 0,
    -- filter=87 channel=39
    2, 4, -6, -4, 9, -3, -9, -6, -6,
    -- filter=87 channel=40
    6, 6, 10, -10, -8, 7, 4, 6, 3,
    -- filter=87 channel=41
    -12, -11, -2, -11, 0, 4, -14, 11, 11,
    -- filter=87 channel=42
    -10, -4, -5, -5, 4, 3, -2, 1, 8,
    -- filter=87 channel=43
    8, 6, -10, 5, 5, -11, -5, -1, 10,
    -- filter=87 channel=44
    6, 11, 18, 3, -9, -2, 11, 9, 0,
    -- filter=87 channel=45
    -5, -9, 6, 6, -10, 0, 3, 9, 5,
    -- filter=87 channel=46
    12, 4, 9, 15, 12, 12, 12, 4, 1,
    -- filter=87 channel=47
    -7, 7, -4, -10, 8, -5, -2, 0, 0,
    -- filter=87 channel=48
    -2, 4, 8, -11, 2, 14, 2, -5, 0,
    -- filter=87 channel=49
    2, -9, 11, -6, 3, -5, 5, 2, -6,
    -- filter=87 channel=50
    22, 23, 15, 23, 22, 11, 8, 5, 11,
    -- filter=87 channel=51
    12, -2, 3, -1, -3, -5, 11, 7, 3,
    -- filter=87 channel=52
    6, 9, -9, -9, -7, 6, 2, -5, 3,
    -- filter=87 channel=53
    15, 9, 24, 6, 9, 19, 17, 23, 22,
    -- filter=87 channel=54
    2, 29, 27, 15, 32, 30, 13, 20, 23,
    -- filter=87 channel=55
    -3, -8, -7, -1, -7, 9, -7, -10, 3,
    -- filter=87 channel=56
    8, 9, -5, -3, 10, -3, -3, 7, 14,
    -- filter=87 channel=57
    8, -6, 0, 2, 1, -5, 3, 2, 6,
    -- filter=87 channel=58
    6, 10, -2, 0, -7, 0, 10, 7, -10,
    -- filter=87 channel=59
    -8, 5, 5, -4, -6, 8, -5, 1, 11,
    -- filter=87 channel=60
    -11, -4, 7, 4, 20, 19, -7, 10, 2,
    -- filter=87 channel=61
    10, 1, -10, -14, -2, 4, -15, 4, 14,
    -- filter=87 channel=62
    1, 4, -6, -7, 9, 0, -14, 6, -6,
    -- filter=87 channel=63
    2, 5, 3, -5, -3, -8, -8, 0, -6,
    -- filter=88 channel=0
    -5, 10, 17, 13, 17, 18, 11, 8, 0,
    -- filter=88 channel=1
    -15, -9, -2, -7, -22, -2, -11, -23, 0,
    -- filter=88 channel=2
    -20, -13, -19, -10, -13, -9, -15, -13, -16,
    -- filter=88 channel=3
    -16, -7, -16, -4, -16, 0, -2, -9, -5,
    -- filter=88 channel=4
    9, 1, 13, 9, 20, 8, 16, 6, 8,
    -- filter=88 channel=5
    -4, 5, -1, -10, 2, 9, -10, 4, 1,
    -- filter=88 channel=6
    0, 4, 6, 4, 2, -3, 12, 0, 7,
    -- filter=88 channel=7
    -1, 7, 10, -4, -5, 9, 8, 6, 14,
    -- filter=88 channel=8
    -12, 2, 0, 12, 10, 16, -2, 19, 6,
    -- filter=88 channel=9
    1, 3, -13, 10, -10, -15, 2, 2, 2,
    -- filter=88 channel=10
    11, 10, 9, -3, 2, 10, 3, 9, 5,
    -- filter=88 channel=11
    -4, -6, -3, -6, 9, 6, 6, -2, 11,
    -- filter=88 channel=12
    -1, 11, 11, -5, 9, 9, 0, 7, -1,
    -- filter=88 channel=13
    -4, 11, 2, 14, 10, 11, -1, 16, 14,
    -- filter=88 channel=14
    10, 4, 9, 7, 5, 11, 9, 11, 15,
    -- filter=88 channel=15
    -7, 4, 15, 1, 19, 2, 11, 17, 14,
    -- filter=88 channel=16
    -4, -12, 0, -6, 1, 4, -4, 7, 3,
    -- filter=88 channel=17
    3, 5, 11, -1, 9, 0, -4, -2, -2,
    -- filter=88 channel=18
    17, 26, 26, 12, 28, 27, 22, 27, 21,
    -- filter=88 channel=19
    -3, -12, 0, -6, -8, -5, 1, 2, 2,
    -- filter=88 channel=20
    -6, 12, 0, -4, 14, 11, 8, 13, 12,
    -- filter=88 channel=21
    0, 0, 2, -2, 11, 4, 5, 11, 3,
    -- filter=88 channel=22
    -5, -1, 8, -6, -7, -1, -10, -6, 0,
    -- filter=88 channel=23
    0, -2, 1, -2, 1, 10, 0, 0, 13,
    -- filter=88 channel=24
    6, 4, 8, 12, 12, -4, 9, 1, 13,
    -- filter=88 channel=25
    -29, -25, -12, -9, -31, -8, -12, -29, -6,
    -- filter=88 channel=26
    -10, 1, 1, 4, 6, 5, 0, 2, 0,
    -- filter=88 channel=27
    -13, -13, 0, -11, -1, -13, -18, -10, -8,
    -- filter=88 channel=28
    4, -3, -1, 15, 10, 4, 11, 13, 17,
    -- filter=88 channel=29
    -18, 5, 2, -2, 5, 13, 5, 0, 12,
    -- filter=88 channel=30
    3, -7, 19, 1, -3, 5, 14, 8, 6,
    -- filter=88 channel=31
    9, 9, 12, 3, 12, -4, 9, -5, 0,
    -- filter=88 channel=32
    -5, -14, -9, -12, -21, -7, 1, -18, 0,
    -- filter=88 channel=33
    6, 6, 5, 5, -3, -7, 7, 10, -6,
    -- filter=88 channel=34
    5, -1, -1, 0, 0, 8, 4, 0, -1,
    -- filter=88 channel=35
    -19, -12, 5, -4, -19, -9, -7, -20, -14,
    -- filter=88 channel=36
    1, -1, 0, -7, 6, 1, -6, 2, 10,
    -- filter=88 channel=37
    -4, -14, -6, -14, -5, -15, -2, -15, 1,
    -- filter=88 channel=38
    -19, -2, -3, -7, 0, -5, -1, 2, 1,
    -- filter=88 channel=39
    9, 5, 1, -10, 6, -2, 9, 4, -5,
    -- filter=88 channel=40
    1, -7, 0, -8, -3, -1, 1, -11, -5,
    -- filter=88 channel=41
    -19, -11, -4, 0, -10, 12, -3, -5, 7,
    -- filter=88 channel=42
    -9, 3, 4, -9, -3, -9, 3, -8, 10,
    -- filter=88 channel=43
    0, -15, -22, -13, -26, -16, -13, -22, -14,
    -- filter=88 channel=44
    -13, -15, 4, -2, -17, -1, 2, -16, -12,
    -- filter=88 channel=45
    -3, -9, -7, -7, 1, 3, 9, -1, -4,
    -- filter=88 channel=46
    2, 12, 14, 10, 7, 10, 0, 0, 6,
    -- filter=88 channel=47
    -9, 8, 3, -7, 4, 4, -1, -9, 9,
    -- filter=88 channel=48
    -6, 8, 2, -10, 7, 7, 1, 5, 0,
    -- filter=88 channel=49
    13, 0, 15, 0, 1, 11, -4, 13, 11,
    -- filter=88 channel=50
    8, 3, 3, 3, -7, -1, 4, 4, 14,
    -- filter=88 channel=51
    3, 24, 20, 20, 10, 26, 13, 10, 16,
    -- filter=88 channel=52
    8, -6, -2, 3, 8, 7, 5, 4, 0,
    -- filter=88 channel=53
    -4, -9, 11, -4, -12, -7, -5, 3, 13,
    -- filter=88 channel=54
    -2, -6, -7, 0, -10, -3, -12, -8, -1,
    -- filter=88 channel=55
    -9, -7, -8, -10, 1, 10, 6, -5, 5,
    -- filter=88 channel=56
    -1, 4, 9, -7, -1, 7, 12, 11, 7,
    -- filter=88 channel=57
    -7, -5, 2, 0, -1, 8, 7, 0, -8,
    -- filter=88 channel=58
    8, 17, 0, 10, 8, 5, 9, 6, 8,
    -- filter=88 channel=59
    -2, -15, -15, -22, -20, -15, -14, -2, 0,
    -- filter=88 channel=60
    -2, 2, 6, 10, 21, 19, 11, 8, 14,
    -- filter=88 channel=61
    -9, -5, 0, 9, 2, 20, -5, 0, 4,
    -- filter=88 channel=62
    1, -12, -6, 1, -13, -8, 2, -5, -7,
    -- filter=88 channel=63
    -4, -5, 8, 6, 8, 0, -6, -1, 9,
    -- filter=89 channel=0
    -9, -2, -5, -3, 3, 2, 1, 3, 0,
    -- filter=89 channel=1
    -10, -15, 0, -7, 4, 0, 7, 10, 5,
    -- filter=89 channel=2
    11, 0, -10, 1, -11, -17, -6, -3, -22,
    -- filter=89 channel=3
    13, 2, -4, 12, 17, 1, 9, 5, 0,
    -- filter=89 channel=4
    6, 3, -3, -1, 9, 11, -9, 9, -1,
    -- filter=89 channel=5
    7, 13, -3, 5, 6, 8, -9, -4, 2,
    -- filter=89 channel=6
    0, 13, -11, -1, -1, -2, 6, -4, -6,
    -- filter=89 channel=7
    5, 0, -8, 2, -3, -4, -9, 0, -7,
    -- filter=89 channel=8
    22, 23, 2, 11, 16, 8, 3, 2, -24,
    -- filter=89 channel=9
    9, 3, -10, 0, 9, -6, -6, 2, -17,
    -- filter=89 channel=10
    -16, -4, -6, -10, -6, 3, 2, -13, 3,
    -- filter=89 channel=11
    -2, 8, 9, 7, 8, 11, 4, 8, -15,
    -- filter=89 channel=12
    10, -2, -3, 2, -3, -2, -5, -6, 4,
    -- filter=89 channel=13
    1, 7, -11, 12, 6, 11, 12, 13, -17,
    -- filter=89 channel=14
    6, 1, 0, -6, -2, -1, -4, -10, 7,
    -- filter=89 channel=15
    23, 25, 5, 18, 23, -10, -4, 0, -23,
    -- filter=89 channel=16
    10, 23, 5, 30, 23, -8, 4, -10, -25,
    -- filter=89 channel=17
    17, 8, 3, 15, 14, 0, 6, 12, -6,
    -- filter=89 channel=18
    9, 12, 8, 12, 16, 9, -1, 8, -5,
    -- filter=89 channel=19
    -7, -4, 7, -3, -2, -8, 8, 2, 6,
    -- filter=89 channel=20
    -11, -7, -1, -1, -10, -2, -4, 0, -1,
    -- filter=89 channel=21
    7, 9, 1, -1, -9, 1, 7, 3, -5,
    -- filter=89 channel=22
    -7, 0, -5, -9, 4, 2, -3, 5, -6,
    -- filter=89 channel=23
    0, -1, -6, -2, 1, -3, -5, 0, -5,
    -- filter=89 channel=24
    6, 11, 7, 8, 17, 2, 8, 9, -10,
    -- filter=89 channel=25
    0, -11, -2, 4, -14, -20, 1, -13, -30,
    -- filter=89 channel=26
    -9, 1, -2, -10, -6, -5, 0, -15, -6,
    -- filter=89 channel=27
    -4, -1, -14, -2, -2, -16, 1, 2, -19,
    -- filter=89 channel=28
    15, 17, 11, 1, 19, 5, -7, 7, -15,
    -- filter=89 channel=29
    28, 32, 5, 34, 33, -2, 11, -2, -36,
    -- filter=89 channel=30
    -12, -22, 3, -20, -13, 0, -2, 6, -3,
    -- filter=89 channel=31
    -3, -2, -3, 4, 6, -2, 5, 10, 9,
    -- filter=89 channel=32
    -4, -18, -8, -10, -11, -6, -2, -11, -1,
    -- filter=89 channel=33
    -8, -2, -1, 5, -5, -1, 1, -1, 1,
    -- filter=89 channel=34
    3, 10, -10, 1, -6, -2, -9, 7, 3,
    -- filter=89 channel=35
    -8, -6, -10, -16, -21, -11, -19, -19, -16,
    -- filter=89 channel=36
    0, 0, 2, 0, -8, 3, -3, -5, -2,
    -- filter=89 channel=37
    5, 13, -8, 16, 9, -8, 1, 9, -14,
    -- filter=89 channel=38
    9, -2, -2, 12, 15, -2, 10, -5, -20,
    -- filter=89 channel=39
    11, -5, -9, 4, 0, 8, -4, 6, 0,
    -- filter=89 channel=40
    -3, -7, 0, 7, 1, -6, 7, -6, 4,
    -- filter=89 channel=41
    11, 27, -10, 9, 17, -5, -11, -18, -34,
    -- filter=89 channel=42
    -7, 1, 0, 8, -2, -6, -6, -8, 1,
    -- filter=89 channel=43
    -8, -27, -16, 2, -9, -1, 6, -12, 4,
    -- filter=89 channel=44
    -11, 1, 6, -17, -7, 2, -10, -7, 2,
    -- filter=89 channel=45
    2, 3, 9, 2, 7, 0, 7, -2, 8,
    -- filter=89 channel=46
    11, -6, -8, 1, -3, -4, -2, -7, -6,
    -- filter=89 channel=47
    1, -1, -1, -10, 9, -1, 0, 10, -3,
    -- filter=89 channel=48
    5, 13, 5, 5, 14, -14, -11, -13, -13,
    -- filter=89 channel=49
    11, -1, 3, 2, -9, -11, 0, -7, -3,
    -- filter=89 channel=50
    1, -14, -2, -11, -15, -3, 4, 12, 0,
    -- filter=89 channel=51
    -9, 5, -9, -5, 3, -3, 4, 12, 0,
    -- filter=89 channel=52
    4, -7, 4, 4, 8, 5, 6, 2, 7,
    -- filter=89 channel=53
    -14, -23, -1, -17, -5, -5, -4, 0, 2,
    -- filter=89 channel=54
    0, 13, 3, -6, -1, -4, -8, -1, -14,
    -- filter=89 channel=55
    -7, 0, 8, 10, -2, 6, -6, 9, 0,
    -- filter=89 channel=56
    3, -2, 4, -10, -7, 4, -5, 5, 0,
    -- filter=89 channel=57
    -9, -8, -9, 0, -1, 8, -2, -3, -6,
    -- filter=89 channel=58
    -6, 5, -2, 0, 3, 8, 9, 11, -4,
    -- filter=89 channel=59
    22, 13, -9, 11, -2, -8, 9, -14, -26,
    -- filter=89 channel=60
    15, 26, 5, 31, 36, -2, 8, -2, -17,
    -- filter=89 channel=61
    4, 0, 1, 0, 25, -3, -5, 7, -17,
    -- filter=89 channel=62
    9, 20, -3, 3, 11, -4, 4, 11, -14,
    -- filter=89 channel=63
    9, -9, 10, -9, 10, 2, -8, 3, -9,
    -- filter=90 channel=0
    14, 11, 1, -5, 17, 16, 8, -2, 18,
    -- filter=90 channel=1
    -4, -14, 3, -12, -23, -12, -14, -21, -10,
    -- filter=90 channel=2
    -17, -24, 0, -29, -26, -11, -17, -14, -8,
    -- filter=90 channel=3
    -9, -19, 8, -25, -4, -7, -17, -5, 0,
    -- filter=90 channel=4
    7, 19, 11, 0, 1, 19, -4, 9, 4,
    -- filter=90 channel=5
    -11, -5, 10, -1, 0, -7, 6, 1, 9,
    -- filter=90 channel=6
    -2, 12, 15, 3, 9, 6, 10, -2, 0,
    -- filter=90 channel=7
    1, 0, 7, 14, 7, 15, 8, -2, 12,
    -- filter=90 channel=8
    2, 6, 14, -2, -1, 6, -1, 0, 18,
    -- filter=90 channel=9
    7, 4, 3, -8, 4, 5, 6, 0, -3,
    -- filter=90 channel=10
    6, 13, 4, 14, 16, 16, 11, -1, 5,
    -- filter=90 channel=11
    -7, -9, 13, 0, -8, 10, -2, -10, -4,
    -- filter=90 channel=12
    -2, 5, 0, -1, -1, 6, -4, 2, -9,
    -- filter=90 channel=13
    15, 19, 17, 9, 18, 8, -2, 2, 10,
    -- filter=90 channel=14
    11, 11, 1, 12, 14, 3, -5, 7, 13,
    -- filter=90 channel=15
    2, 3, 27, 8, 13, 24, 8, -2, 21,
    -- filter=90 channel=16
    -5, -8, 14, -19, -10, 9, -9, -5, 0,
    -- filter=90 channel=17
    9, 1, 5, -6, -5, 11, 0, 8, 5,
    -- filter=90 channel=18
    14, 19, 14, 23, 21, 29, 22, 30, 14,
    -- filter=90 channel=19
    2, 0, 5, 1, -10, -3, -9, -5, -11,
    -- filter=90 channel=20
    16, 0, 15, -2, 3, 16, -1, 2, 19,
    -- filter=90 channel=21
    -3, -3, -3, 6, 3, 5, -2, -6, -7,
    -- filter=90 channel=22
    6, -5, 8, 5, -2, 4, 6, 2, -9,
    -- filter=90 channel=23
    13, 10, 1, -6, 12, -2, 0, 4, -1,
    -- filter=90 channel=24
    14, 4, 16, -4, -3, 14, 2, 6, 5,
    -- filter=90 channel=25
    -29, -25, -4, -34, -38, -4, -18, -26, -13,
    -- filter=90 channel=26
    6, 0, 7, 2, 8, 10, -2, 2, 22,
    -- filter=90 channel=27
    -20, -5, 1, -6, -23, -10, -19, -9, 3,
    -- filter=90 channel=28
    0, 10, 1, 9, -2, 3, -3, -4, 17,
    -- filter=90 channel=29
    -10, 2, 12, -7, 7, 15, -15, -4, 25,
    -- filter=90 channel=30
    9, 16, 28, 16, 14, 23, 6, 10, 27,
    -- filter=90 channel=31
    0, 2, 10, 7, -6, 8, 1, 3, 10,
    -- filter=90 channel=32
    -4, -12, -11, -10, -7, -16, -16, -16, -15,
    -- filter=90 channel=33
    4, -6, 3, 9, 2, 9, -5, 6, 3,
    -- filter=90 channel=34
    10, 8, 14, 8, 4, 9, 7, 2, 9,
    -- filter=90 channel=35
    -14, -16, -13, -18, -21, -14, -18, -13, 1,
    -- filter=90 channel=36
    0, 6, 9, 11, 7, -3, 7, 9, 8,
    -- filter=90 channel=37
    -10, -5, 1, -10, -9, 4, 0, -7, -14,
    -- filter=90 channel=38
    1, -15, -4, -24, -11, -5, -10, -3, 8,
    -- filter=90 channel=39
    0, 5, 9, 7, 9, 3, -9, -3, -9,
    -- filter=90 channel=40
    0, 2, 2, -7, 1, -3, 3, -7, 4,
    -- filter=90 channel=41
    -2, 2, 14, -15, -8, 0, -14, -6, 7,
    -- filter=90 channel=42
    -8, -7, -2, -3, -1, 5, -8, 4, 2,
    -- filter=90 channel=43
    3, -1, 16, 8, 8, 15, 2, 14, 9,
    -- filter=90 channel=44
    -4, -15, 0, 1, -15, 4, -15, -5, -12,
    -- filter=90 channel=45
    -10, 9, -10, -6, 0, -9, 3, -7, 2,
    -- filter=90 channel=46
    12, 2, 10, 0, 18, 8, 5, 0, 5,
    -- filter=90 channel=47
    -1, 9, 7, -7, 0, -2, 0, 10, -9,
    -- filter=90 channel=48
    -7, -5, 1, 1, 2, 2, 8, 4, 15,
    -- filter=90 channel=49
    -2, 17, 13, 13, 7, 2, 18, 20, 19,
    -- filter=90 channel=50
    13, 12, 19, 7, 9, 13, 6, 20, 6,
    -- filter=90 channel=51
    18, 9, 6, 11, 18, 21, 15, 22, 22,
    -- filter=90 channel=52
    -7, -4, -8, 7, -1, 4, -3, 8, -3,
    -- filter=90 channel=53
    -1, 0, 5, -6, -7, 5, 11, 1, 10,
    -- filter=90 channel=54
    -1, -8, -1, -11, -14, -11, -11, -17, -15,
    -- filter=90 channel=55
    -7, 2, 0, -10, 4, -4, -10, 3, 10,
    -- filter=90 channel=56
    0, 6, 5, 3, -3, 16, 10, 9, 7,
    -- filter=90 channel=57
    9, 0, -1, -8, -1, 5, -6, -4, 6,
    -- filter=90 channel=58
    -2, 0, 7, 4, -2, -2, 0, 15, 15,
    -- filter=90 channel=59
    -24, -17, 0, -9, -13, 8, -18, -2, 4,
    -- filter=90 channel=60
    8, 4, 23, 4, 13, 10, -13, -1, 23,
    -- filter=90 channel=61
    6, 8, 4, -3, 13, 10, -7, 3, 6,
    -- filter=90 channel=62
    -3, -16, 2, -10, -17, -3, -4, -15, -8,
    -- filter=90 channel=63
    4, 3, 2, 8, 7, 0, -8, -5, -3,
    -- filter=91 channel=0
    -14, -1, -19, 6, 0, 0, 9, 1, -8,
    -- filter=91 channel=1
    -7, -3, -3, -4, -9, 15, -3, 17, 5,
    -- filter=91 channel=2
    -4, 4, 0, -6, 19, 19, 5, 13, 18,
    -- filter=91 channel=3
    6, 9, 9, 6, 13, 3, 12, 11, 9,
    -- filter=91 channel=4
    3, 0, -1, -2, 2, -4, -11, 1, 0,
    -- filter=91 channel=5
    -7, 3, 6, 0, 8, 18, 5, -5, -3,
    -- filter=91 channel=6
    -5, -10, -8, -2, 10, 2, 7, -5, -5,
    -- filter=91 channel=7
    0, -8, 9, 6, 5, 0, 1, 4, 3,
    -- filter=91 channel=8
    -15, -19, -18, 2, 0, 14, 7, 17, 14,
    -- filter=91 channel=9
    -1, 10, -5, 0, 10, 15, 3, 7, 0,
    -- filter=91 channel=10
    6, -1, -4, -7, -17, 0, -4, 0, -10,
    -- filter=91 channel=11
    -8, -1, -16, 5, -8, 6, 2, 15, 10,
    -- filter=91 channel=12
    8, 8, 0, 3, 5, -3, -5, -5, 7,
    -- filter=91 channel=13
    0, -11, -11, 9, 7, 5, 0, 23, 11,
    -- filter=91 channel=14
    -7, -4, -10, -8, -8, -2, -8, -4, 11,
    -- filter=91 channel=15
    -6, 2, -16, 15, 17, 3, 0, 23, 6,
    -- filter=91 channel=16
    -5, -19, -12, -6, 14, 23, -4, 28, 18,
    -- filter=91 channel=17
    -6, 0, -13, -6, 6, 12, 9, 15, 6,
    -- filter=91 channel=18
    3, 6, -8, 6, 2, -7, 10, -6, -11,
    -- filter=91 channel=19
    0, 9, -5, 2, 13, 13, 7, 10, 6,
    -- filter=91 channel=20
    -11, -4, 0, -2, -2, -7, 5, -3, -6,
    -- filter=91 channel=21
    0, 0, 5, 4, 10, 4, 0, 0, -7,
    -- filter=91 channel=22
    0, 0, 2, -7, -9, 9, 2, -9, 2,
    -- filter=91 channel=23
    -10, -16, 5, 2, -15, 0, 7, -2, -5,
    -- filter=91 channel=24
    -10, -4, -1, 0, -4, 4, -11, 6, 1,
    -- filter=91 channel=25
    -3, -8, 2, 5, 8, 8, 0, 20, 26,
    -- filter=91 channel=26
    1, -4, 2, -1, 7, 6, 9, 10, 0,
    -- filter=91 channel=27
    -15, -2, -16, 8, 3, -1, 10, -1, 19,
    -- filter=91 channel=28
    -4, 0, -1, 6, 3, 18, -7, 3, 10,
    -- filter=91 channel=29
    -18, -14, -22, 19, 10, 17, 18, 33, 27,
    -- filter=91 channel=30
    7, 1, 2, -4, -12, -12, -7, 0, -1,
    -- filter=91 channel=31
    0, 1, 3, -3, 0, 7, 0, 3, 8,
    -- filter=91 channel=32
    -6, -4, -3, -3, 3, 0, 2, -9, -2,
    -- filter=91 channel=33
    7, -8, 3, 7, -5, -6, 5, -5, 0,
    -- filter=91 channel=34
    -9, 10, -2, 7, -1, 8, -5, 0, 5,
    -- filter=91 channel=35
    -5, 0, -9, -5, -4, 1, -14, -7, 4,
    -- filter=91 channel=36
    -8, 6, 1, 0, 2, 7, 2, 1, 0,
    -- filter=91 channel=37
    -7, -11, 3, -6, 2, -5, 2, 5, 14,
    -- filter=91 channel=38
    -19, -14, -21, -12, 8, -5, 0, 16, 25,
    -- filter=91 channel=39
    8, 0, -9, -6, -1, 0, -4, 5, 0,
    -- filter=91 channel=40
    -10, -8, 9, 6, 0, -2, 7, -8, 4,
    -- filter=91 channel=41
    1, -5, -20, -5, 21, 19, 0, 22, 24,
    -- filter=91 channel=42
    -1, 10, -6, -5, -4, -9, 0, -6, -5,
    -- filter=91 channel=43
    0, -16, 0, 3, -5, -4, 14, 13, 4,
    -- filter=91 channel=44
    7, 10, 3, -9, 1, 1, 5, 1, 9,
    -- filter=91 channel=45
    -6, -7, 0, 7, 0, 6, -6, 9, -10,
    -- filter=91 channel=46
    -10, 4, 1, 1, 10, -6, 4, 5, -9,
    -- filter=91 channel=47
    5, 0, -8, -1, -1, 7, -3, 4, -4,
    -- filter=91 channel=48
    -13, 5, 0, 2, 15, -3, -2, 16, 1,
    -- filter=91 channel=49
    9, -3, 3, -6, -5, 13, -4, -14, -1,
    -- filter=91 channel=50
    8, 5, -12, -9, -16, -2, 0, 1, -1,
    -- filter=91 channel=51
    -4, -6, -3, -1, -13, -8, -2, -10, -9,
    -- filter=91 channel=52
    -5, -7, 0, -4, -10, -4, 3, -4, 6,
    -- filter=91 channel=53
    -7, -6, -9, -3, -15, -3, 0, -9, -1,
    -- filter=91 channel=54
    -12, -1, -9, -8, 17, 7, -8, 12, 4,
    -- filter=91 channel=55
    3, 2, -6, -3, -4, -8, -9, -4, -8,
    -- filter=91 channel=56
    -4, -8, 5, -5, 1, 9, 0, -6, -10,
    -- filter=91 channel=57
    10, -1, 2, 9, -9, -1, 9, 0, 4,
    -- filter=91 channel=58
    2, 3, 7, -5, 1, 0, 8, 3, 7,
    -- filter=91 channel=59
    3, -1, -12, 9, -2, 15, -1, 7, 20,
    -- filter=91 channel=60
    -20, -9, -17, 10, 5, 10, 9, 18, 29,
    -- filter=91 channel=61
    -20, -17, -23, -13, -3, -11, 7, -5, 19,
    -- filter=91 channel=62
    4, 4, 3, 3, 15, 7, -3, 11, 12,
    -- filter=91 channel=63
    -8, -9, -8, 3, 4, 10, -5, -10, -4,
    -- filter=92 channel=0
    -7, -6, 0, -13, -6, 11, -6, -3, 13,
    -- filter=92 channel=1
    -3, 8, 10, -8, -3, -1, 3, 2, -12,
    -- filter=92 channel=2
    4, -1, 4, -7, -17, 3, -3, -1, 7,
    -- filter=92 channel=3
    2, -1, 4, -6, -3, 4, 9, 5, -1,
    -- filter=92 channel=4
    -7, 3, -3, -1, -2, -1, 2, 3, 0,
    -- filter=92 channel=5
    -4, 6, 13, 6, -7, -7, 9, -1, 0,
    -- filter=92 channel=6
    -8, 0, 0, -7, -7, -3, -1, -2, 0,
    -- filter=92 channel=7
    11, -4, 1, 3, -2, 4, 10, 0, -5,
    -- filter=92 channel=8
    -2, 8, 16, -4, -14, 4, 0, -6, -2,
    -- filter=92 channel=9
    3, -1, -8, -1, -3, 9, 5, 3, -8,
    -- filter=92 channel=10
    -8, -7, 11, 5, -6, 4, -4, -10, -3,
    -- filter=92 channel=11
    3, 0, 9, -3, 2, 12, 1, -9, 8,
    -- filter=92 channel=12
    2, -1, -6, 1, 8, 1, -5, 0, 3,
    -- filter=92 channel=13
    1, 13, 14, 5, 8, 12, -16, -13, 13,
    -- filter=92 channel=14
    2, 3, 8, 2, -2, 12, -3, 1, 8,
    -- filter=92 channel=15
    8, -2, 20, -5, -6, 17, 7, -6, 12,
    -- filter=92 channel=16
    -6, 5, 13, -6, -20, 9, 11, -18, -7,
    -- filter=92 channel=17
    2, 6, -3, -9, -17, 7, 6, -10, -8,
    -- filter=92 channel=18
    9, 3, -6, -6, 9, 5, 7, 4, -3,
    -- filter=92 channel=19
    1, 0, -4, 13, 0, -6, 8, -2, -14,
    -- filter=92 channel=20
    1, 1, 10, 2, -1, 15, -7, 11, -1,
    -- filter=92 channel=21
    4, -8, 0, 10, 1, 3, -3, 1, -7,
    -- filter=92 channel=22
    7, 1, 4, 8, 0, 2, -3, -9, 0,
    -- filter=92 channel=23
    2, -3, 1, 0, -11, 8, -9, 3, 8,
    -- filter=92 channel=24
    3, 0, -3, 5, -8, 2, 5, 5, 6,
    -- filter=92 channel=25
    -8, 5, 16, 3, -9, -5, -7, -2, -8,
    -- filter=92 channel=26
    5, -1, 14, 0, 8, 17, -10, 13, 3,
    -- filter=92 channel=27
    -7, -1, 17, 0, -16, 4, 11, -15, -11,
    -- filter=92 channel=28
    -11, -10, 14, -6, -5, -6, 12, -9, -14,
    -- filter=92 channel=29
    1, -1, 24, -16, -20, 16, -13, -7, 0,
    -- filter=92 channel=30
    8, 1, 3, 29, 10, 15, 11, 3, 0,
    -- filter=92 channel=31
    0, -4, 4, 2, 9, 9, -7, -3, 9,
    -- filter=92 channel=32
    4, -3, 3, 5, -7, -3, -2, 3, -9,
    -- filter=92 channel=33
    7, -1, -7, 1, 6, -6, 6, 8, -2,
    -- filter=92 channel=34
    -4, -1, 1, 6, 7, 0, -3, -2, 3,
    -- filter=92 channel=35
    -3, 0, 17, -10, -9, 11, -3, 0, -6,
    -- filter=92 channel=36
    -7, -3, -1, 0, -9, 6, -10, 3, 8,
    -- filter=92 channel=37
    -3, 11, -4, 1, 3, 13, -4, -2, 11,
    -- filter=92 channel=38
    6, 4, 4, -6, -1, 2, -3, -9, 9,
    -- filter=92 channel=39
    -9, -5, 2, -2, 7, -5, 4, 6, 0,
    -- filter=92 channel=40
    6, -5, 3, -4, 7, 0, -1, -7, -4,
    -- filter=92 channel=41
    -4, -9, 21, -2, -4, 21, -1, -4, 4,
    -- filter=92 channel=42
    -2, 0, 0, 3, 4, 8, 0, 5, -5,
    -- filter=92 channel=43
    0, 13, 5, 8, 22, 19, 0, 0, 12,
    -- filter=92 channel=44
    -3, 4, 1, 13, 10, 1, 7, -1, 1,
    -- filter=92 channel=45
    4, 10, 7, -7, -7, -1, -8, -5, 9,
    -- filter=92 channel=46
    3, 6, -1, -2, 3, 10, 5, -6, 7,
    -- filter=92 channel=47
    3, -8, -2, 5, 2, 10, 9, -8, 5,
    -- filter=92 channel=48
    5, -7, 13, 5, 1, 10, 2, -12, 2,
    -- filter=92 channel=49
    4, 0, -2, -7, 0, 9, 4, 2, -1,
    -- filter=92 channel=50
    16, 6, 12, 8, 16, -6, 12, -2, 9,
    -- filter=92 channel=51
    -9, -8, -6, -7, 8, 8, -10, -2, 1,
    -- filter=92 channel=52
    9, 0, 5, -1, -1, -7, 8, 0, 6,
    -- filter=92 channel=53
    14, 15, -3, 12, -2, 5, 20, 12, 13,
    -- filter=92 channel=54
    0, -5, 10, 1, 6, -2, 5, 0, -2,
    -- filter=92 channel=55
    4, 1, -1, -5, 2, 2, 4, 0, 7,
    -- filter=92 channel=56
    4, 11, -2, -1, 7, -4, 12, 5, -7,
    -- filter=92 channel=57
    -3, -2, 8, -4, 7, -1, -4, 8, -9,
    -- filter=92 channel=58
    -6, -10, 4, -3, -5, -6, -8, 10, -7,
    -- filter=92 channel=59
    -6, -6, 10, -13, 2, 12, -11, -17, -2,
    -- filter=92 channel=60
    -5, 0, 29, -5, -12, 16, 3, -25, 11,
    -- filter=92 channel=61
    6, 2, 8, 2, 0, 1, 9, -18, 1,
    -- filter=92 channel=62
    9, 0, -1, -2, -14, 12, -6, -3, -9,
    -- filter=92 channel=63
    2, 9, 4, 0, 6, 5, -6, -1, 7,
    -- filter=93 channel=0
    -10, 3, 5, 7, 4, 6, 17, 10, 8,
    -- filter=93 channel=1
    6, -9, -14, 9, 2, -1, 8, 6, 4,
    -- filter=93 channel=2
    -2, -6, 5, 9, 7, 0, 5, 2, -11,
    -- filter=93 channel=3
    4, 0, -6, -2, 10, 5, -2, -3, 2,
    -- filter=93 channel=4
    -8, -13, 5, 13, -3, 1, 7, 8, 12,
    -- filter=93 channel=5
    -9, -6, -6, -6, -11, 9, -10, -8, 4,
    -- filter=93 channel=6
    2, -5, 2, 5, -2, 9, 9, -3, 8,
    -- filter=93 channel=7
    -2, 1, -9, -7, -11, 8, -10, -4, 11,
    -- filter=93 channel=8
    -3, 0, -9, -1, 22, 17, -1, 3, 2,
    -- filter=93 channel=9
    -23, -44, -34, -34, -55, -41, -38, -47, -37,
    -- filter=93 channel=10
    6, 16, 8, 2, 21, 11, 12, 5, 1,
    -- filter=93 channel=11
    -8, 0, -9, 8, 13, 9, 7, 18, 9,
    -- filter=93 channel=12
    8, 4, -5, 8, -4, 7, 8, -7, 1,
    -- filter=93 channel=13
    -1, -17, -18, -7, -7, 0, 7, 10, 2,
    -- filter=93 channel=14
    -3, -8, 7, 4, 1, 5, 3, 1, 0,
    -- filter=93 channel=15
    -18, 0, -4, 9, 14, 10, 8, -3, -6,
    -- filter=93 channel=16
    -25, -26, -14, 6, 4, 7, 8, 10, 10,
    -- filter=93 channel=17
    -15, -5, 3, 8, 13, 4, 3, 4, 18,
    -- filter=93 channel=18
    -2, -12, -3, -2, -1, 11, 7, -9, 1,
    -- filter=93 channel=19
    -8, -10, -1, -8, -19, -6, -1, -18, 6,
    -- filter=93 channel=20
    -11, -3, 3, -5, -11, -12, 0, -3, -7,
    -- filter=93 channel=21
    -8, 5, 6, -2, -6, 4, -4, 3, -3,
    -- filter=93 channel=22
    6, 4, 10, 6, -3, 7, -8, 2, 4,
    -- filter=93 channel=23
    6, 11, 1, 13, 20, 7, 19, 27, 15,
    -- filter=93 channel=24
    -4, -8, 4, -8, -2, -6, 13, 13, 0,
    -- filter=93 channel=25
    2, -5, 2, 2, 16, 12, 8, 1, 2,
    -- filter=93 channel=26
    0, 2, 10, 3, 5, -1, 10, 3, 6,
    -- filter=93 channel=27
    -5, 3, 0, 23, 20, 21, 18, 12, 9,
    -- filter=93 channel=28
    -12, -21, -15, -12, -5, -7, -8, -12, 0,
    -- filter=93 channel=29
    -15, -32, -25, -9, -6, -2, -3, -9, -1,
    -- filter=93 channel=30
    -11, -6, 4, 4, -8, 11, -10, 7, 15,
    -- filter=93 channel=31
    9, -5, 4, 3, -1, 9, -6, -3, 10,
    -- filter=93 channel=32
    13, 3, -1, 7, 15, 14, 3, 2, 11,
    -- filter=93 channel=33
    -7, 0, 1, -8, 1, -10, 1, 8, -6,
    -- filter=93 channel=34
    2, -7, -8, 0, -1, 6, 6, -7, -1,
    -- filter=93 channel=35
    12, 25, 10, 26, 37, 18, 20, 28, 10,
    -- filter=93 channel=36
    8, 8, 0, 0, 12, 8, 8, -4, -6,
    -- filter=93 channel=37
    -3, -10, -6, 3, -5, -6, -2, 0, 2,
    -- filter=93 channel=38
    -2, -12, -12, 7, 9, 12, 24, 21, 14,
    -- filter=93 channel=39
    5, -1, -3, -4, 6, 0, 8, 0, 8,
    -- filter=93 channel=40
    -3, 5, -6, 1, 9, 14, 9, 9, 0,
    -- filter=93 channel=41
    -17, -15, -13, 16, 19, 18, 16, 12, 20,
    -- filter=93 channel=42
    -3, 0, 3, 8, -6, 0, 5, 0, 1,
    -- filter=93 channel=43
    -10, -2, 4, -12, -8, 11, 5, 12, 24,
    -- filter=93 channel=44
    11, 7, -4, 2, 14, 7, -5, 0, 2,
    -- filter=93 channel=45
    -5, 8, -1, 9, 9, 7, 2, -9, -4,
    -- filter=93 channel=46
    -15, 0, -9, -8, -8, -4, -11, 3, 1,
    -- filter=93 channel=47
    5, -6, 1, 4, -5, -5, -10, 2, 2,
    -- filter=93 channel=48
    -13, -7, 1, 0, -15, 5, -11, -13, -3,
    -- filter=93 channel=49
    18, 24, 6, 23, 26, 27, 12, 4, 11,
    -- filter=93 channel=50
    0, -6, 11, 1, -13, -6, 9, -2, 13,
    -- filter=93 channel=51
    14, 8, 4, 1, 9, 13, 18, 19, 5,
    -- filter=93 channel=52
    5, 6, -8, -1, 8, -1, -2, -6, -5,
    -- filter=93 channel=53
    7, 4, -8, -3, -5, 6, 7, -2, -1,
    -- filter=93 channel=54
    -11, -30, -28, -20, -29, -14, -22, -33, -18,
    -- filter=93 channel=55
    -8, 9, 3, 5, -6, -9, 7, -8, 4,
    -- filter=93 channel=56
    -1, -8, 8, 0, 0, -2, -7, -5, 0,
    -- filter=93 channel=57
    -1, 8, -9, 3, -9, 0, 0, 10, 9,
    -- filter=93 channel=58
    -7, 0, 13, -10, -4, -5, -6, 6, -8,
    -- filter=93 channel=59
    -8, -9, 5, 5, 15, 5, 8, 17, 14,
    -- filter=93 channel=60
    -8, -16, -20, 3, 13, 17, 8, 27, 16,
    -- filter=93 channel=61
    -12, -14, 1, 0, 14, 18, 5, 12, 10,
    -- filter=93 channel=62
    4, 0, 4, 1, 13, 8, 11, 0, -3,
    -- filter=93 channel=63
    -4, -10, -8, -3, -8, 10, -2, 0, -3,
    -- filter=94 channel=0
    8, 0, 0, -2, 5, -7, -6, -5, -3,
    -- filter=94 channel=1
    4, 5, -10, 3, -6, -5, 9, 0, -8,
    -- filter=94 channel=2
    -5, -5, 0, 4, -2, 8, 4, 4, 3,
    -- filter=94 channel=3
    4, 0, -2, 10, -1, -6, -7, 6, 9,
    -- filter=94 channel=4
    -2, 0, 6, -4, -1, 1, -2, -5, -9,
    -- filter=94 channel=5
    1, -6, 6, -10, -3, 5, -8, 9, 3,
    -- filter=94 channel=6
    7, -2, 0, -8, -2, 5, -1, -7, 2,
    -- filter=94 channel=7
    -5, -5, 10, -2, 5, -4, -8, 9, -3,
    -- filter=94 channel=8
    -10, 2, 0, 8, 2, -3, 5, -5, 8,
    -- filter=94 channel=9
    0, -8, 1, 1, 1, -1, -7, 7, 4,
    -- filter=94 channel=10
    1, 7, -2, 2, 1, 5, -4, 3, 6,
    -- filter=94 channel=11
    -9, -5, -1, 6, 9, 0, -4, -7, 3,
    -- filter=94 channel=12
    -5, 9, -5, -10, -2, -1, 10, -9, -8,
    -- filter=94 channel=13
    7, 2, -5, -1, -10, -1, -4, -6, -1,
    -- filter=94 channel=14
    -5, 8, 2, -5, -4, -8, 6, 1, -4,
    -- filter=94 channel=15
    0, -3, -6, -3, -6, -2, -10, 7, 2,
    -- filter=94 channel=16
    7, -4, 6, 7, 9, -6, 3, -2, -8,
    -- filter=94 channel=17
    6, -2, -10, -1, 0, 3, 6, 6, -7,
    -- filter=94 channel=18
    -1, 5, -5, 7, -4, 0, 0, -1, 3,
    -- filter=94 channel=19
    8, 3, 8, 0, 5, 0, 0, -10, -1,
    -- filter=94 channel=20
    -1, 3, 5, 0, 9, 1, 3, 5, -9,
    -- filter=94 channel=21
    -3, 2, -5, 0, 10, 6, -1, -8, 4,
    -- filter=94 channel=22
    -3, -1, -4, 6, -10, 0, 10, 7, -8,
    -- filter=94 channel=23
    -8, -3, -2, 5, 1, -8, 9, 1, -10,
    -- filter=94 channel=24
    -6, -6, 3, 7, -8, 2, -4, 1, -8,
    -- filter=94 channel=25
    10, -5, 3, -9, 0, 3, 0, 5, -7,
    -- filter=94 channel=26
    -8, -7, -10, -9, 9, 6, -8, -1, 8,
    -- filter=94 channel=27
    -9, 2, 0, 0, -6, -5, -7, 4, -7,
    -- filter=94 channel=28
    -7, 4, -11, -10, 0, -5, 9, 0, 3,
    -- filter=94 channel=29
    -10, -1, 1, 3, -10, 3, -3, 3, -1,
    -- filter=94 channel=30
    2, 6, -6, 4, 1, 9, -3, 1, 6,
    -- filter=94 channel=31
    9, 1, -8, -6, 1, -1, 2, 7, -9,
    -- filter=94 channel=32
    4, 10, 6, -8, -2, 8, -5, -5, -10,
    -- filter=94 channel=33
    -6, 2, -7, -3, -4, 4, -1, 7, -4,
    -- filter=94 channel=34
    -1, 9, 1, -6, 4, 1, 7, -2, 6,
    -- filter=94 channel=35
    -1, 0, -4, -5, 2, -10, -5, 7, -1,
    -- filter=94 channel=36
    5, -9, -1, -6, 5, -2, -7, -10, 4,
    -- filter=94 channel=37
    1, -5, 7, 0, 8, -4, -3, 8, 0,
    -- filter=94 channel=38
    10, 1, -9, 7, -9, 8, -3, -9, 7,
    -- filter=94 channel=39
    -8, 3, 7, -6, -7, 1, -9, -5, 0,
    -- filter=94 channel=40
    4, -10, -5, 5, -7, -1, 0, -4, 7,
    -- filter=94 channel=41
    0, -7, 7, -9, -9, -8, -10, 1, 7,
    -- filter=94 channel=42
    0, 9, -10, 1, 4, 5, -5, 0, -8,
    -- filter=94 channel=43
    -7, -9, 8, -8, 0, -8, -9, 5, -5,
    -- filter=94 channel=44
    -2, -2, -8, -1, 0, -6, 2, -3, 5,
    -- filter=94 channel=45
    -6, -7, 10, -9, -10, 9, 1, 0, -2,
    -- filter=94 channel=46
    8, -7, -4, 7, 7, 5, -6, -3, 7,
    -- filter=94 channel=47
    0, -7, -1, -10, -6, -10, -6, 8, 2,
    -- filter=94 channel=48
    -4, 9, 4, 1, 8, 0, 0, 6, -4,
    -- filter=94 channel=49
    0, 6, -5, 9, -4, 9, 5, 7, -4,
    -- filter=94 channel=50
    2, 0, 0, 3, 2, -2, -6, 0, 1,
    -- filter=94 channel=51
    -6, -6, 7, -5, 1, 8, 3, 9, 2,
    -- filter=94 channel=52
    -3, -2, -4, -10, 7, -8, 0, 7, 4,
    -- filter=94 channel=53
    3, -7, -3, -3, 2, -6, 2, -6, 2,
    -- filter=94 channel=54
    7, -8, 1, -8, 2, 4, 3, 1, -2,
    -- filter=94 channel=55
    1, -3, -9, 8, -9, 7, -8, -1, -3,
    -- filter=94 channel=56
    8, -4, -1, 6, 0, -6, 8, -2, 4,
    -- filter=94 channel=57
    10, 5, -4, 0, 8, 10, -10, -3, 6,
    -- filter=94 channel=58
    -9, 6, 8, 5, -9, -8, 3, -5, -10,
    -- filter=94 channel=59
    -2, -5, 8, -1, 6, 1, -9, 7, 3,
    -- filter=94 channel=60
    -5, -7, -2, 6, 3, -2, -8, 8, 1,
    -- filter=94 channel=61
    -6, 0, -6, -3, 3, -6, 0, -3, 7,
    -- filter=94 channel=62
    10, 1, 7, 0, 3, -7, -10, -3, -2,
    -- filter=94 channel=63
    -6, 2, -6, 8, -3, -4, 6, -1, -3,
    -- filter=95 channel=0
    -1, 6, -2, 8, 9, 10, -3, -12, -5,
    -- filter=95 channel=1
    -2, -6, 5, 2, 10, -2, 0, -11, -8,
    -- filter=95 channel=2
    -9, -3, -6, -6, -13, -7, 4, -6, 2,
    -- filter=95 channel=3
    0, -6, 0, 9, -4, -6, 7, 6, 4,
    -- filter=95 channel=4
    1, 9, 1, 3, 6, 10, 10, 2, -11,
    -- filter=95 channel=5
    -10, 5, -6, -4, -6, -3, -5, -1, 5,
    -- filter=95 channel=6
    2, 7, -6, 2, 0, -1, 5, -2, 1,
    -- filter=95 channel=7
    8, 6, -9, 8, -5, -8, 4, 1, 8,
    -- filter=95 channel=8
    -2, 14, -4, -3, -7, 9, -7, -11, 0,
    -- filter=95 channel=9
    -7, -6, -3, 0, -8, 12, 5, 1, 11,
    -- filter=95 channel=10
    6, 9, 8, 7, -6, 5, 0, -10, -10,
    -- filter=95 channel=11
    -6, 11, 10, -9, 2, -1, 0, 3, -14,
    -- filter=95 channel=12
    10, 1, -9, 8, 7, 4, -3, 0, -1,
    -- filter=95 channel=13
    5, -1, 6, 0, -8, 11, 3, -1, -7,
    -- filter=95 channel=14
    -7, -4, 10, -4, 2, 3, 1, -2, 5,
    -- filter=95 channel=15
    5, 5, -2, 7, -5, 2, 4, -12, -8,
    -- filter=95 channel=16
    -6, 11, 7, -7, -8, 8, 0, -7, -11,
    -- filter=95 channel=17
    -1, 13, 5, -8, 10, -7, 3, 2, -9,
    -- filter=95 channel=18
    4, -7, -7, 4, 3, -8, -4, 3, -10,
    -- filter=95 channel=19
    -9, -1, 0, 5, 9, 7, -8, -3, 6,
    -- filter=95 channel=20
    6, -7, -4, 0, 4, 0, -6, 0, 11,
    -- filter=95 channel=21
    5, -5, 5, 1, -7, -4, 0, 2, -3,
    -- filter=95 channel=22
    4, 2, -7, -9, -1, 4, 2, 0, -6,
    -- filter=95 channel=23
    -8, 5, 2, -3, -4, -4, 10, -1, -12,
    -- filter=95 channel=24
    -6, -3, -7, 9, -5, 4, 1, -2, -3,
    -- filter=95 channel=25
    -4, -4, 3, 8, -13, -4, 7, -12, -12,
    -- filter=95 channel=26
    2, 8, 8, -2, 7, 0, 0, 9, -6,
    -- filter=95 channel=27
    -6, 9, 2, 0, 6, 0, 4, 3, -10,
    -- filter=95 channel=28
    -10, -8, 4, 3, -9, -7, 3, -5, 7,
    -- filter=95 channel=29
    5, 0, 8, 10, 3, -6, -3, 4, -5,
    -- filter=95 channel=30
    -10, 8, 1, -1, 3, 8, 7, 16, 6,
    -- filter=95 channel=31
    -1, 8, 4, 2, 3, -8, 8, 2, 9,
    -- filter=95 channel=32
    4, -3, -7, 9, 0, -4, -3, -3, -4,
    -- filter=95 channel=33
    -3, 8, 7, 5, -9, -5, 2, 4, -7,
    -- filter=95 channel=34
    -6, -4, 8, -6, 9, 3, -6, -1, -2,
    -- filter=95 channel=35
    0, 3, 2, 0, -3, -10, 0, 0, 5,
    -- filter=95 channel=36
    1, 0, -5, 1, -7, -2, 10, -1, 4,
    -- filter=95 channel=37
    -3, 8, 3, -6, 0, -4, 9, 5, 4,
    -- filter=95 channel=38
    8, 4, -4, -5, -9, 0, 10, -7, -2,
    -- filter=95 channel=39
    2, 8, -2, -3, 4, 7, 0, 7, 1,
    -- filter=95 channel=40
    11, 0, 9, -3, 9, -7, 0, -5, -7,
    -- filter=95 channel=41
    -7, 6, 3, -3, 9, -8, 6, -11, 6,
    -- filter=95 channel=42
    -9, 4, 1, -7, -6, 0, -3, -8, 3,
    -- filter=95 channel=43
    -8, -1, 3, 8, 8, -1, 2, 9, 0,
    -- filter=95 channel=44
    -9, 7, -6, -4, -1, -6, -2, 11, 0,
    -- filter=95 channel=45
    2, 0, 7, 9, 0, 6, 1, 6, -10,
    -- filter=95 channel=46
    5, -4, -5, 11, -8, -3, -9, -4, -3,
    -- filter=95 channel=47
    -3, 6, 8, -2, -2, 2, -8, -6, 7,
    -- filter=95 channel=48
    2, 7, -9, -7, 6, -3, -2, -8, -1,
    -- filter=95 channel=49
    -1, 10, 0, 1, -6, -3, -7, -10, -11,
    -- filter=95 channel=50
    -2, 2, 2, -8, 1, 9, 4, -1, 2,
    -- filter=95 channel=51
    -5, 7, 0, 2, 8, 11, 4, -6, -7,
    -- filter=95 channel=52
    -5, -7, -6, -8, -9, 7, 0, -10, 6,
    -- filter=95 channel=53
    4, -8, -8, -4, -2, 0, 6, 3, -7,
    -- filter=95 channel=54
    -4, 11, 0, 0, 10, 9, -9, 12, 6,
    -- filter=95 channel=55
    -4, -8, 5, 0, -4, -7, -1, 0, -2,
    -- filter=95 channel=56
    0, 8, -8, -2, -6, -6, -2, 9, -7,
    -- filter=95 channel=57
    -10, 7, -10, -7, 4, 7, 2, -6, 4,
    -- filter=95 channel=58
    6, 0, -1, -3, -3, 9, -1, -1, 10,
    -- filter=95 channel=59
    0, 9, 6, 5, 1, 7, 8, -8, -5,
    -- filter=95 channel=60
    6, 13, 3, 13, 2, -2, -5, -7, 3,
    -- filter=95 channel=61
    -5, 13, 9, 5, 9, -5, 12, -1, -13,
    -- filter=95 channel=62
    4, 1, -3, -1, -3, -3, 10, -2, -10,
    -- filter=95 channel=63
    -4, 1, -10, 0, 2, 2, 4, -6, 5,
    -- filter=96 channel=0
    -5, 0, 5, -4, 4, 3, -1, -4, 0,
    -- filter=96 channel=1
    1, 3, 4, 16, 0, 2, 10, -8, -2,
    -- filter=96 channel=2
    13, -2, -6, -4, 7, 7, -3, 5, -9,
    -- filter=96 channel=3
    12, 6, 0, 7, -5, -1, -4, 8, 6,
    -- filter=96 channel=4
    11, -8, -3, 9, 0, 0, 0, -8, 7,
    -- filter=96 channel=5
    -1, 9, 6, 4, -2, -7, -5, -3, 2,
    -- filter=96 channel=6
    -6, 9, -7, 2, 10, -3, 11, 5, 7,
    -- filter=96 channel=7
    9, 0, -7, 2, -10, 1, -5, 8, -2,
    -- filter=96 channel=8
    12, 5, -1, 5, -9, -8, -3, 6, 3,
    -- filter=96 channel=9
    -6, -2, 0, -4, -5, 9, -9, -5, 0,
    -- filter=96 channel=10
    8, -1, 5, 2, 8, -2, 9, -7, -4,
    -- filter=96 channel=11
    5, -4, 4, 2, 1, 3, -5, 1, 5,
    -- filter=96 channel=12
    -8, -7, 0, 10, 0, 6, 6, 6, -6,
    -- filter=96 channel=13
    4, 2, -5, -2, -9, -4, -2, -1, -1,
    -- filter=96 channel=14
    -3, -6, -6, 9, 7, -2, 3, -9, 3,
    -- filter=96 channel=15
    12, 2, 3, 12, -4, 1, -2, 1, 6,
    -- filter=96 channel=16
    6, -4, -2, 0, 11, -3, 17, -6, -8,
    -- filter=96 channel=17
    -2, 6, 0, -5, 9, -1, 9, 2, 8,
    -- filter=96 channel=18
    -10, -9, -2, 6, -6, 8, -8, 0, 11,
    -- filter=96 channel=19
    3, 4, 6, 5, -2, 11, -5, 8, 2,
    -- filter=96 channel=20
    -2, -12, -9, -1, -2, 7, 0, 6, -7,
    -- filter=96 channel=21
    2, 2, 4, 7, -2, -7, 3, 9, 7,
    -- filter=96 channel=22
    1, -2, 5, -3, 7, 5, -4, -1, -6,
    -- filter=96 channel=23
    -3, -8, 10, -6, 5, -7, -2, 2, -4,
    -- filter=96 channel=24
    1, 0, 7, 8, -6, 3, 6, -4, 0,
    -- filter=96 channel=25
    4, 10, 0, -4, 10, -7, 13, -6, 8,
    -- filter=96 channel=26
    -2, -4, -4, -4, -3, 0, 1, 0, -10,
    -- filter=96 channel=27
    6, 2, 0, 15, 8, -5, -4, -4, 6,
    -- filter=96 channel=28
    15, -2, 2, 4, -3, 4, 0, 4, 0,
    -- filter=96 channel=29
    7, -4, -10, 13, 7, 0, 13, -8, -7,
    -- filter=96 channel=30
    -8, -8, 0, -2, -4, -14, -12, -4, 0,
    -- filter=96 channel=31
    0, -8, 8, -3, -5, 9, -9, 9, 10,
    -- filter=96 channel=32
    5, -9, -8, -8, 4, -9, -9, 1, -3,
    -- filter=96 channel=33
    -5, 5, 8, -9, 9, 6, -2, -6, 7,
    -- filter=96 channel=34
    3, 0, -1, -3, -6, -5, -1, -12, -8,
    -- filter=96 channel=35
    -4, -8, -4, 12, 1, -11, 6, 5, -6,
    -- filter=96 channel=36
    0, 0, -2, -4, 8, 6, 2, 8, 10,
    -- filter=96 channel=37
    10, -9, -8, 7, 5, -9, -7, 0, 3,
    -- filter=96 channel=38
    16, 10, -9, 0, 3, -5, -5, 0, 7,
    -- filter=96 channel=39
    -9, 1, -5, -1, -10, 8, -2, -3, -8,
    -- filter=96 channel=40
    7, 9, -5, -4, -10, -11, 0, -8, -11,
    -- filter=96 channel=41
    13, -9, -12, 5, -10, -12, 8, 8, -13,
    -- filter=96 channel=42
    2, 8, -7, -3, 10, 8, -1, -3, 0,
    -- filter=96 channel=43
    -1, 0, 4, -3, 7, 1, 0, 3, 4,
    -- filter=96 channel=44
    6, 2, -7, 11, -4, -2, 4, 1, 0,
    -- filter=96 channel=45
    0, -3, -1, -8, -8, 0, 2, 0, 1,
    -- filter=96 channel=46
    -7, -10, -10, -14, 5, 0, -9, -9, -9,
    -- filter=96 channel=47
    -4, 10, -8, 10, -9, -8, 8, 0, 10,
    -- filter=96 channel=48
    9, -6, -1, 4, -4, 3, -8, 2, 8,
    -- filter=96 channel=49
    0, 8, 5, 1, -2, -4, -4, 8, 1,
    -- filter=96 channel=50
    4, -7, 4, -4, 8, -8, 0, -13, -10,
    -- filter=96 channel=51
    4, 9, 3, -8, 9, 0, -1, -3, -9,
    -- filter=96 channel=52
    -10, -6, -8, 4, 7, 8, -7, -8, -8,
    -- filter=96 channel=53
    -5, -6, -7, 0, -7, 6, -2, -10, -3,
    -- filter=96 channel=54
    1, -8, -3, 4, -5, 6, 2, 8, 6,
    -- filter=96 channel=55
    3, 8, -6, 8, 4, 9, -1, 0, 7,
    -- filter=96 channel=56
    -8, 5, -3, 3, 7, -8, 1, -6, 1,
    -- filter=96 channel=57
    4, 3, 2, -2, 4, -4, 10, 9, -4,
    -- filter=96 channel=58
    3, 10, 9, 5, 10, -8, 2, -4, 9,
    -- filter=96 channel=59
    6, -5, -8, -7, 5, -10, 11, -5, 0,
    -- filter=96 channel=60
    -5, -4, -4, 11, -10, -5, 5, -1, -13,
    -- filter=96 channel=61
    12, 7, -11, 0, -1, 6, 2, -4, 0,
    -- filter=96 channel=62
    -3, 1, 5, -4, -1, -5, 9, 10, 6,
    -- filter=96 channel=63
    -10, -9, 1, -7, 0, -7, 10, 2, -5,
    -- filter=97 channel=0
    0, 16, 0, -5, 6, 3, -13, -10, -7,
    -- filter=97 channel=1
    5, 12, 3, 12, 10, 7, 0, 4, 5,
    -- filter=97 channel=2
    0, 11, 3, 1, -10, -7, -1, -4, -10,
    -- filter=97 channel=3
    4, -5, 5, -13, -7, -5, -11, -7, -7,
    -- filter=97 channel=4
    12, 8, 16, -12, 3, -6, -2, 2, 0,
    -- filter=97 channel=5
    -5, 0, 8, 2, -13, -2, 2, 3, -8,
    -- filter=97 channel=6
    5, 11, 9, -6, 0, -9, -12, 1, -6,
    -- filter=97 channel=7
    -2, 5, -6, -1, -8, -7, 2, 0, -1,
    -- filter=97 channel=8
    9, 18, 13, -5, -5, -1, -13, -3, 0,
    -- filter=97 channel=9
    -4, 2, 4, 6, 5, 0, -9, -16, -12,
    -- filter=97 channel=10
    0, 0, -4, 10, 16, 8, 11, 0, -6,
    -- filter=97 channel=11
    10, 0, 15, 3, 9, -3, -1, -8, 0,
    -- filter=97 channel=12
    2, -9, 7, -1, -3, 4, 7, -9, -5,
    -- filter=97 channel=13
    8, 3, 16, 13, 6, -2, -17, -9, -8,
    -- filter=97 channel=14
    -5, 3, -9, -5, 8, -9, -2, 2, 3,
    -- filter=97 channel=15
    14, 16, 22, -14, -11, -4, -14, -13, -6,
    -- filter=97 channel=16
    26, 24, 21, -9, -7, -7, -9, -18, -7,
    -- filter=97 channel=17
    16, 18, 10, 2, 4, -4, -14, -7, -4,
    -- filter=97 channel=18
    13, -1, 2, 6, -4, 12, -8, 7, 8,
    -- filter=97 channel=19
    -8, 5, 6, 4, 1, -10, 10, 2, -12,
    -- filter=97 channel=20
    4, 6, 4, -4, -2, -8, 8, -4, -2,
    -- filter=97 channel=21
    5, 9, 9, -4, -8, 2, 8, 3, -1,
    -- filter=97 channel=22
    0, -5, -5, 7, -2, -4, 0, 2, -3,
    -- filter=97 channel=23
    0, 12, 12, -3, -2, -5, 0, -7, 9,
    -- filter=97 channel=24
    10, 17, 0, 8, 7, 5, 1, -8, -9,
    -- filter=97 channel=25
    9, 10, 6, -1, -11, -13, -4, -2, 2,
    -- filter=97 channel=26
    9, 3, -1, -9, 2, -3, 5, 1, 7,
    -- filter=97 channel=27
    16, 0, 0, -2, -8, -17, -14, -6, -1,
    -- filter=97 channel=28
    20, 12, 19, -10, -11, -9, -5, -3, 4,
    -- filter=97 channel=29
    30, 19, 11, -16, -12, -10, -9, -12, -1,
    -- filter=97 channel=30
    -6, -8, -4, 6, -7, -7, -7, -16, 1,
    -- filter=97 channel=31
    4, 2, -9, -2, 6, 9, -8, -8, 7,
    -- filter=97 channel=32
    -7, 8, 7, 13, -3, 7, 0, 1, -13,
    -- filter=97 channel=33
    10, 1, 4, 6, -7, -9, -4, -7, 7,
    -- filter=97 channel=34
    -4, 2, -3, 6, -9, 5, 6, -5, 2,
    -- filter=97 channel=35
    0, 8, -4, -5, 0, -4, 7, 0, 2,
    -- filter=97 channel=36
    0, 1, 7, 2, 10, -6, 7, -6, 0,
    -- filter=97 channel=37
    4, 1, 10, -6, -6, 5, 0, 4, -3,
    -- filter=97 channel=38
    5, 17, 6, -4, 1, -5, -20, -22, -17,
    -- filter=97 channel=39
    -6, -3, 7, 0, -7, 1, 1, 4, -9,
    -- filter=97 channel=40
    7, 1, -7, -8, 1, -11, 5, 4, 3,
    -- filter=97 channel=41
    23, 21, 25, -7, -20, -19, -18, -18, -9,
    -- filter=97 channel=42
    1, 10, 6, -9, -5, -6, 8, -2, -8,
    -- filter=97 channel=43
    12, 21, 2, 28, 25, 23, 1, 5, 2,
    -- filter=97 channel=44
    0, 4, 0, 5, 2, -4, -3, -1, -10,
    -- filter=97 channel=45
    -7, 7, 0, -2, 2, 1, -3, 0, 8,
    -- filter=97 channel=46
    -1, -1, 0, -3, -8, -3, -7, 7, -10,
    -- filter=97 channel=47
    -7, -1, 6, 10, 1, 8, 6, 8, 4,
    -- filter=97 channel=48
    11, 8, -3, -1, -1, -9, -13, -5, -2,
    -- filter=97 channel=49
    14, 7, -1, -4, -17, -15, 11, 4, -7,
    -- filter=97 channel=50
    9, 0, 4, 10, 13, 13, -5, -10, 3,
    -- filter=97 channel=51
    -2, 0, -5, 9, 13, 13, -4, 4, 10,
    -- filter=97 channel=52
    -4, -5, 7, -3, -1, -8, -6, -7, -6,
    -- filter=97 channel=53
    4, 5, -8, 0, -5, 5, -4, -14, -16,
    -- filter=97 channel=54
    5, 0, -3, -7, -4, -9, -16, -7, -5,
    -- filter=97 channel=55
    3, -6, 2, -5, -8, -5, 5, -10, -4,
    -- filter=97 channel=56
    8, -4, 8, 5, -6, 0, -7, 8, -10,
    -- filter=97 channel=57
    -9, -2, 3, -3, 9, 0, 4, -1, 2,
    -- filter=97 channel=58
    0, 3, 6, 2, -3, -4, 3, 12, -3,
    -- filter=97 channel=59
    16, 16, 15, 2, 1, -11, -8, -11, 2,
    -- filter=97 channel=60
    32, 15, 20, 0, 0, 7, -15, -23, -4,
    -- filter=97 channel=61
    15, 17, 5, 1, -9, 3, -22, -6, -12,
    -- filter=97 channel=62
    0, 2, 6, 0, -2, -11, -6, -3, -4,
    -- filter=97 channel=63
    -6, -4, 3, -8, -8, 3, 2, 8, 9,
    -- filter=98 channel=0
    -6, 10, -13, 9, 3, -6, -3, 5, -1,
    -- filter=98 channel=1
    -6, 2, 6, 0, -6, 10, -12, 9, -2,
    -- filter=98 channel=2
    0, 9, -3, 5, 4, 5, -3, -11, -26,
    -- filter=98 channel=3
    3, 26, 12, 8, 24, 17, 19, 12, 2,
    -- filter=98 channel=4
    -1, -5, -13, 5, -2, 0, -12, 2, -13,
    -- filter=98 channel=5
    -7, -1, 0, -4, -7, 14, 6, 4, -2,
    -- filter=98 channel=6
    1, 0, -7, 1, 9, 1, 0, -10, -19,
    -- filter=98 channel=7
    -10, 1, -2, -12, -1, 2, -9, -9, -13,
    -- filter=98 channel=8
    -2, 11, 10, 15, 28, 2, -15, -5, -21,
    -- filter=98 channel=9
    -9, -12, -20, -11, 2, -17, 0, -19, -10,
    -- filter=98 channel=10
    -14, 0, 0, -16, -7, 0, 0, -8, 10,
    -- filter=98 channel=11
    -14, 3, -1, -3, 4, 4, -5, -5, 8,
    -- filter=98 channel=12
    -2, -2, -7, 9, 2, 9, -7, 9, -1,
    -- filter=98 channel=13
    6, -9, -12, 1, -3, -15, -8, -5, -10,
    -- filter=98 channel=14
    -12, -13, 2, -8, 4, -9, 0, -7, -11,
    -- filter=98 channel=15
    9, 21, -10, -1, 23, -6, -19, -12, -15,
    -- filter=98 channel=16
    14, 2, -15, 7, 30, 0, -1, -14, -33,
    -- filter=98 channel=17
    6, 15, 17, 8, 19, 14, -14, 0, 4,
    -- filter=98 channel=18
    -7, 0, -10, -14, -10, -12, -9, -21, -9,
    -- filter=98 channel=19
    -19, -16, 3, -20, -14, -2, -14, -1, -12,
    -- filter=98 channel=20
    -16, 0, -6, -7, -9, -19, -13, -19, -19,
    -- filter=98 channel=21
    12, 0, -7, 0, 4, 9, 5, 2, -3,
    -- filter=98 channel=22
    -7, 1, 0, 0, -5, 3, 9, 10, 4,
    -- filter=98 channel=23
    0, 7, 1, -14, 1, -4, 1, 0, -1,
    -- filter=98 channel=24
    -7, 5, 1, -9, 8, 10, 0, 13, 1,
    -- filter=98 channel=25
    0, 12, 5, 9, 18, 0, 1, -3, -2,
    -- filter=98 channel=26
    -7, -18, -20, -7, 0, -4, 0, -7, -20,
    -- filter=98 channel=27
    19, 19, 7, 8, 22, 5, -1, 0, -10,
    -- filter=98 channel=28
    -13, 0, -14, -11, 4, 5, -12, -16, -15,
    -- filter=98 channel=29
    0, 12, -18, 20, 16, -5, -1, -6, -39,
    -- filter=98 channel=30
    -17, -18, -8, -29, -13, -11, -30, -10, -13,
    -- filter=98 channel=31
    -2, 6, 6, 6, 7, 2, 2, -9, 7,
    -- filter=98 channel=32
    -11, -1, -6, -10, 2, -4, -1, 9, -1,
    -- filter=98 channel=33
    -7, -6, 6, -2, 6, 3, 9, -9, 0,
    -- filter=98 channel=34
    3, 6, -5, -7, -12, -8, -13, -13, -10,
    -- filter=98 channel=35
    6, 5, 4, -2, 15, 13, -1, -3, 0,
    -- filter=98 channel=36
    -9, 9, 5, 5, -8, 9, 2, 0, 0,
    -- filter=98 channel=37
    1, 5, 13, 10, 16, 14, 13, 10, 12,
    -- filter=98 channel=38
    10, 10, 0, 9, 28, 16, -4, 17, -14,
    -- filter=98 channel=39
    -8, -2, 4, -3, 3, -8, -1, -6, 0,
    -- filter=98 channel=40
    10, 14, 8, 1, 0, 5, -5, -6, 8,
    -- filter=98 channel=41
    16, 19, 15, 22, 37, 21, 1, 10, -19,
    -- filter=98 channel=42
    1, -7, 0, 1, 0, -7, 8, -5, 3,
    -- filter=98 channel=43
    -24, -28, -26, -8, -6, -13, -14, -2, -5,
    -- filter=98 channel=44
    -8, 1, -1, -17, -8, -1, -17, -11, -7,
    -- filter=98 channel=45
    -9, -7, -7, -6, 7, 0, 3, -6, -7,
    -- filter=98 channel=46
    0, 1, -10, -9, -2, -22, -6, -12, -21,
    -- filter=98 channel=47
    6, -3, 6, 2, 3, 6, 4, 10, 9,
    -- filter=98 channel=48
    -5, 0, -9, 3, -2, -3, 6, -8, -6,
    -- filter=98 channel=49
    -7, 17, 2, 4, -1, -4, -9, -14, -1,
    -- filter=98 channel=50
    -14, -24, -1, -9, -27, -3, -8, -4, -18,
    -- filter=98 channel=51
    -14, 2, -7, -12, -6, 5, -5, -8, 0,
    -- filter=98 channel=52
    4, -1, -3, -7, -8, 4, -3, -1, -7,
    -- filter=98 channel=53
    -22, -4, -7, -17, -10, -10, -10, -4, 4,
    -- filter=98 channel=54
    2, 11, 8, 0, -1, 11, 0, 5, -4,
    -- filter=98 channel=55
    3, 10, 6, -9, 5, 0, 4, -1, -5,
    -- filter=98 channel=56
    5, -12, -3, 0, 2, -9, -10, 6, 7,
    -- filter=98 channel=57
    -4, -3, -7, -8, 0, 1, 7, -9, 0,
    -- filter=98 channel=58
    -9, -14, -10, -18, -5, -13, -1, -1, -2,
    -- filter=98 channel=59
    23, 30, 16, 11, 15, 16, 0, 6, -7,
    -- filter=98 channel=60
    17, 28, 7, 21, 44, 21, 6, 4, -19,
    -- filter=98 channel=61
    -3, 2, 10, -1, 32, 19, -10, 18, 6,
    -- filter=98 channel=62
    1, 26, 14, 6, 25, 2, 15, 3, -5,
    -- filter=98 channel=63
    -5, 4, 7, -9, -4, 1, 0, 5, 1,
    -- filter=99 channel=0
    5, 16, 10, 6, 18, 25, 7, 15, 13,
    -- filter=99 channel=1
    -31, -36, -21, -30, -38, -17, -24, -26, -20,
    -- filter=99 channel=2
    -25, -25, -8, -21, -27, -12, -16, -20, -33,
    -- filter=99 channel=3
    -8, 13, 14, 4, 0, 19, -9, -7, 0,
    -- filter=99 channel=4
    7, 5, 10, 13, 27, 20, -5, 3, 2,
    -- filter=99 channel=5
    1, 0, 16, 12, 13, 9, 7, 5, 15,
    -- filter=99 channel=6
    -14, 8, -1, -9, -1, -7, -11, -13, -8,
    -- filter=99 channel=7
    12, 2, 4, -2, 4, 2, 5, 12, 9,
    -- filter=99 channel=8
    -4, 25, 27, -6, 34, 30, -10, 6, 21,
    -- filter=99 channel=9
    6, 5, 12, -4, 11, 0, -14, 11, 3,
    -- filter=99 channel=10
    4, -6, 0, -14, -6, 0, 3, 2, 7,
    -- filter=99 channel=11
    0, -1, -1, -7, 0, 11, -10, -2, 0,
    -- filter=99 channel=12
    0, -5, 0, 0, 2, 6, 1, -4, 1,
    -- filter=99 channel=13
    -2, 20, 17, 8, 30, 16, 8, 15, 14,
    -- filter=99 channel=14
    0, -6, 3, -2, -6, 2, 13, -3, 13,
    -- filter=99 channel=15
    3, 28, 22, -4, 21, 34, -13, 20, 14,
    -- filter=99 channel=16
    -17, -7, -3, -18, 12, 1, -20, 6, 0,
    -- filter=99 channel=17
    -6, 1, 27, 0, 12, 16, -1, 3, 19,
    -- filter=99 channel=18
    14, 33, 24, 13, 39, 27, 21, 15, 10,
    -- filter=99 channel=19
    -10, -21, -21, -16, -10, -13, -16, -7, -4,
    -- filter=99 channel=20
    3, 2, 10, 0, 2, 0, 12, 10, -7,
    -- filter=99 channel=21
    6, -9, -2, 8, 5, 0, -1, -4, -1,
    -- filter=99 channel=22
    0, 8, -8, 9, 0, -7, 0, 5, -1,
    -- filter=99 channel=23
    -20, -15, -9, -15, -1, -6, -9, 0, 0,
    -- filter=99 channel=24
    -7, 1, 6, -3, 19, 10, -8, 5, 16,
    -- filter=99 channel=25
    -34, -32, -29, -35, -32, -33, -24, -41, -25,
    -- filter=99 channel=26
    3, 7, -5, 1, -6, -7, -5, -10, -8,
    -- filter=99 channel=27
    -20, -5, 5, -24, -23, -6, -15, -19, 3,
    -- filter=99 channel=28
    -5, 2, 3, 0, 13, 14, -8, -1, -7,
    -- filter=99 channel=29
    -8, 25, 6, -4, 27, 14, 0, 5, 6,
    -- filter=99 channel=30
    -3, 6, 2, 5, 0, 0, 9, -9, 4,
    -- filter=99 channel=31
    2, 11, 10, -5, 11, 7, 4, -5, 2,
    -- filter=99 channel=32
    -21, -10, -7, -7, -22, -14, -5, -10, -7,
    -- filter=99 channel=33
    5, -7, 0, 1, 4, -9, 8, 8, -8,
    -- filter=99 channel=34
    6, 10, 12, -3, 14, 0, 0, 5, 5,
    -- filter=99 channel=35
    -32, -27, -6, -25, -35, -8, -28, -30, -13,
    -- filter=99 channel=36
    -2, 4, -2, 1, -2, 6, 8, 1, 10,
    -- filter=99 channel=37
    -2, 10, -1, -8, 8, 2, -10, -6, -9,
    -- filter=99 channel=38
    -5, -9, 4, -21, 5, 11, -9, 0, 9,
    -- filter=99 channel=39
    -9, 1, 5, 5, 3, -1, 2, -8, 10,
    -- filter=99 channel=40
    -3, -1, -3, -10, -4, -6, -13, -16, 0,
    -- filter=99 channel=41
    -15, 7, 13, 1, 11, 27, -1, 8, 5,
    -- filter=99 channel=42
    -9, -8, 0, 0, 0, 4, -6, -6, -10,
    -- filter=99 channel=43
    -28, -44, -40, -25, -33, -23, -25, -26, -16,
    -- filter=99 channel=44
    -13, -16, -4, -22, -15, 0, -5, -14, -2,
    -- filter=99 channel=45
    -9, 0, 8, 8, 2, 1, 8, 2, -8,
    -- filter=99 channel=46
    3, 9, 4, 21, 11, -1, 17, 2, -2,
    -- filter=99 channel=47
    0, -6, -3, -2, -4, 0, 2, -8, 0,
    -- filter=99 channel=48
    3, 19, 0, 9, 15, 2, -1, -5, 7,
    -- filter=99 channel=49
    -10, 8, 19, 5, 18, 17, -4, 4, 6,
    -- filter=99 channel=50
    6, -2, -1, 11, -16, -2, 10, -2, -2,
    -- filter=99 channel=51
    17, 5, 6, 0, 26, 7, 13, 23, 23,
    -- filter=99 channel=52
    -8, 1, 1, 1, -6, 0, 1, -7, 2,
    -- filter=99 channel=53
    -11, -13, 0, -7, -21, 7, 0, -16, 0,
    -- filter=99 channel=54
    6, 10, 15, 8, 13, 6, 0, -6, 2,
    -- filter=99 channel=55
    -5, 4, -5, 6, 0, -7, -4, 5, -3,
    -- filter=99 channel=56
    0, 0, 4, 4, 3, 4, 1, -1, 5,
    -- filter=99 channel=57
    -2, -5, -4, -2, 0, -6, -4, 0, 3,
    -- filter=99 channel=58
    -2, 4, -9, -8, -1, 0, 1, -5, 8,
    -- filter=99 channel=59
    0, 2, 14, -22, 2, 7, -13, -14, -2,
    -- filter=99 channel=60
    9, 35, 38, 9, 42, 47, 5, 28, 37,
    -- filter=99 channel=61
    1, 7, 12, -5, 18, 31, -5, 11, 21,
    -- filter=99 channel=62
    -11, 5, -3, -12, -7, 13, 0, -7, 6,
    -- filter=99 channel=63
    -3, 7, 2, -6, -5, -4, 8, -3, -4,
    -- filter=100 channel=0
    11, -1, 14, 8, 2, 8, 2, -13, 7,
    -- filter=100 channel=1
    0, -8, 3, 5, 4, -5, 2, 3, -4,
    -- filter=100 channel=2
    5, -2, -1, 0, -16, 6, -7, -4, 7,
    -- filter=100 channel=3
    5, -5, -4, -6, -1, 10, 8, 0, 2,
    -- filter=100 channel=4
    9, 0, 8, 4, 3, 3, -6, -1, 9,
    -- filter=100 channel=5
    4, 6, 0, -1, 11, 0, -1, -4, -4,
    -- filter=100 channel=6
    0, -9, -4, -6, 4, -1, 0, -13, -5,
    -- filter=100 channel=7
    2, 6, 3, -1, 16, 5, -6, 7, -7,
    -- filter=100 channel=8
    5, -6, 2, 1, -21, -4, 3, 4, 12,
    -- filter=100 channel=9
    7, -11, 7, -3, -5, -8, 6, 3, 0,
    -- filter=100 channel=10
    3, -3, -12, 5, 2, -6, 5, -5, -9,
    -- filter=100 channel=11
    9, -7, 6, 7, -14, -12, 14, -7, -3,
    -- filter=100 channel=12
    7, -4, 6, -3, 8, -2, 3, -1, -4,
    -- filter=100 channel=13
    -9, 0, 12, -6, -8, 14, 1, -11, 9,
    -- filter=100 channel=14
    12, 13, -2, 9, -1, -5, -5, 0, 6,
    -- filter=100 channel=15
    -6, -20, 5, 9, -9, 18, 15, 1, 12,
    -- filter=100 channel=16
    7, -18, 4, -5, -5, 15, 1, -13, 0,
    -- filter=100 channel=17
    3, -7, -6, 19, -1, 3, 1, -4, -3,
    -- filter=100 channel=18
    -2, -3, 9, 0, -5, -4, -9, -4, 2,
    -- filter=100 channel=19
    6, 1, 0, -1, -1, -7, -5, -7, -11,
    -- filter=100 channel=20
    -3, 12, 16, -5, 9, 16, -7, -3, 0,
    -- filter=100 channel=21
    -9, 1, 2, -2, -3, -1, -4, -4, 4,
    -- filter=100 channel=22
    4, -9, 6, -1, 10, -8, -1, 9, -1,
    -- filter=100 channel=23
    8, 4, -5, 6, 0, -13, -1, 0, 1,
    -- filter=100 channel=24
    13, -8, 3, 5, 6, 0, 7, 4, 0,
    -- filter=100 channel=25
    -1, -16, 11, -3, -16, 13, 14, -1, 5,
    -- filter=100 channel=26
    7, -2, 6, -3, 2, 18, 8, -5, 0,
    -- filter=100 channel=27
    -2, -10, 9, 15, -3, 1, 18, -12, 1,
    -- filter=100 channel=28
    8, 1, 0, 9, -17, -6, 5, -2, -13,
    -- filter=100 channel=29
    -2, -13, 22, 0, -27, 22, -5, -16, 12,
    -- filter=100 channel=30
    22, 16, 14, 30, 9, 3, 18, 23, -4,
    -- filter=100 channel=31
    -8, 4, -2, 3, -2, 0, 0, -3, 10,
    -- filter=100 channel=32
    10, 8, -8, 0, -9, -2, 2, 4, -10,
    -- filter=100 channel=33
    -4, 2, -7, -6, -1, 0, -1, 1, -5,
    -- filter=100 channel=34
    -4, 11, 3, 0, 3, 1, 2, 2, 1,
    -- filter=100 channel=35
    2, -18, 0, 13, -5, -7, 19, -14, -2,
    -- filter=100 channel=36
    5, -1, -4, 0, 8, 5, -5, 1, 4,
    -- filter=100 channel=37
    -6, 2, 10, 13, 5, -2, 8, 0, 1,
    -- filter=100 channel=38
    3, -16, 3, 11, -5, 9, 16, -14, 5,
    -- filter=100 channel=39
    8, 6, 9, 5, 4, 4, 4, -2, -1,
    -- filter=100 channel=40
    -1, 1, 3, 2, 0, -1, -7, 6, -9,
    -- filter=100 channel=41
    13, -19, 0, 19, -22, 1, 0, -15, 3,
    -- filter=100 channel=42
    10, 9, 3, 6, 5, -8, -8, -2, 10,
    -- filter=100 channel=43
    3, 1, -2, -5, -6, -4, -8, -3, 0,
    -- filter=100 channel=44
    1, 0, 2, 13, -3, -11, 6, 10, -8,
    -- filter=100 channel=45
    -10, 9, 7, 8, 10, 7, 0, 10, 1,
    -- filter=100 channel=46
    8, -2, 11, -1, -4, 20, 7, -5, 20,
    -- filter=100 channel=47
    -9, 9, -4, -7, 4, -9, 8, -9, -5,
    -- filter=100 channel=48
    -5, -1, 16, -11, 4, 14, -6, -9, -5,
    -- filter=100 channel=49
    1, -8, 4, 4, -14, 0, -4, 4, -8,
    -- filter=100 channel=50
    15, 2, -9, 12, 3, 8, 4, 17, 8,
    -- filter=100 channel=51
    2, 0, -3, 4, -4, 4, 6, 0, 3,
    -- filter=100 channel=52
    -3, 3, -1, -5, -6, -5, 1, -7, -4,
    -- filter=100 channel=53
    7, 19, 0, 7, 5, -10, 13, 1, -6,
    -- filter=100 channel=54
    9, -11, 3, 8, 0, 0, 9, -4, -4,
    -- filter=100 channel=55
    -5, -9, 0, -10, -2, 5, -9, 0, 3,
    -- filter=100 channel=56
    3, 9, 11, -5, 1, 0, -8, 11, -4,
    -- filter=100 channel=57
    -3, -4, -6, 10, -3, 6, 9, -4, 0,
    -- filter=100 channel=58
    0, -5, 9, -7, 5, 10, -7, 7, -10,
    -- filter=100 channel=59
    -3, -1, 0, -4, -13, 9, 7, -15, 0,
    -- filter=100 channel=60
    -4, -15, 1, 15, -15, 8, 4, -4, 7,
    -- filter=100 channel=61
    15, -7, 3, 19, -12, -1, 5, -12, -9,
    -- filter=100 channel=62
    8, 1, 11, 15, -2, -5, 1, -6, -8,
    -- filter=100 channel=63
    5, -4, -10, -1, -6, -9, 4, 0, -2,
    -- filter=101 channel=0
    -8, 2, 3, 1, -5, 3, 16, 13, 14,
    -- filter=101 channel=1
    10, 7, -1, -7, -10, -14, -4, 3, 3,
    -- filter=101 channel=2
    -18, -10, -7, 3, 1, 11, 2, 0, 10,
    -- filter=101 channel=3
    5, -9, -13, -8, -3, 7, 0, 15, -2,
    -- filter=101 channel=4
    -4, -19, -10, -7, 0, 1, 10, 7, 9,
    -- filter=101 channel=5
    -4, 2, 0, -1, 10, -6, 6, 9, 14,
    -- filter=101 channel=6
    -4, -13, -17, -3, 0, -4, -1, -3, 3,
    -- filter=101 channel=7
    -4, 1, -11, 5, 6, -7, -6, 8, 4,
    -- filter=101 channel=8
    -18, -29, -24, -2, 3, 7, 15, 19, 14,
    -- filter=101 channel=9
    1, -3, 2, -4, 6, -7, 14, 9, 11,
    -- filter=101 channel=10
    -2, -5, -5, -9, 3, -3, -10, -8, -6,
    -- filter=101 channel=11
    3, -15, 0, 3, -19, -15, 0, 11, 14,
    -- filter=101 channel=12
    2, -1, 3, 0, -8, 9, 6, -2, 1,
    -- filter=101 channel=13
    -13, -4, 2, -8, -17, -17, 16, 17, 16,
    -- filter=101 channel=14
    1, -10, -8, 0, 6, 3, -6, -2, 3,
    -- filter=101 channel=15
    -22, -27, -23, 12, 13, 12, 6, 10, 11,
    -- filter=101 channel=16
    -18, -36, -15, -10, -14, 2, 21, 19, 22,
    -- filter=101 channel=17
    -15, -20, -14, 0, 5, -4, 5, 23, 20,
    -- filter=101 channel=18
    0, 0, -11, 4, 7, 15, 0, 4, 5,
    -- filter=101 channel=19
    10, -7, -8, -10, 4, -4, 0, -4, 6,
    -- filter=101 channel=20
    7, -5, 8, -2, 0, 0, 3, 8, 0,
    -- filter=101 channel=21
    0, 3, -4, 7, 11, 6, 0, -1, -3,
    -- filter=101 channel=22
    0, -4, 5, 5, -6, 10, -6, 1, 4,
    -- filter=101 channel=23
    -8, 5, 4, 1, -5, -1, -9, 7, 6,
    -- filter=101 channel=24
    10, -15, -15, -4, -11, -10, 4, 13, 18,
    -- filter=101 channel=25
    -13, -12, -21, -2, 3, -2, 17, 14, 10,
    -- filter=101 channel=26
    -8, -4, -4, 2, 0, 8, -1, -3, -3,
    -- filter=101 channel=27
    -14, -15, -27, -5, 0, 0, 19, 16, 9,
    -- filter=101 channel=28
    -20, -13, -14, -2, 1, -6, 1, 21, 18,
    -- filter=101 channel=29
    -17, -32, -18, 3, 6, -9, 20, 34, 33,
    -- filter=101 channel=30
    2, -8, -4, -4, -3, 0, -15, -12, 10,
    -- filter=101 channel=31
    8, -2, 1, 6, 8, -7, 3, 8, 0,
    -- filter=101 channel=32
    9, 2, 1, 1, 0, 5, -9, 3, -5,
    -- filter=101 channel=33
    3, 9, -6, -9, 3, 5, 4, -7, 9,
    -- filter=101 channel=34
    0, 2, 0, 3, 1, 7, 4, 8, -5,
    -- filter=101 channel=35
    -10, -6, -11, 0, -3, 3, -4, 0, 13,
    -- filter=101 channel=36
    -1, -3, 7, 8, 9, 7, 0, 3, 4,
    -- filter=101 channel=37
    0, -1, -1, 0, -6, 2, 4, 16, 0,
    -- filter=101 channel=38
    -3, -23, -20, -2, -18, -4, 4, 14, 20,
    -- filter=101 channel=39
    -3, 2, 2, 5, -1, 3, 8, -8, -1,
    -- filter=101 channel=40
    -4, 1, -11, 0, -4, -3, -5, -2, 8,
    -- filter=101 channel=41
    -29, -39, -30, 4, 5, 0, 30, 37, 32,
    -- filter=101 channel=42
    9, -4, 8, 3, 6, 10, -8, 0, 0,
    -- filter=101 channel=43
    16, 29, 39, 2, -2, 13, 21, 26, 30,
    -- filter=101 channel=44
    2, 8, -5, -5, 4, -4, 8, 1, 8,
    -- filter=101 channel=45
    -6, -9, -2, 4, -7, 10, -6, -1, 6,
    -- filter=101 channel=46
    -15, -12, -3, 7, 6, 0, 8, 6, 0,
    -- filter=101 channel=47
    -4, -8, 3, -2, -8, -6, -8, -4, 4,
    -- filter=101 channel=48
    -19, -12, 3, -3, -3, 0, 13, 0, 9,
    -- filter=101 channel=49
    -12, -5, -8, 20, 21, 20, 11, 13, 12,
    -- filter=101 channel=50
    10, 2, 1, 6, 0, -2, -3, 2, -1,
    -- filter=101 channel=51
    -6, 14, 10, -6, -6, 6, 5, 8, 5,
    -- filter=101 channel=52
    4, 2, 6, 4, 1, -10, -8, -5, -7,
    -- filter=101 channel=53
    12, 11, 6, -5, 5, -8, -4, -4, 5,
    -- filter=101 channel=54
    -15, -8, -12, 6, 5, 6, -4, 9, 15,
    -- filter=101 channel=55
    2, -8, 7, 2, -9, -9, -10, 8, 1,
    -- filter=101 channel=56
    3, -1, -8, -9, -6, 9, 3, 9, -5,
    -- filter=101 channel=57
    9, 6, -9, -7, 5, -6, 2, -5, 5,
    -- filter=101 channel=58
    4, 0, 7, -2, 3, 1, -6, -9, -11,
    -- filter=101 channel=59
    -7, -26, -15, 8, 8, -6, 5, 24, 9,
    -- filter=101 channel=60
    -24, -36, -28, 3, -6, -1, 34, 31, 33,
    -- filter=101 channel=61
    -17, -5, -3, -3, -2, -3, 4, 9, 29,
    -- filter=101 channel=62
    -11, -17, -7, 7, 3, 9, 13, 5, 19,
    -- filter=101 channel=63
    9, -4, -10, 9, 9, 1, 2, -1, -9,
    -- filter=102 channel=0
    8, 0, 6, 3, -5, 9, 0, 8, 6,
    -- filter=102 channel=1
    1, -9, 1, -7, -6, -3, 0, -10, 0,
    -- filter=102 channel=2
    9, 8, -6, 6, 0, -5, -5, -1, -6,
    -- filter=102 channel=3
    2, -10, 8, -8, -1, 2, -1, 0, 8,
    -- filter=102 channel=4
    -8, -2, 6, 6, -6, 1, 0, -1, 9,
    -- filter=102 channel=5
    -5, 0, 7, -5, 1, 8, 2, -5, -4,
    -- filter=102 channel=6
    -6, 4, -10, 10, -4, 3, 3, 0, -8,
    -- filter=102 channel=7
    -5, -7, 10, 1, -2, 8, -4, 0, 0,
    -- filter=102 channel=8
    -8, -9, 0, -9, -6, -4, -6, 0, -7,
    -- filter=102 channel=9
    -3, -1, -4, 4, 5, 4, 1, -4, -6,
    -- filter=102 channel=10
    0, -7, 7, 0, 5, 4, 2, 7, 2,
    -- filter=102 channel=11
    -6, -7, -2, 7, -8, 1, -4, 1, 5,
    -- filter=102 channel=12
    -1, 2, 2, -4, 8, 8, 1, -6, 10,
    -- filter=102 channel=13
    -5, 9, 8, 6, 10, -8, 6, 2, -5,
    -- filter=102 channel=14
    2, 0, -6, -7, -3, -4, -2, -10, -2,
    -- filter=102 channel=15
    2, 2, 4, 0, 6, 5, -4, -8, -2,
    -- filter=102 channel=16
    -6, 1, -1, 2, -4, -1, -9, -8, 5,
    -- filter=102 channel=17
    5, 0, 3, -7, 1, 2, 8, -7, 9,
    -- filter=102 channel=18
    -4, -5, -8, -4, -9, 3, 3, -9, 4,
    -- filter=102 channel=19
    -7, 9, 8, 7, -7, -2, -3, 0, -5,
    -- filter=102 channel=20
    -10, 9, 10, -6, -1, -4, 3, -8, 3,
    -- filter=102 channel=21
    -8, -7, 0, -4, -1, -1, 0, 7, -3,
    -- filter=102 channel=22
    3, -6, -5, 8, 9, -3, -7, -10, -1,
    -- filter=102 channel=23
    -5, 0, 3, 7, -6, -1, 5, 1, 9,
    -- filter=102 channel=24
    -3, 2, 10, 7, -10, -9, 3, 9, -3,
    -- filter=102 channel=25
    -7, -8, -10, 9, 4, 0, -3, -3, -2,
    -- filter=102 channel=26
    -3, -7, 0, 8, -6, 3, 5, 8, 7,
    -- filter=102 channel=27
    0, 1, -7, 7, -9, -2, 1, 9, -1,
    -- filter=102 channel=28
    -1, -8, -4, -7, 0, -4, -5, -2, -7,
    -- filter=102 channel=29
    -9, -4, -3, -7, 6, -10, -6, 0, -1,
    -- filter=102 channel=30
    -5, 0, 1, 0, -6, -5, -7, -3, -6,
    -- filter=102 channel=31
    8, -4, -10, 8, 5, 9, 8, -6, 3,
    -- filter=102 channel=32
    8, -7, 0, 7, -2, -3, 0, -5, 4,
    -- filter=102 channel=33
    8, -1, 0, 9, 0, -10, 0, -1, 6,
    -- filter=102 channel=34
    3, -10, -1, 5, 4, -4, 8, -8, -1,
    -- filter=102 channel=35
    0, 6, -4, -1, 10, 6, 0, -7, -2,
    -- filter=102 channel=36
    -6, -4, 0, -2, -4, 5, -4, 6, 0,
    -- filter=102 channel=37
    -8, 0, -7, 0, 7, 7, 1, -4, -8,
    -- filter=102 channel=38
    -4, 9, 7, -9, -5, 2, -1, -10, -7,
    -- filter=102 channel=39
    3, 0, -8, 5, -9, -2, -2, 7, 8,
    -- filter=102 channel=40
    8, 0, 0, 1, -5, 9, 0, -8, 0,
    -- filter=102 channel=41
    -5, -9, 6, 5, 1, 0, -7, 0, -6,
    -- filter=102 channel=42
    7, 3, 7, -1, 4, -5, -1, -2, 3,
    -- filter=102 channel=43
    -10, 7, 3, 7, 2, -4, -6, 0, 0,
    -- filter=102 channel=44
    -1, -3, -9, 0, 7, 1, -3, -3, 2,
    -- filter=102 channel=45
    -5, -7, 3, -6, 3, 1, -4, 5, -8,
    -- filter=102 channel=46
    7, 8, -10, -3, -3, -7, 6, 7, -3,
    -- filter=102 channel=47
    0, -2, -3, -1, -4, -8, -2, 0, 0,
    -- filter=102 channel=48
    -5, -10, 1, 10, -6, 1, 8, 0, 3,
    -- filter=102 channel=49
    7, 1, 9, -2, -5, -6, -4, -10, -7,
    -- filter=102 channel=50
    -6, 1, 7, -4, -1, -4, 6, -10, -2,
    -- filter=102 channel=51
    -8, -1, 1, -10, -4, -9, 4, 3, 10,
    -- filter=102 channel=52
    9, 6, 0, 5, 6, -6, -3, 4, -8,
    -- filter=102 channel=53
    -8, -8, -9, -3, -8, -7, 4, 3, 0,
    -- filter=102 channel=54
    1, -3, 9, -4, 9, 9, 1, 6, 5,
    -- filter=102 channel=55
    6, -5, -3, 9, -4, 6, -3, -8, -4,
    -- filter=102 channel=56
    -3, -5, 0, 0, 10, -10, 2, -10, -2,
    -- filter=102 channel=57
    0, -8, -4, -5, 6, -5, -9, -1, -7,
    -- filter=102 channel=58
    9, 4, -5, 0, 9, -2, 5, 0, -1,
    -- filter=102 channel=59
    -6, -4, -6, 1, -2, 8, -1, 1, -10,
    -- filter=102 channel=60
    -3, 0, 3, 10, -4, -6, 1, 3, 1,
    -- filter=102 channel=61
    -7, -3, -8, 10, 6, 7, 9, -2, -1,
    -- filter=102 channel=62
    3, 2, -8, 4, -8, 6, 8, -2, -4,
    -- filter=102 channel=63
    -3, -3, 1, 0, -9, 0, 0, -2, -9,
    -- filter=103 channel=0
    7, 22, 7, 4, 12, 10, 8, 5, 10,
    -- filter=103 channel=1
    -10, -2, 6, 0, 4, -3, -10, -7, -13,
    -- filter=103 channel=2
    -1, -1, 2, 0, -16, -15, -5, -14, -8,
    -- filter=103 channel=3
    -7, 7, 4, 2, -14, -9, -3, -12, 2,
    -- filter=103 channel=4
    0, 8, 14, -4, 17, 13, -5, -3, 6,
    -- filter=103 channel=5
    -16, -14, -11, -11, -19, -10, -2, -6, 3,
    -- filter=103 channel=6
    11, 3, 7, 0, -1, -2, -10, -4, 2,
    -- filter=103 channel=7
    -5, -15, 5, -7, -5, 6, -9, -7, 6,
    -- filter=103 channel=8
    22, 28, 17, 2, 0, 12, 3, 5, -11,
    -- filter=103 channel=9
    -21, -36, -42, -28, -35, -44, -14, -44, -43,
    -- filter=103 channel=10
    9, 21, 0, 7, 12, 17, -6, 25, 9,
    -- filter=103 channel=11
    -4, 11, 20, 10, 0, 15, 2, -5, -5,
    -- filter=103 channel=12
    8, -6, 1, 4, -7, -1, -8, -6, -5,
    -- filter=103 channel=13
    15, 13, 6, 3, 1, -5, 1, 1, -11,
    -- filter=103 channel=14
    -5, -4, 7, 0, -13, -1, -5, -15, -10,
    -- filter=103 channel=15
    4, 5, 10, 0, -5, 14, -3, 2, -15,
    -- filter=103 channel=16
    19, 16, 8, -1, -4, -16, -3, -25, -16,
    -- filter=103 channel=17
    0, 11, 22, -8, 7, -1, 4, 3, -4,
    -- filter=103 channel=18
    11, 5, 0, 12, 3, 0, 4, 9, -9,
    -- filter=103 channel=19
    -19, -28, -11, -10, -24, -15, -1, -26, -6,
    -- filter=103 channel=20
    -9, -21, -17, -20, -16, -19, -17, -13, -18,
    -- filter=103 channel=21
    0, -5, 0, 4, -2, -1, 0, -5, 11,
    -- filter=103 channel=22
    -2, 4, 0, 1, -9, 1, -6, 5, -1,
    -- filter=103 channel=23
    4, 8, 7, 20, 20, 32, -1, 22, 9,
    -- filter=103 channel=24
    13, 9, 16, 8, 14, 16, -11, -3, -1,
    -- filter=103 channel=25
    0, -4, 0, -18, -8, -6, -1, -11, -6,
    -- filter=103 channel=26
    -10, -17, -12, -14, 3, -7, -2, -16, 4,
    -- filter=103 channel=27
    5, 25, 18, -7, 14, 3, 4, 1, 6,
    -- filter=103 channel=28
    0, 5, 3, 5, -18, -9, -13, -17, -16,
    -- filter=103 channel=29
    5, 11, -4, -20, -7, -12, -12, -21, -21,
    -- filter=103 channel=30
    -21, -13, -1, -34, -34, 0, -24, -26, -4,
    -- filter=103 channel=31
    -5, 1, 0, 1, 3, -4, 0, 12, -5,
    -- filter=103 channel=32
    -5, -7, 13, -5, -7, 9, -11, 3, 15,
    -- filter=103 channel=33
    4, -10, -9, -10, 1, -4, 3, -5, 7,
    -- filter=103 channel=34
    -9, -1, 1, -6, -7, 6, -15, -15, -13,
    -- filter=103 channel=35
    9, 28, 15, 12, 21, 29, 3, 21, 21,
    -- filter=103 channel=36
    -4, -7, 5, 6, 7, 9, 11, 10, 13,
    -- filter=103 channel=37
    -12, -8, -1, -18, -17, 0, -16, -10, -14,
    -- filter=103 channel=38
    20, 16, 7, 13, 20, 15, 6, 10, -11,
    -- filter=103 channel=39
    -8, 9, 0, 0, 1, 10, 9, -5, 8,
    -- filter=103 channel=40
    -6, -5, -5, 0, 4, -6, 2, 9, -2,
    -- filter=103 channel=41
    23, 11, 12, -10, 5, 3, -9, -2, -11,
    -- filter=103 channel=42
    7, 6, 4, 5, 2, 9, -2, 8, -1,
    -- filter=103 channel=43
    -1, 0, 5, 4, 6, 12, -10, -13, 6,
    -- filter=103 channel=44
    -5, 1, -10, -1, -9, -1, -1, -1, 4,
    -- filter=103 channel=45
    -9, -1, -8, 2, -6, 3, -8, -10, -10,
    -- filter=103 channel=46
    -7, -12, -13, -17, -9, 0, -6, -16, -12,
    -- filter=103 channel=47
    -2, 7, 9, -3, 2, -6, 2, 1, -4,
    -- filter=103 channel=48
    -7, 1, -8, -11, -6, -15, 4, -12, -6,
    -- filter=103 channel=49
    5, 27, 25, 12, 12, 16, 14, 18, 16,
    -- filter=103 channel=50
    -7, -21, -6, -12, -12, 0, -23, -18, 3,
    -- filter=103 channel=51
    7, 22, 13, 8, 31, 16, 13, 30, 10,
    -- filter=103 channel=52
    -2, 1, 5, -8, 6, 5, 0, 4, 1,
    -- filter=103 channel=53
    -12, -22, 3, -21, -5, 0, -16, -17, 2,
    -- filter=103 channel=54
    -17, -28, -30, -13, -30, -37, -12, -24, -24,
    -- filter=103 channel=55
    -5, 7, -4, -9, -7, 4, -9, 1, 7,
    -- filter=103 channel=56
    -10, -3, 1, -2, -5, -7, -12, 4, -4,
    -- filter=103 channel=57
    -10, -7, -8, 5, -2, -6, 5, 3, 7,
    -- filter=103 channel=58
    1, 6, -7, 0, -9, 3, 5, -3, 4,
    -- filter=103 channel=59
    -2, 19, 14, 2, -2, 9, 0, -6, -4,
    -- filter=103 channel=60
    21, 36, 16, 2, 12, 14, -8, 7, 0,
    -- filter=103 channel=61
    5, 29, 20, 20, 19, 24, -3, 9, 4,
    -- filter=103 channel=62
    -4, -5, 6, 1, -10, -3, -6, -1, -16,
    -- filter=103 channel=63
    -2, 8, -6, -10, -9, -7, -1, -8, 0,
    -- filter=104 channel=0
    0, 16, 5, 16, 6, 6, 10, 12, 20,
    -- filter=104 channel=1
    -10, -6, -4, -2, -17, -3, -2, -15, -13,
    -- filter=104 channel=2
    -12, -20, -7, -15, -16, -12, -18, -17, -18,
    -- filter=104 channel=3
    -15, -10, -14, -4, 2, -7, -2, -1, -12,
    -- filter=104 channel=4
    6, 6, 10, 11, 19, 9, 11, 16, 17,
    -- filter=104 channel=5
    3, -11, -4, 8, -2, -7, -9, 2, -6,
    -- filter=104 channel=6
    -10, -6, 2, -2, 2, -4, 1, -1, -7,
    -- filter=104 channel=7
    -5, 5, 1, 2, -15, 0, -9, -5, 8,
    -- filter=104 channel=8
    7, 6, -3, 9, 25, 17, 7, 18, 18,
    -- filter=104 channel=9
    -2, -15, -18, -1, -26, -34, -4, -10, -14,
    -- filter=104 channel=10
    5, 4, 0, 3, 16, 10, -2, 6, 0,
    -- filter=104 channel=11
    7, 0, 0, 0, 12, 11, -6, 8, 8,
    -- filter=104 channel=12
    6, -2, -2, 5, -10, -2, 1, -7, 9,
    -- filter=104 channel=13
    -1, 17, 4, 13, 3, -1, 18, 5, -2,
    -- filter=104 channel=14
    -3, 3, 6, -14, 2, -9, -2, -2, 0,
    -- filter=104 channel=15
    12, 3, 0, 16, 20, 13, 14, 9, -2,
    -- filter=104 channel=16
    0, 0, -13, -3, -6, -7, -5, 9, -18,
    -- filter=104 channel=17
    13, 12, 7, 13, 1, 16, 14, 8, 16,
    -- filter=104 channel=18
    7, 13, 13, 12, 17, 20, 15, 22, 3,
    -- filter=104 channel=19
    -9, -9, -8, -20, -11, -23, -13, -22, -7,
    -- filter=104 channel=20
    -10, -5, -16, -13, -3, -13, -14, -15, -18,
    -- filter=104 channel=21
    -3, -8, 10, 2, -11, 6, -1, -5, 4,
    -- filter=104 channel=22
    -9, 4, 2, -8, 1, 9, 9, 5, 4,
    -- filter=104 channel=23
    3, 2, 12, 0, 15, 17, 0, 0, 5,
    -- filter=104 channel=24
    -2, 7, 0, 12, 4, 14, 10, 18, 19,
    -- filter=104 channel=25
    -12, -16, -21, -16, -21, -25, -13, -25, -22,
    -- filter=104 channel=26
    -18, -16, 1, -22, -4, -6, -17, -20, -14,
    -- filter=104 channel=27
    5, -10, -12, -10, 6, -5, -1, 0, 7,
    -- filter=104 channel=28
    3, 11, 11, -2, 5, -3, 2, 13, 3,
    -- filter=104 channel=29
    1, 0, -13, -3, -12, -9, 2, 1, -1,
    -- filter=104 channel=30
    -13, -29, -12, -33, -34, -5, -33, -18, -6,
    -- filter=104 channel=31
    -7, 10, 5, -4, 0, 11, -6, 5, 1,
    -- filter=104 channel=32
    -18, -15, -3, -23, -6, -4, -12, -17, -2,
    -- filter=104 channel=33
    10, -8, 5, 1, -9, 8, 9, -7, -3,
    -- filter=104 channel=34
    0, -2, -4, -10, -7, -5, 2, 2, 2,
    -- filter=104 channel=35
    -8, -4, 1, -15, 8, 13, -16, -8, -2,
    -- filter=104 channel=36
    0, -7, -4, 7, -5, -3, -2, -9, -7,
    -- filter=104 channel=37
    -12, -3, 0, 2, -7, -20, -11, -5, 0,
    -- filter=104 channel=38
    0, -2, 4, 0, -1, 8, 0, 10, 0,
    -- filter=104 channel=39
    1, 4, -8, 0, -9, -9, 4, -5, 8,
    -- filter=104 channel=40
    -12, -12, 6, -10, -8, -11, 1, -12, -5,
    -- filter=104 channel=41
    -4, 0, -8, 0, 12, -5, 6, 15, 13,
    -- filter=104 channel=42
    8, -6, 8, -7, -4, -7, -3, -5, -4,
    -- filter=104 channel=43
    -32, -29, -20, -20, -22, -25, -28, -18, -15,
    -- filter=104 channel=44
    -17, -6, 0, -20, -23, -11, -9, -25, -16,
    -- filter=104 channel=45
    -7, -7, -10, 5, 3, 0, -6, 3, -6,
    -- filter=104 channel=46
    -7, -3, -3, 3, -15, -10, 2, -14, -6,
    -- filter=104 channel=47
    -7, 2, -1, 3, -6, -4, -6, -2, 3,
    -- filter=104 channel=48
    -4, -6, 4, 7, 4, -6, 3, 8, 0,
    -- filter=104 channel=49
    -2, 5, 16, 15, 16, 20, 12, 18, 20,
    -- filter=104 channel=50
    -14, -6, -10, -13, -12, -2, -4, -10, -8,
    -- filter=104 channel=51
    18, 28, 10, 14, 32, 28, 16, 12, 8,
    -- filter=104 channel=52
    4, 4, -3, 5, 1, 0, 8, -4, 0,
    -- filter=104 channel=53
    -14, -14, -7, -24, -18, -9, -27, -18, -1,
    -- filter=104 channel=54
    -18, -6, -15, -5, -25, -18, -10, -20, -24,
    -- filter=104 channel=55
    -3, 7, 5, 10, 5, 3, 5, 4, -9,
    -- filter=104 channel=56
    -10, 1, -2, 6, 3, -8, -5, -5, -4,
    -- filter=104 channel=57
    -4, -3, -10, 10, 5, 9, 0, -8, -9,
    -- filter=104 channel=58
    0, -5, -8, -5, -8, 4, -8, 0, 4,
    -- filter=104 channel=59
    -1, -3, 3, -11, 0, 0, 2, -12, -3,
    -- filter=104 channel=60
    11, 22, 13, 18, 20, 4, 11, 29, 18,
    -- filter=104 channel=61
    6, 9, 10, 19, 29, 16, 8, 20, 24,
    -- filter=104 channel=62
    2, 0, 1, 7, -15, 2, -1, 0, -10,
    -- filter=104 channel=63
    -1, 0, 6, 0, -7, -2, 3, 1, 0,
    -- filter=105 channel=0
    -9, -13, -15, 7, -9, 2, -9, 6, -4,
    -- filter=105 channel=1
    -9, -4, -4, 5, 4, -11, -6, -11, -8,
    -- filter=105 channel=2
    4, -11, 0, -7, 2, 0, -8, 1, -8,
    -- filter=105 channel=3
    -3, -6, 14, -4, 7, 8, -2, 8, -1,
    -- filter=105 channel=4
    -3, -5, 4, 9, -6, -7, -6, -7, -9,
    -- filter=105 channel=5
    7, 4, 10, 1, 0, 10, 11, -2, 4,
    -- filter=105 channel=6
    -5, 11, 3, 1, -8, -12, -9, -6, -9,
    -- filter=105 channel=7
    -6, -3, -3, 8, 3, -2, 6, 8, 3,
    -- filter=105 channel=8
    5, -9, -7, 5, -2, 3, -12, -13, -9,
    -- filter=105 channel=9
    14, 47, 40, 25, 49, 48, 10, 31, 46,
    -- filter=105 channel=10
    0, -2, -9, 1, 0, -9, -5, 4, 2,
    -- filter=105 channel=11
    -2, 0, -1, 7, -9, -1, -3, -6, -3,
    -- filter=105 channel=12
    -2, -3, 2, -4, 0, -4, 8, 11, 8,
    -- filter=105 channel=13
    -8, 8, 14, -2, 0, 6, 6, -2, -2,
    -- filter=105 channel=14
    9, 5, 10, 11, -8, 6, 7, -1, -9,
    -- filter=105 channel=15
    -2, 14, -3, 10, -4, 6, -1, -9, -10,
    -- filter=105 channel=16
    3, 9, 7, -4, 9, 3, -14, 6, -17,
    -- filter=105 channel=17
    -6, -9, -3, -1, -3, 0, 10, 4, -2,
    -- filter=105 channel=18
    11, 22, 18, 19, 14, 7, 16, 14, 0,
    -- filter=105 channel=19
    0, 8, -1, 0, 14, 0, 9, 7, 2,
    -- filter=105 channel=20
    11, 17, 9, 2, 18, 10, 11, 23, 8,
    -- filter=105 channel=21
    11, 11, 2, 2, 11, 5, -4, 12, -2,
    -- filter=105 channel=22
    6, 5, 4, -9, -4, 0, 4, 5, 7,
    -- filter=105 channel=23
    -12, -18, -8, -1, -17, -12, 0, -15, -12,
    -- filter=105 channel=24
    -1, 5, 0, 7, 4, 0, 8, 7, 7,
    -- filter=105 channel=25
    -15, -4, -2, -10, -8, -22, -3, -3, -11,
    -- filter=105 channel=26
    9, 11, -10, 4, -9, -3, 6, 2, -3,
    -- filter=105 channel=27
    -15, -4, -15, -9, -12, -20, -15, -16, -12,
    -- filter=105 channel=28
    12, 14, 15, 6, 21, 4, 8, 14, 12,
    -- filter=105 channel=29
    -4, 16, 8, 6, 20, 8, 1, 12, 0,
    -- filter=105 channel=30
    0, 0, -1, 6, 0, -7, 7, 1, 0,
    -- filter=105 channel=31
    11, 1, -2, 9, -1, 0, 8, 11, 13,
    -- filter=105 channel=32
    -4, -3, -3, 6, -7, 7, 11, 0, -7,
    -- filter=105 channel=33
    4, 6, 5, 2, 9, -6, -10, 9, -9,
    -- filter=105 channel=34
    8, -5, -1, 0, -6, -3, 0, 4, -8,
    -- filter=105 channel=35
    1, -19, -24, -6, -24, -18, -14, -17, -12,
    -- filter=105 channel=36
    -3, 8, 5, -7, -3, 9, -2, 7, 1,
    -- filter=105 channel=37
    -5, -1, 2, 3, 2, 9, 9, 6, 13,
    -- filter=105 channel=38
    0, -17, -2, 1, -17, -9, -15, -7, -22,
    -- filter=105 channel=39
    -3, 3, 0, 7, 10, 3, 7, 0, -7,
    -- filter=105 channel=40
    6, -8, 6, 7, -6, -5, -4, -1, 0,
    -- filter=105 channel=41
    -1, 6, 0, -3, -3, -11, 6, -11, -20,
    -- filter=105 channel=42
    -1, 8, -2, 9, 10, 8, 7, -10, 3,
    -- filter=105 channel=43
    -20, -4, 1, -12, -7, 5, 0, -1, -13,
    -- filter=105 channel=44
    -3, -2, -2, 0, -12, -1, 6, -10, 1,
    -- filter=105 channel=45
    2, 0, 1, -6, 0, -3, 8, -8, 0,
    -- filter=105 channel=46
    -5, 0, -1, 12, 6, -5, 0, 7, -5,
    -- filter=105 channel=47
    8, -6, -1, -1, 7, -9, 5, 10, -2,
    -- filter=105 channel=48
    -4, -2, -1, 10, 7, 1, -7, 4, 8,
    -- filter=105 channel=49
    5, 5, -3, 6, 1, -2, 0, 1, -14,
    -- filter=105 channel=50
    -3, 8, -4, 0, 1, 14, 14, 10, 10,
    -- filter=105 channel=51
    14, 1, -9, -5, -4, 5, -4, -4, 0,
    -- filter=105 channel=52
    -4, -3, -1, -8, 10, 3, 3, -2, -7,
    -- filter=105 channel=53
    5, 1, -12, 6, 0, -3, 7, -7, 0,
    -- filter=105 channel=54
    13, 35, 29, 27, 37, 25, 18, 14, 15,
    -- filter=105 channel=55
    1, -7, -10, 0, 7, 1, -10, 8, 0,
    -- filter=105 channel=56
    5, -3, -2, 3, -2, 5, -9, -5, -1,
    -- filter=105 channel=57
    -4, 0, 0, 4, 5, -5, -1, -1, -9,
    -- filter=105 channel=58
    9, 8, -3, 7, 9, 6, 9, 17, 11,
    -- filter=105 channel=59
    -3, 9, 12, -6, 6, -7, -3, 0, -8,
    -- filter=105 channel=60
    -5, -8, 6, 9, -5, -2, -6, -3, -19,
    -- filter=105 channel=61
    7, -7, -5, -2, -1, -12, 2, 1, -13,
    -- filter=105 channel=62
    0, 6, 8, 4, -7, -3, 3, 5, 6,
    -- filter=105 channel=63
    -5, -8, 7, 4, -9, 3, -6, 8, 9,
    -- filter=106 channel=0
    5, 0, 7, 0, -5, -6, -7, 1, -7,
    -- filter=106 channel=1
    14, 3, 2, 13, -1, 1, -4, -3, 4,
    -- filter=106 channel=2
    2, -4, -5, 9, -8, -12, -6, 2, -9,
    -- filter=106 channel=3
    1, -12, 5, -11, -8, 5, 2, -12, 0,
    -- filter=106 channel=4
    9, -7, 10, 2, 1, 6, 8, -3, 5,
    -- filter=106 channel=5
    0, 9, -6, -3, 12, -6, 12, -5, -5,
    -- filter=106 channel=6
    2, 9, 5, 3, 3, 7, 5, 10, 9,
    -- filter=106 channel=7
    -1, -6, 1, -4, 4, 0, 12, 11, 4,
    -- filter=106 channel=8
    -2, 0, 0, -5, 6, -6, 11, 3, -8,
    -- filter=106 channel=9
    13, 12, 7, 21, 18, 30, 7, 10, 23,
    -- filter=106 channel=10
    10, 0, 6, 8, 0, 0, 0, -4, -6,
    -- filter=106 channel=11
    -1, -4, 0, 6, 5, -7, 0, 1, -4,
    -- filter=106 channel=12
    10, -9, 9, 1, 10, 0, 0, 10, 3,
    -- filter=106 channel=13
    -2, 5, -4, -8, 3, 14, 2, 0, -3,
    -- filter=106 channel=14
    -4, 1, 4, 10, -5, -9, -2, -7, -7,
    -- filter=106 channel=15
    0, 0, 9, 2, -2, 3, 10, 7, 0,
    -- filter=106 channel=16
    -7, -12, -7, 6, -8, -4, 12, -10, -6,
    -- filter=106 channel=17
    11, 2, -7, 0, 8, -3, 8, -6, -5,
    -- filter=106 channel=18
    6, 9, 17, 2, 5, 7, 16, 17, 6,
    -- filter=106 channel=19
    14, -4, 6, 13, 9, 0, 7, 4, 0,
    -- filter=106 channel=20
    8, 1, -5, -2, 5, 7, -7, 6, -5,
    -- filter=106 channel=21
    -8, 5, -3, 4, -8, 7, -2, 6, 5,
    -- filter=106 channel=22
    -10, 0, -2, -5, -7, 0, 3, -10, -5,
    -- filter=106 channel=23
    10, -3, 4, -8, -4, -5, 13, 7, -5,
    -- filter=106 channel=24
    6, -9, -5, 12, -8, 6, -4, -5, -2,
    -- filter=106 channel=25
    1, -11, -10, 9, -10, 4, -1, -3, -1,
    -- filter=106 channel=26
    -3, -6, 0, 0, 5, -5, 8, 3, -2,
    -- filter=106 channel=27
    8, -6, 0, -6, -14, 0, 5, -9, -10,
    -- filter=106 channel=28
    3, 0, 7, 15, 16, 9, 11, -5, 2,
    -- filter=106 channel=29
    -8, 1, 2, 11, 6, -4, 10, 4, -13,
    -- filter=106 channel=30
    0, 2, -12, 7, 4, -6, 12, 5, 3,
    -- filter=106 channel=31
    7, 3, -4, -1, 10, -1, -1, 9, 6,
    -- filter=106 channel=32
    -2, -10, -7, 7, -1, 3, 3, -4, 2,
    -- filter=106 channel=33
    2, -8, -5, 5, -1, -5, 3, 7, 4,
    -- filter=106 channel=34
    -6, 0, -9, -2, -6, -8, 9, 2, 6,
    -- filter=106 channel=35
    3, -2, -6, -5, 0, -6, 7, -2, -17,
    -- filter=106 channel=36
    -1, 10, 10, 7, -7, -3, -7, -4, 1,
    -- filter=106 channel=37
    2, -3, -8, -1, 6, 2, 7, -3, -1,
    -- filter=106 channel=38
    5, -8, -4, 1, -15, -2, -4, -14, -6,
    -- filter=106 channel=39
    0, 0, 5, 2, -1, -7, 0, -2, -8,
    -- filter=106 channel=40
    -8, 2, 2, -5, 1, 3, -10, 7, -2,
    -- filter=106 channel=41
    -7, 0, 3, 11, -1, -4, -5, -15, -15,
    -- filter=106 channel=42
    9, 0, 0, -9, 10, 4, -2, -1, 9,
    -- filter=106 channel=43
    5, -3, 5, 0, -12, -5, 8, 5, -2,
    -- filter=106 channel=44
    -3, 7, -5, -5, 2, -2, 13, 4, 1,
    -- filter=106 channel=45
    7, -5, 0, 4, 0, -6, 4, 3, -5,
    -- filter=106 channel=46
    -4, 1, -5, 7, 2, -6, 6, -1, -9,
    -- filter=106 channel=47
    0, -5, -9, -10, 4, -4, -6, 2, -8,
    -- filter=106 channel=48
    -3, -2, -8, 1, -6, 11, -9, 6, 7,
    -- filter=106 channel=49
    11, 4, -7, -2, -5, 6, -5, 9, 5,
    -- filter=106 channel=50
    11, 8, 8, -4, 12, -3, 2, 0, 2,
    -- filter=106 channel=51
    11, 0, -4, 7, 8, -3, 0, -6, 0,
    -- filter=106 channel=52
    10, -7, -3, 5, 9, 0, 1, 1, -1,
    -- filter=106 channel=53
    1, 4, -9, 6, 7, -14, 5, -8, -12,
    -- filter=106 channel=54
    12, 0, 16, 14, 17, 9, 14, 7, 0,
    -- filter=106 channel=55
    -6, -9, -10, -9, -7, -2, -8, -9, 8,
    -- filter=106 channel=56
    -8, 0, 2, -8, 3, 3, 8, 0, 9,
    -- filter=106 channel=57
    7, -9, 5, 6, 8, 9, 6, -2, -6,
    -- filter=106 channel=58
    9, 6, 1, 5, 2, -2, 0, 15, 10,
    -- filter=106 channel=59
    2, -13, -1, -11, -4, -4, -2, -4, -11,
    -- filter=106 channel=60
    2, -6, 7, 0, 0, -2, 4, -15, -4,
    -- filter=106 channel=61
    13, -7, -3, 0, -5, 0, 12, -3, 1,
    -- filter=106 channel=62
    7, -13, -7, 7, 7, -1, -4, -13, -3,
    -- filter=106 channel=63
    -5, 10, 8, 0, 10, -3, 3, -3, -9,
    -- filter=107 channel=0
    -5, -15, -15, -9, 0, -16, -2, -18, 2,
    -- filter=107 channel=1
    -4, 10, 16, 12, 15, 26, 9, 8, 23,
    -- filter=107 channel=2
    5, 18, 23, 11, 11, 24, 15, 5, 17,
    -- filter=107 channel=3
    7, 4, 9, 8, 14, 10, -5, 6, 8,
    -- filter=107 channel=4
    -10, 0, -12, 3, -4, -13, -1, -16, -4,
    -- filter=107 channel=5
    -5, -3, 15, -6, 1, 9, -6, 4, -4,
    -- filter=107 channel=6
    0, 12, 3, 7, 10, 14, 8, 3, 1,
    -- filter=107 channel=7
    1, -7, 7, -3, -4, 7, 9, 4, 4,
    -- filter=107 channel=8
    -12, 0, -3, -16, -11, -9, -6, -18, -4,
    -- filter=107 channel=9
    17, 43, 39, 19, 46, 57, 10, 39, 45,
    -- filter=107 channel=10
    5, 3, 0, 1, 6, -3, 12, -4, 3,
    -- filter=107 channel=11
    2, 0, 6, -4, 0, -4, -2, 2, 1,
    -- filter=107 channel=12
    -7, -3, 7, 8, 0, -1, -5, 0, 4,
    -- filter=107 channel=13
    -7, 3, 3, -3, -4, 6, 0, 5, -7,
    -- filter=107 channel=14
    7, -4, 5, 0, -3, 4, 10, 2, -9,
    -- filter=107 channel=15
    -13, -2, 2, -8, -9, 2, -3, -6, 0,
    -- filter=107 channel=16
    -11, 9, 17, -13, 11, 16, 4, 1, 11,
    -- filter=107 channel=17
    -8, 0, -10, -7, -6, -12, -3, -12, -10,
    -- filter=107 channel=18
    -6, -3, 9, 7, 3, 3, 0, 0, 2,
    -- filter=107 channel=19
    9, 11, 7, 4, 33, 19, 20, 15, 13,
    -- filter=107 channel=20
    14, 5, 7, 7, 27, 21, 20, 8, 11,
    -- filter=107 channel=21
    -2, 0, 0, 2, 4, 3, 1, -6, 10,
    -- filter=107 channel=22
    0, -6, 1, 5, 2, 0, 0, 9, -5,
    -- filter=107 channel=23
    8, 0, -7, 1, -10, -4, -1, 4, 0,
    -- filter=107 channel=24
    -10, -6, -9, -19, -17, -4, -8, 0, -6,
    -- filter=107 channel=25
    -3, 4, 28, 6, 23, 27, 18, 22, 12,
    -- filter=107 channel=26
    8, 13, 16, 10, 0, 0, 4, 7, 17,
    -- filter=107 channel=27
    -2, -7, -6, -5, 0, 10, 0, 4, 8,
    -- filter=107 channel=28
    10, 0, 8, -1, 2, 12, -10, 6, 3,
    -- filter=107 channel=29
    1, 17, 6, 6, 19, 10, -6, -4, 7,
    -- filter=107 channel=30
    12, 4, 5, 10, 3, 18, 3, 21, 12,
    -- filter=107 channel=31
    9, 0, -8, -1, -4, -5, 2, 4, 8,
    -- filter=107 channel=32
    15, 7, 8, 10, 14, 7, 6, 6, 12,
    -- filter=107 channel=33
    10, -5, 0, 9, 0, -9, 2, 2, -8,
    -- filter=107 channel=34
    0, 5, 4, 11, 10, 2, -5, -8, -2,
    -- filter=107 channel=35
    -6, -12, -4, -15, -10, -9, 4, -6, 0,
    -- filter=107 channel=36
    1, 11, 6, 0, -9, 1, 11, -4, 7,
    -- filter=107 channel=37
    -2, 12, 14, 8, 18, 16, -2, 11, 17,
    -- filter=107 channel=38
    3, 4, 6, -12, 1, 4, 0, -7, 4,
    -- filter=107 channel=39
    -5, 6, -1, 1, 0, 6, 6, 6, -2,
    -- filter=107 channel=40
    -3, -5, -8, 6, 0, 2, 10, 2, 2,
    -- filter=107 channel=41
    -17, -11, 1, -11, -14, -2, 2, -5, -19,
    -- filter=107 channel=42
    9, 3, -9, -10, -8, 0, -6, -6, 0,
    -- filter=107 channel=43
    16, 9, 16, 12, 20, 15, 17, 19, 1,
    -- filter=107 channel=44
    -2, 5, 21, 6, 18, 9, 11, 20, 6,
    -- filter=107 channel=45
    -7, -1, 5, -1, 10, -5, -9, -2, 8,
    -- filter=107 channel=46
    10, 2, 15, 3, 8, 9, 2, 13, 13,
    -- filter=107 channel=47
    4, -3, 0, -7, -4, -5, 2, 0, 4,
    -- filter=107 channel=48
    5, 3, 12, 4, 2, 0, 8, 10, 7,
    -- filter=107 channel=49
    -6, -2, -14, -1, -8, -16, -10, -5, 1,
    -- filter=107 channel=50
    11, 4, 3, 5, 6, 9, 21, 6, 11,
    -- filter=107 channel=51
    -4, -16, -11, -16, -14, -10, 1, -9, -13,
    -- filter=107 channel=52
    2, 6, 8, 0, 10, -8, -4, 5, 2,
    -- filter=107 channel=53
    5, 5, 15, 2, 14, 18, 14, 0, 9,
    -- filter=107 channel=54
    11, 35, 19, 16, 22, 26, -1, 19, 26,
    -- filter=107 channel=55
    0, -7, -7, -9, 8, -5, 4, 1, 10,
    -- filter=107 channel=56
    -5, -7, 12, 3, 2, -3, -3, 8, -3,
    -- filter=107 channel=57
    -1, 7, -4, -2, -3, 1, 1, 3, 3,
    -- filter=107 channel=58
    8, 2, 11, 5, 9, 13, 17, 13, 18,
    -- filter=107 channel=59
    1, -4, 10, -2, 7, 10, -6, -8, 2,
    -- filter=107 channel=60
    -12, -21, -15, -19, -17, -16, -5, -13, -18,
    -- filter=107 channel=61
    -22, -28, -11, -14, -24, -14, -9, -24, -13,
    -- filter=107 channel=62
    -2, -3, 1, 1, 6, 14, -4, 1, -1,
    -- filter=107 channel=63
    -9, -6, -2, 4, 0, -4, -7, 5, 0,
    -- filter=108 channel=0
    6, -4, -7, 7, -13, 0, 0, -3, -5,
    -- filter=108 channel=1
    0, 7, 8, 3, 5, -3, -5, 7, 2,
    -- filter=108 channel=2
    3, 1, -11, 0, -9, -12, -1, -3, 4,
    -- filter=108 channel=3
    10, 4, 10, 6, -4, 4, 1, -1, 0,
    -- filter=108 channel=4
    6, -2, -2, 11, 1, -13, 0, -7, -4,
    -- filter=108 channel=5
    0, 4, -7, -6, 8, -8, -6, 13, -1,
    -- filter=108 channel=6
    -7, -9, 7, 7, -12, 9, -8, -10, -5,
    -- filter=108 channel=7
    1, -5, 0, -4, 13, -9, 8, -3, 9,
    -- filter=108 channel=8
    16, -1, -10, 18, -14, -4, 0, -10, -1,
    -- filter=108 channel=9
    19, 0, 4, 11, 2, 16, -1, -2, 4,
    -- filter=108 channel=10
    0, 9, 4, 4, 0, 9, 5, 12, 8,
    -- filter=108 channel=11
    7, -3, -12, 16, 11, -15, 4, 1, -13,
    -- filter=108 channel=12
    -9, 7, -3, -5, 6, -8, -8, -7, 9,
    -- filter=108 channel=13
    10, -2, 4, 3, -18, -6, -6, 2, -7,
    -- filter=108 channel=14
    0, 13, -2, -6, 2, 7, 13, 14, 9,
    -- filter=108 channel=15
    9, 2, -6, 11, -18, -1, 10, -13, 1,
    -- filter=108 channel=16
    0, -3, -18, 0, 1, -9, 12, -4, -14,
    -- filter=108 channel=17
    3, -7, -15, -1, -6, -9, -3, -5, -14,
    -- filter=108 channel=18
    10, 5, -7, 7, 3, -2, -7, -9, -4,
    -- filter=108 channel=19
    -8, 0, -3, -8, 13, -6, 8, 8, -14,
    -- filter=108 channel=20
    -6, -9, 8, 6, -11, 7, 2, -6, 5,
    -- filter=108 channel=21
    2, 0, 0, 0, 0, 0, -4, -9, 3,
    -- filter=108 channel=22
    -9, -9, -3, -2, 4, 7, 0, 8, -6,
    -- filter=108 channel=23
    5, 4, -8, 5, 13, -4, -4, 2, 11,
    -- filter=108 channel=24
    11, -5, -7, -2, -2, -4, 8, -10, -6,
    -- filter=108 channel=25
    12, 5, 0, 4, 10, -9, 0, -6, 5,
    -- filter=108 channel=26
    12, -7, -1, 10, 8, 0, -1, 12, 3,
    -- filter=108 channel=27
    -2, -2, 4, 16, 1, -9, 7, 9, 10,
    -- filter=108 channel=28
    5, 0, -9, 0, -4, -12, -7, 2, -19,
    -- filter=108 channel=29
    10, -19, 0, 10, -8, -19, -1, -5, -14,
    -- filter=108 channel=30
    17, 11, -1, 20, 27, 6, 12, 9, 9,
    -- filter=108 channel=31
    -8, 3, 11, -5, 8, -1, 7, 1, -3,
    -- filter=108 channel=32
    9, 11, 14, 8, 15, 14, 11, 16, 14,
    -- filter=108 channel=33
    9, -2, -4, -10, 0, 0, 5, 2, -7,
    -- filter=108 channel=34
    3, -5, 11, -6, -5, -7, 11, -7, -4,
    -- filter=108 channel=35
    15, 0, 2, 0, 16, 10, 5, -1, 17,
    -- filter=108 channel=36
    0, -3, 4, 3, 0, -2, 10, 9, -5,
    -- filter=108 channel=37
    0, 4, 4, 6, 0, 5, 6, -7, -7,
    -- filter=108 channel=38
    11, 2, -5, 8, -2, -3, 9, 1, -7,
    -- filter=108 channel=39
    8, 4, -3, 5, -7, -10, 3, 0, 9,
    -- filter=108 channel=40
    10, 8, -8, 2, 8, -4, 6, -4, 0,
    -- filter=108 channel=41
    9, -3, -10, 14, -4, -19, 11, -1, 4,
    -- filter=108 channel=42
    4, 7, -1, 3, 8, 0, 5, -10, 8,
    -- filter=108 channel=43
    2, 11, 13, -1, 10, 16, 10, 5, 7,
    -- filter=108 channel=44
    13, 4, 6, 2, 12, 5, 9, 15, -2,
    -- filter=108 channel=45
    -7, 2, -10, 7, 8, 10, 0, -8, 6,
    -- filter=108 channel=46
    5, 11, 4, -3, -8, -5, 2, 9, 6,
    -- filter=108 channel=47
    7, -7, 0, 0, -6, 4, -8, 7, 7,
    -- filter=108 channel=48
    1, 4, 8, -5, -2, -9, 1, -10, 2,
    -- filter=108 channel=49
    11, 3, -4, 7, -3, -10, 5, 14, 10,
    -- filter=108 channel=50
    0, 0, 0, 4, 22, 6, 4, -1, -2,
    -- filter=108 channel=51
    10, 1, 0, 6, -1, 4, -7, -3, 7,
    -- filter=108 channel=52
    -9, 10, -3, -6, 1, -7, 1, -2, 7,
    -- filter=108 channel=53
    11, 8, -1, 5, 9, 0, 7, 26, 9,
    -- filter=108 channel=54
    14, 14, 7, 6, 12, 6, 15, 7, 12,
    -- filter=108 channel=55
    -10, 0, 6, 6, -6, 2, -3, 0, -5,
    -- filter=108 channel=56
    11, -3, 5, -3, -7, 10, 0, -8, 0,
    -- filter=108 channel=57
    -6, -1, -8, -2, -10, -6, 9, 3, 4,
    -- filter=108 channel=58
    -8, 5, -6, 0, -9, 10, -6, -2, 10,
    -- filter=108 channel=59
    8, -8, 3, 14, 4, 3, 1, -1, 12,
    -- filter=108 channel=60
    9, -14, -7, 18, -2, -19, 14, -4, -5,
    -- filter=108 channel=61
    12, 0, -8, 16, 2, -15, 5, -8, -1,
    -- filter=108 channel=62
    4, -7, -13, 13, -3, -1, 3, -4, 6,
    -- filter=108 channel=63
    -6, 3, -8, -4, -10, 8, 8, -10, -9,
    -- filter=109 channel=0
    -7, -6, 0, 3, 2, -7, -9, -3, 12,
    -- filter=109 channel=1
    -16, -2, -9, -27, 4, 17, -11, 16, 15,
    -- filter=109 channel=2
    -12, -1, 2, -20, 3, 9, -21, 10, 15,
    -- filter=109 channel=3
    15, 11, 20, 16, 24, 29, 14, 12, 24,
    -- filter=109 channel=4
    -13, 1, 2, -5, 12, 10, -6, 7, 2,
    -- filter=109 channel=5
    13, 4, 13, 1, 15, 0, 9, 11, 2,
    -- filter=109 channel=6
    -16, -12, -11, 3, 11, 12, -1, -12, -8,
    -- filter=109 channel=7
    14, -5, 6, -5, 4, 3, 2, 3, -5,
    -- filter=109 channel=8
    -4, 1, 0, 6, 6, 18, 0, 17, 6,
    -- filter=109 channel=9
    6, -6, -11, 3, 6, -16, -1, 1, -6,
    -- filter=109 channel=10
    -14, -10, 3, -4, -12, -1, -16, 0, 2,
    -- filter=109 channel=11
    -19, -18, 0, -9, 10, -3, 4, 8, 11,
    -- filter=109 channel=12
    4, -6, 1, -3, -3, 8, -6, -7, 8,
    -- filter=109 channel=13
    -15, -8, -6, -3, 11, -6, 2, 5, -7,
    -- filter=109 channel=14
    2, -2, 13, 4, 5, -2, 13, 9, 10,
    -- filter=109 channel=15
    -9, -12, 0, 5, 11, -6, -8, 12, -4,
    -- filter=109 channel=16
    -2, -1, 0, 3, 6, 14, 9, 10, 16,
    -- filter=109 channel=17
    6, -3, -2, 6, 18, 2, 8, 1, 10,
    -- filter=109 channel=18
    0, -7, -8, 7, 1, -22, -1, 3, -13,
    -- filter=109 channel=19
    -5, -2, 1, -8, -2, 0, 5, 5, -4,
    -- filter=109 channel=20
    0, 8, -10, 4, 10, 3, -3, -5, 3,
    -- filter=109 channel=21
    3, 11, 0, 12, -5, 4, -7, 6, -7,
    -- filter=109 channel=22
    7, -5, 5, 6, -7, -2, 5, -2, 4,
    -- filter=109 channel=23
    -4, -9, 12, -13, -10, -3, -8, -2, 8,
    -- filter=109 channel=24
    0, -14, -10, -9, 9, 0, 3, -2, 2,
    -- filter=109 channel=25
    -22, -3, 18, -17, 16, 10, -1, 16, 23,
    -- filter=109 channel=26
    -5, -1, 0, -4, -4, -1, -3, 11, 10,
    -- filter=109 channel=27
    -5, -5, 17, -19, 9, 22, 0, 16, 16,
    -- filter=109 channel=28
    -4, 3, -14, -8, 13, 0, -4, -4, -5,
    -- filter=109 channel=29
    -15, -10, -10, 20, 13, 6, 9, 21, -3,
    -- filter=109 channel=30
    2, -1, 10, 7, 8, 5, -6, 17, 12,
    -- filter=109 channel=31
    11, -2, 7, 8, -8, -4, 9, -7, -1,
    -- filter=109 channel=32
    -8, -4, 17, -20, -3, 1, -13, 7, 17,
    -- filter=109 channel=33
    -6, 1, -5, 1, -4, -8, -8, 3, -9,
    -- filter=109 channel=34
    9, 5, -9, 9, -4, -6, 1, -4, 2,
    -- filter=109 channel=35
    -24, 4, 18, -14, 6, 22, -30, -7, 21,
    -- filter=109 channel=36
    3, 10, 3, 6, -4, 8, 0, 10, -1,
    -- filter=109 channel=37
    0, 14, 0, 19, 22, 10, 4, 22, 11,
    -- filter=109 channel=38
    -23, -4, 0, -4, 3, 3, 0, 21, 20,
    -- filter=109 channel=39
    10, 0, 0, 2, 11, -4, 5, -9, -7,
    -- filter=109 channel=40
    -3, 6, 9, 5, -9, -1, 6, 2, 0,
    -- filter=109 channel=41
    -1, -1, 12, 3, 14, 7, 14, 13, 21,
    -- filter=109 channel=42
    7, 0, 9, -4, 9, 0, 7, 8, 6,
    -- filter=109 channel=43
    -30, -44, -30, -21, -36, -35, -8, -12, -22,
    -- filter=109 channel=44
    5, 3, 20, 0, 11, 8, -5, 15, 3,
    -- filter=109 channel=45
    -3, -5, 7, 0, 8, 0, 7, -4, 6,
    -- filter=109 channel=46
    3, 5, 5, 8, 14, 9, 8, -1, -6,
    -- filter=109 channel=47
    9, 6, 0, -7, -9, 0, -7, -3, 8,
    -- filter=109 channel=48
    1, -4, -15, 4, 6, 4, 5, 4, -8,
    -- filter=109 channel=49
    -11, 5, 12, -6, 2, 9, -16, 4, -2,
    -- filter=109 channel=50
    2, -10, 4, -7, 0, 0, 3, -7, 0,
    -- filter=109 channel=51
    -7, 1, -1, -19, -9, 6, -15, -8, 4,
    -- filter=109 channel=52
    -1, -8, -1, 0, 7, 8, -8, 0, 2,
    -- filter=109 channel=53
    2, -5, 4, -8, 8, 10, -3, -3, 14,
    -- filter=109 channel=54
    11, -1, 7, 16, 15, -3, 16, 7, 6,
    -- filter=109 channel=55
    -9, -1, 0, -2, 8, 9, -10, -2, -7,
    -- filter=109 channel=56
    0, -4, -8, -6, 7, 2, 4, 1, -2,
    -- filter=109 channel=57
    1, 10, -10, -9, -9, 3, -4, 1, 3,
    -- filter=109 channel=58
    0, 4, 2, -1, -13, 3, -10, -8, -11,
    -- filter=109 channel=59
    5, 0, 9, 3, 22, 19, 4, 30, 19,
    -- filter=109 channel=60
    -15, -8, -14, -4, 25, 1, 23, 22, 20,
    -- filter=109 channel=61
    -2, -7, -6, 0, 8, 19, -11, 9, 12,
    -- filter=109 channel=62
    8, 20, 12, 0, 26, 19, 18, 17, 24,
    -- filter=109 channel=63
    -8, 2, -2, 1, 5, 2, 5, -8, -3,
    -- filter=110 channel=0
    12, 15, 4, -2, 0, 10, 13, 18, 10,
    -- filter=110 channel=1
    -11, 0, -2, -18, -19, -7, -15, -6, -2,
    -- filter=110 channel=2
    4, -13, -12, -19, -24, -15, -19, -22, -26,
    -- filter=110 channel=3
    -3, 8, 4, 5, -1, 5, 0, 2, -5,
    -- filter=110 channel=4
    -1, 19, -2, 0, 7, 6, 4, 10, 8,
    -- filter=110 channel=5
    8, 0, 8, -7, -4, -2, 1, -8, 6,
    -- filter=110 channel=6
    3, 5, -5, 5, 0, -9, 6, -9, 3,
    -- filter=110 channel=7
    2, 4, -5, 6, 4, 0, 2, 11, -3,
    -- filter=110 channel=8
    8, 15, 3, 10, 8, 0, 6, 1, -5,
    -- filter=110 channel=9
    -3, -4, 11, 0, 4, 11, -13, -2, 9,
    -- filter=110 channel=10
    -1, 5, -7, 7, -5, -4, 6, -2, 0,
    -- filter=110 channel=11
    -4, 8, 8, 2, 4, 5, -4, -2, -7,
    -- filter=110 channel=12
    0, 4, -10, 1, 2, -9, -4, 1, 8,
    -- filter=110 channel=13
    1, 13, 6, 4, 8, 14, -2, -4, -5,
    -- filter=110 channel=14
    9, 11, 0, 8, 2, 1, 5, -6, 13,
    -- filter=110 channel=15
    9, 18, 20, 2, 20, 2, -8, 10, 7,
    -- filter=110 channel=16
    -3, 7, 3, 5, -2, -1, -16, -16, -5,
    -- filter=110 channel=17
    0, 17, 10, -8, 13, 6, -9, 7, 8,
    -- filter=110 channel=18
    10, 1, 18, 14, 4, 18, 15, 6, 15,
    -- filter=110 channel=19
    -15, -13, -9, -13, -4, 1, -6, -15, -9,
    -- filter=110 channel=20
    1, -7, 5, -7, -3, 6, -7, 1, -1,
    -- filter=110 channel=21
    -5, -9, -2, 1, -2, 0, 10, 7, -3,
    -- filter=110 channel=22
    -1, 8, 1, 9, 5, -2, -5, 4, 5,
    -- filter=110 channel=23
    -9, -8, 0, 11, 8, -2, -7, 4, -11,
    -- filter=110 channel=24
    11, 9, 10, 6, 6, 1, -1, 11, 15,
    -- filter=110 channel=25
    0, -20, -23, -5, -30, -29, -5, -21, -14,
    -- filter=110 channel=26
    -2, 1, 11, -8, 8, -5, 8, -4, 4,
    -- filter=110 channel=27
    0, -5, 2, -7, -16, -18, -11, -18, -5,
    -- filter=110 channel=28
    -1, 11, 11, -7, 2, 8, -5, -10, 5,
    -- filter=110 channel=29
    0, 10, 7, -6, 10, 1, -19, -6, -13,
    -- filter=110 channel=30
    -3, 10, -5, 11, 1, -7, 8, 7, 1,
    -- filter=110 channel=31
    8, 6, -6, -3, 10, 10, -4, 0, 7,
    -- filter=110 channel=32
    -4, -15, -16, 2, -2, -11, 0, -17, -17,
    -- filter=110 channel=33
    -1, 7, 3, 7, 9, -8, -6, -5, -7,
    -- filter=110 channel=34
    5, -6, 1, -7, 7, -5, 0, 12, -4,
    -- filter=110 channel=35
    0, -10, -15, 6, 1, -18, 6, -5, -16,
    -- filter=110 channel=36
    -9, 1, -5, -5, -10, 1, 10, 0, 7,
    -- filter=110 channel=37
    0, 4, -1, 0, 9, -2, -8, 5, 1,
    -- filter=110 channel=38
    8, -8, -10, -6, -6, 1, -14, -3, -13,
    -- filter=110 channel=39
    9, 9, -7, 7, 4, 7, 4, 6, -7,
    -- filter=110 channel=40
    -3, 7, 6, 7, 4, 3, 6, -4, -3,
    -- filter=110 channel=41
    16, 1, 6, 5, -1, 1, -5, 4, 2,
    -- filter=110 channel=42
    10, 6, -7, 2, 4, -1, -3, -5, 2,
    -- filter=110 channel=43
    6, -6, 5, 8, 0, 1, -2, -9, -8,
    -- filter=110 channel=44
    -3, -15, -5, -4, -14, -5, -12, -11, -13,
    -- filter=110 channel=45
    9, 4, -9, 10, 3, 10, 9, -2, 4,
    -- filter=110 channel=46
    0, -4, 0, 5, 1, -5, 7, 4, 12,
    -- filter=110 channel=47
    -4, 5, 4, 3, -5, 5, 0, 10, 6,
    -- filter=110 channel=48
    -8, 10, 6, -5, -3, -4, -4, -10, 6,
    -- filter=110 channel=49
    -4, 6, -6, -4, 4, 11, 8, 3, 4,
    -- filter=110 channel=50
    3, -2, 8, -4, -9, 1, -5, 5, 8,
    -- filter=110 channel=51
    18, 18, -4, 18, 1, -2, 4, 15, 6,
    -- filter=110 channel=52
    6, 10, -2, 7, 5, -9, 2, 0, 5,
    -- filter=110 channel=53
    11, 0, 1, -6, -1, -8, -4, -3, 9,
    -- filter=110 channel=54
    -8, 14, 7, 6, -4, 1, -5, -6, 3,
    -- filter=110 channel=55
    2, -2, -6, -4, -2, 2, 5, -7, -1,
    -- filter=110 channel=56
    -6, 2, 7, 4, -5, 7, 0, 4, 2,
    -- filter=110 channel=57
    -2, 3, -2, -10, 1, 10, 5, 0, -4,
    -- filter=110 channel=58
    8, 2, 1, -5, 5, -10, -5, -7, -3,
    -- filter=110 channel=59
    0, 7, -4, 4, 2, -13, -11, -15, -15,
    -- filter=110 channel=60
    19, 28, 19, 16, 24, 17, -5, 13, 3,
    -- filter=110 channel=61
    17, 14, 6, 13, 16, 6, -3, 16, 15,
    -- filter=110 channel=62
    -6, -7, 6, 5, -10, 10, -7, -2, -1,
    -- filter=110 channel=63
    6, -10, 9, 5, 5, 1, 8, 9, 3,
    -- filter=111 channel=0
    8, 4, 2, -3, 6, -4, -8, -5, -9,
    -- filter=111 channel=1
    9, 7, -2, 2, 2, -4, -10, -7, 2,
    -- filter=111 channel=2
    -8, -10, -1, -6, 6, -1, 1, -5, 10,
    -- filter=111 channel=3
    10, -1, -3, 9, -1, 1, 7, 6, 4,
    -- filter=111 channel=4
    10, -5, 8, 4, 3, -7, -3, -4, -2,
    -- filter=111 channel=5
    -4, -3, 4, -5, 6, 1, 12, -7, -3,
    -- filter=111 channel=6
    0, -10, 8, 2, -10, 0, -3, -6, 6,
    -- filter=111 channel=7
    0, -6, 7, 0, 0, 7, 8, 5, 0,
    -- filter=111 channel=8
    7, -3, -11, 14, -6, -7, 10, 9, -3,
    -- filter=111 channel=9
    13, -11, -7, 18, -2, 1, 7, 0, -4,
    -- filter=111 channel=10
    -2, 5, 12, 5, -7, 10, -5, 2, 6,
    -- filter=111 channel=11
    -7, 0, 7, -4, -6, -4, 5, 0, 2,
    -- filter=111 channel=12
    5, -2, -2, 7, -8, -5, 0, 7, -4,
    -- filter=111 channel=13
    0, -10, -3, 1, 8, -12, -4, 6, 6,
    -- filter=111 channel=14
    11, 11, 6, 2, 8, 11, 4, 6, -9,
    -- filter=111 channel=15
    12, 4, 4, -7, -11, -14, 14, 8, -7,
    -- filter=111 channel=16
    -1, -4, -12, -5, 6, -12, 0, 8, 1,
    -- filter=111 channel=17
    -5, 4, -6, 5, -7, -8, 7, 9, -3,
    -- filter=111 channel=18
    10, 7, 0, 7, 7, -2, 1, 4, 7,
    -- filter=111 channel=19
    9, 11, 6, 1, -6, -7, 12, 9, 4,
    -- filter=111 channel=20
    2, 3, 5, -5, 1, -9, 3, -8, -6,
    -- filter=111 channel=21
    -2, 0, 10, 4, 0, 1, -4, 1, 3,
    -- filter=111 channel=22
    -2, 0, 9, 7, 4, 5, -4, 1, 6,
    -- filter=111 channel=23
    -2, 4, 16, -3, 0, 11, -8, 2, 1,
    -- filter=111 channel=24
    12, 0, -4, 3, 1, -8, 13, 8, -1,
    -- filter=111 channel=25
    -5, 5, 5, 0, -2, 11, -8, 4, -2,
    -- filter=111 channel=26
    -4, 0, 0, 10, 6, 8, 0, 5, 0,
    -- filter=111 channel=27
    -3, 12, -6, -7, -9, -2, -8, -6, 13,
    -- filter=111 channel=28
    -5, -11, -4, -1, -1, -14, 12, -3, -7,
    -- filter=111 channel=29
    0, 1, -3, 13, -7, -11, 5, -6, -7,
    -- filter=111 channel=30
    8, 3, 7, 21, 2, 13, 3, 14, -4,
    -- filter=111 channel=31
    0, 2, 0, 6, -1, -4, -5, -8, 0,
    -- filter=111 channel=32
    4, 1, 11, -6, 0, 1, 0, 0, 4,
    -- filter=111 channel=33
    0, -3, 1, 6, -1, 0, 8, 2, 9,
    -- filter=111 channel=34
    -7, -4, 0, 6, 10, -9, 0, -7, -4,
    -- filter=111 channel=35
    -2, 10, 15, -5, -6, 3, -13, 0, 10,
    -- filter=111 channel=36
    -10, 7, 12, -10, 9, -5, -3, 1, -6,
    -- filter=111 channel=37
    3, -1, 2, 5, -3, 0, 14, -4, 6,
    -- filter=111 channel=38
    -5, 3, -8, 2, 6, -12, 9, -7, -1,
    -- filter=111 channel=39
    7, 3, 3, 6, -8, 7, -2, -10, 10,
    -- filter=111 channel=40
    -9, -2, -5, 1, -9, -1, -5, 2, 11,
    -- filter=111 channel=41
    1, -8, 1, 7, 8, 3, -7, 10, 9,
    -- filter=111 channel=42
    7, -7, 2, 4, -7, 1, 8, 1, -10,
    -- filter=111 channel=43
    -10, -3, 4, 0, -3, 3, 0, 2, -11,
    -- filter=111 channel=44
    9, 13, 1, 11, -4, 5, 2, 6, -5,
    -- filter=111 channel=45
    -3, 8, 5, -3, -2, -5, 3, 8, -5,
    -- filter=111 channel=46
    10, 2, -3, 11, -4, -7, 11, 4, 1,
    -- filter=111 channel=47
    0, -3, 9, 7, 7, -1, -9, 4, 1,
    -- filter=111 channel=48
    -2, -8, -5, -3, -6, -2, 12, 5, 9,
    -- filter=111 channel=49
    11, -5, -7, 0, 5, 0, -9, -6, 5,
    -- filter=111 channel=50
    2, 12, 11, 5, 0, 9, 1, 13, 8,
    -- filter=111 channel=51
    -7, 7, -4, -9, 9, 14, 2, 1, 11,
    -- filter=111 channel=52
    9, -7, 6, -10, 1, 4, 3, 0, -2,
    -- filter=111 channel=53
    15, 4, 3, 13, 12, 0, 1, 0, 0,
    -- filter=111 channel=54
    13, -9, -3, 2, -6, 1, 3, 7, -4,
    -- filter=111 channel=55
    4, -3, -8, -4, 0, 2, -8, 4, 2,
    -- filter=111 channel=56
    8, 0, -5, 10, 10, 2, 4, 2, 0,
    -- filter=111 channel=57
    -8, 2, 9, 3, 0, 9, 9, -9, 3,
    -- filter=111 channel=58
    -3, 5, 7, -10, 5, -1, 5, -1, -1,
    -- filter=111 channel=59
    1, -11, 8, 8, -4, -1, -7, -5, 0,
    -- filter=111 channel=60
    9, -1, -14, 3, 0, -6, 0, 2, -11,
    -- filter=111 channel=61
    11, -6, -7, 3, 4, 6, 5, -7, -7,
    -- filter=111 channel=62
    9, 8, 0, 8, -7, -8, 12, 0, 7,
    -- filter=111 channel=63
    -10, 6, -4, 10, 0, -7, 0, -5, -1,
    -- filter=112 channel=0
    6, 0, -7, -14, 11, 16, 5, -7, 4,
    -- filter=112 channel=1
    10, -8, 12, -6, 11, 11, -6, 0, 11,
    -- filter=112 channel=2
    -8, -5, 16, -3, 0, 19, 1, -7, 12,
    -- filter=112 channel=3
    -4, 19, 17, 0, 6, 13, 3, 15, -1,
    -- filter=112 channel=4
    -10, 1, 2, -12, -7, 8, -16, -1, -6,
    -- filter=112 channel=5
    3, -3, 9, 2, -5, -9, -8, 6, -1,
    -- filter=112 channel=6
    4, -5, -6, -12, 2, -4, -4, -1, 12,
    -- filter=112 channel=7
    -10, -7, -11, -6, -2, -1, 10, -4, -10,
    -- filter=112 channel=8
    -14, 0, 0, -6, -8, 15, -18, -13, 2,
    -- filter=112 channel=9
    -6, -13, -2, 2, -18, -6, 4, -6, -15,
    -- filter=112 channel=10
    7, -1, -1, 2, 10, -1, 3, -3, -4,
    -- filter=112 channel=11
    3, -3, 7, -9, 3, 0, -18, -1, 13,
    -- filter=112 channel=12
    3, 2, -3, -2, 3, 10, -2, 8, 0,
    -- filter=112 channel=13
    -1, -2, -6, 4, 5, 5, 0, -6, 11,
    -- filter=112 channel=14
    0, -2, -2, -1, -6, 2, -9, 6, -2,
    -- filter=112 channel=15
    3, -4, 16, -9, 3, 11, -18, 3, 2,
    -- filter=112 channel=16
    0, 10, 6, -13, 0, 5, -13, 5, 9,
    -- filter=112 channel=17
    0, 8, 5, -11, -4, 0, -6, -3, 13,
    -- filter=112 channel=18
    -6, -9, 0, 9, 0, 3, 8, 1, -3,
    -- filter=112 channel=19
    -8, 1, -2, 9, 0, 0, -8, -8, 5,
    -- filter=112 channel=20
    6, -3, -4, 10, 0, 6, 9, 4, -11,
    -- filter=112 channel=21
    -5, -7, 9, -5, -5, 0, -7, -5, -6,
    -- filter=112 channel=22
    8, 9, 0, -4, -2, 6, 5, 10, -9,
    -- filter=112 channel=23
    0, -1, 3, 4, 0, -4, -5, 4, 7,
    -- filter=112 channel=24
    -4, -8, -7, 0, 5, 5, -4, -14, 12,
    -- filter=112 channel=25
    0, 10, 19, -14, 11, 19, -3, -2, 24,
    -- filter=112 channel=26
    0, -6, -9, -2, 7, -7, 0, 0, 0,
    -- filter=112 channel=27
    -13, -5, 19, -13, -1, 25, -16, -2, 17,
    -- filter=112 channel=28
    -7, 7, -7, -2, -14, 8, -3, -4, 5,
    -- filter=112 channel=29
    -9, 4, 3, -5, 5, 10, -13, 6, 8,
    -- filter=112 channel=30
    6, -2, 0, -9, -18, -14, -3, -16, 0,
    -- filter=112 channel=31
    6, 4, -8, -4, -7, 4, 0, -6, 7,
    -- filter=112 channel=32
    -2, -4, 9, 2, 0, -5, 4, -5, -1,
    -- filter=112 channel=33
    -1, -1, -4, 0, -1, 9, -6, 5, 4,
    -- filter=112 channel=34
    -8, -4, -3, 3, 3, 6, -6, 0, 4,
    -- filter=112 channel=35
    0, 4, 21, 3, 11, 14, 0, 11, 12,
    -- filter=112 channel=36
    6, 0, -5, 3, 2, -6, 4, 1, -5,
    -- filter=112 channel=37
    7, -3, 0, 10, 7, -4, 4, 10, 7,
    -- filter=112 channel=38
    0, -6, 4, 1, 11, 10, -18, 7, 23,
    -- filter=112 channel=39
    -9, -9, 6, -3, -4, 7, -6, -9, 0,
    -- filter=112 channel=40
    -9, 1, 9, 7, 5, 1, 5, 4, 8,
    -- filter=112 channel=41
    1, 5, 16, -13, 8, 12, -20, 10, 17,
    -- filter=112 channel=42
    0, -2, -2, -2, 0, -8, -6, 0, -4,
    -- filter=112 channel=43
    -4, 1, -2, 13, 12, 1, -4, -4, 1,
    -- filter=112 channel=44
    -2, -8, 0, -9, -9, -3, -1, 0, 6,
    -- filter=112 channel=45
    -3, -1, 7, -8, 3, -3, -7, 5, -2,
    -- filter=112 channel=46
    10, 4, -6, -6, -4, 7, 10, 9, -8,
    -- filter=112 channel=47
    5, 3, 3, 5, -8, 7, -3, 8, -8,
    -- filter=112 channel=48
    6, 6, 9, 7, 8, 10, 0, 0, 2,
    -- filter=112 channel=49
    3, -4, 7, -14, -10, 2, -6, -9, -2,
    -- filter=112 channel=50
    -7, 0, 0, -4, -5, -3, 0, 5, -1,
    -- filter=112 channel=51
    -3, -8, 7, -4, -3, -3, -1, -8, 7,
    -- filter=112 channel=52
    -3, -2, -7, -7, -2, -7, 1, 0, 0,
    -- filter=112 channel=53
    -9, -9, 3, 4, 4, 8, -7, -12, -4,
    -- filter=112 channel=54
    -10, 0, 0, 2, -13, -8, -8, -10, -17,
    -- filter=112 channel=55
    6, 0, 8, 0, -3, -9, -6, -1, 4,
    -- filter=112 channel=56
    6, -3, 6, 7, 8, 4, 0, -2, -7,
    -- filter=112 channel=57
    8, 2, -6, 2, 9, -9, 6, -7, 6,
    -- filter=112 channel=58
    -4, 0, 0, -6, 10, 0, 13, 0, 0,
    -- filter=112 channel=59
    6, 7, 18, -8, 17, 22, 3, 8, 25,
    -- filter=112 channel=60
    3, 5, 11, -20, -8, 24, -17, 1, 21,
    -- filter=112 channel=61
    -13, -6, 4, -11, 7, 17, -4, 1, 18,
    -- filter=112 channel=62
    12, 1, 3, 7, 4, 8, -10, 11, 15,
    -- filter=112 channel=63
    1, -7, 8, 1, 3, 2, 2, 6, 7,
    -- filter=113 channel=0
    11, 14, 2, -6, 1, 10, -12, 1, -1,
    -- filter=113 channel=1
    -5, 0, 13, -3, 0, 0, -12, 0, -5,
    -- filter=113 channel=2
    -2, 4, 16, -16, -14, -1, -1, -9, -14,
    -- filter=113 channel=3
    -2, 9, 13, -3, 7, 8, 5, 5, 0,
    -- filter=113 channel=4
    8, 15, 7, 0, 9, -2, -15, -1, -7,
    -- filter=113 channel=5
    1, 2, 5, -3, 0, 9, 0, 3, 7,
    -- filter=113 channel=6
    7, 2, 7, -12, 6, -6, -6, 2, -13,
    -- filter=113 channel=7
    7, 10, 3, 4, 3, -3, 11, -7, -5,
    -- filter=113 channel=8
    4, 22, 6, -5, 8, -2, -9, -15, -19,
    -- filter=113 channel=9
    -10, -9, -11, 0, -6, -2, -5, -6, -18,
    -- filter=113 channel=10
    1, -11, 4, 1, 10, -1, 8, 4, 4,
    -- filter=113 channel=11
    2, 17, 6, -11, 1, 2, -2, 1, -1,
    -- filter=113 channel=12
    1, 9, -6, -4, 2, -9, -3, 5, -8,
    -- filter=113 channel=13
    19, 1, 13, 9, 13, 2, -8, -4, -13,
    -- filter=113 channel=14
    4, -1, 4, -7, 8, 3, 3, 0, 11,
    -- filter=113 channel=15
    20, 11, 15, -4, 1, 0, -22, -9, -9,
    -- filter=113 channel=16
    15, 17, 14, -4, 14, 6, -10, -22, -4,
    -- filter=113 channel=17
    5, 21, 16, -11, -7, -4, -15, -15, -10,
    -- filter=113 channel=18
    -7, 0, 1, -5, -5, 6, 0, -1, -9,
    -- filter=113 channel=19
    0, -5, 0, -2, -3, 6, -2, -10, 6,
    -- filter=113 channel=20
    0, 7, 7, 3, 8, -6, -10, -3, 1,
    -- filter=113 channel=21
    -9, -9, 3, 10, -1, -9, 11, 8, -9,
    -- filter=113 channel=22
    -2, -6, 5, 1, 0, 4, -4, -1, -8,
    -- filter=113 channel=23
    -9, 10, 10, -2, -5, 6, -10, 2, 10,
    -- filter=113 channel=24
    13, 12, 10, 2, 9, 2, -8, -10, -7,
    -- filter=113 channel=25
    -3, 14, 4, 2, -6, 2, -5, -7, -14,
    -- filter=113 channel=26
    0, -4, 5, 10, -5, -2, 9, 10, 12,
    -- filter=113 channel=27
    7, 5, 15, -18, -2, 1, -18, -8, -14,
    -- filter=113 channel=28
    15, 19, 14, 5, 7, -1, 3, -9, -7,
    -- filter=113 channel=29
    29, 29, 21, -7, 15, 14, -10, -21, -10,
    -- filter=113 channel=30
    -4, 2, 8, 0, 3, 7, 9, 4, 4,
    -- filter=113 channel=31
    -7, -8, 4, 6, -8, 2, -8, -9, 1,
    -- filter=113 channel=32
    -7, 2, -12, -7, -5, -2, -6, 0, 5,
    -- filter=113 channel=33
    3, -9, 8, 4, 3, -7, 0, 7, 8,
    -- filter=113 channel=34
    -1, -3, 0, -7, -7, 10, 0, -6, -9,
    -- filter=113 channel=35
    4, 13, 2, -12, 2, 4, -11, -8, 3,
    -- filter=113 channel=36
    -3, -4, -11, 7, 2, 2, -4, -3, 1,
    -- filter=113 channel=37
    12, 8, 10, -4, 0, 10, -6, -11, 4,
    -- filter=113 channel=38
    2, 24, 6, 4, 8, 15, -17, -7, -2,
    -- filter=113 channel=39
    1, 6, -4, -4, 8, -1, 2, -7, -4,
    -- filter=113 channel=40
    8, -4, 10, -4, -4, -9, 5, -6, 3,
    -- filter=113 channel=41
    4, 28, 8, 0, 0, 5, -5, -7, -13,
    -- filter=113 channel=42
    4, 0, 10, 0, 7, 10, 1, 5, 6,
    -- filter=113 channel=43
    -6, -11, -5, 7, 8, 14, 2, -5, 5,
    -- filter=113 channel=44
    -2, -2, -3, -3, 3, -4, -1, 2, -11,
    -- filter=113 channel=45
    -3, 9, 10, 0, 8, -7, 3, -6, 4,
    -- filter=113 channel=46
    0, -3, 0, 0, 5, -7, 9, 11, 0,
    -- filter=113 channel=47
    -3, -4, 9, 0, 5, -9, -1, 5, 3,
    -- filter=113 channel=48
    12, 15, -1, -3, 6, -5, 0, -3, 6,
    -- filter=113 channel=49
    4, 15, 13, -13, -15, -1, -11, 3, 3,
    -- filter=113 channel=50
    -2, 1, -6, -2, 3, 7, 0, 0, 3,
    -- filter=113 channel=51
    3, 10, -13, 6, 7, -6, 0, 10, 9,
    -- filter=113 channel=52
    -3, -3, 10, 7, -9, 0, 2, 0, 2,
    -- filter=113 channel=53
    4, 6, 0, -5, 7, -6, 0, -9, -10,
    -- filter=113 channel=54
    5, -6, 4, -4, -17, -16, 1, -18, -1,
    -- filter=113 channel=55
    7, 10, 5, -8, 4, -7, 0, -1, 0,
    -- filter=113 channel=56
    4, 1, -2, 1, 11, 8, 7, -6, -7,
    -- filter=113 channel=57
    0, -5, -5, 8, 4, -8, 5, -4, 7,
    -- filter=113 channel=58
    0, 7, 7, -1, 7, 8, 5, 0, 2,
    -- filter=113 channel=59
    4, 8, 22, 1, -2, 5, -7, -4, -9,
    -- filter=113 channel=60
    24, 26, 21, -8, 8, 10, -6, 0, -14,
    -- filter=113 channel=61
    15, 12, 18, 6, 0, 3, -7, -18, -17,
    -- filter=113 channel=62
    14, 6, 14, 0, 9, 2, -13, -7, 0,
    -- filter=113 channel=63
    7, 6, 3, 8, 0, -4, -9, 3, 3,
    -- filter=114 channel=0
    -14, -23, -18, -7, -12, -20, -13, -10, -5,
    -- filter=114 channel=1
    2, 23, 19, 8, 36, 35, 29, 44, 41,
    -- filter=114 channel=2
    7, 44, 29, 29, 52, 38, 14, 43, 29,
    -- filter=114 channel=3
    29, 32, 23, 32, 42, 26, 30, 22, 13,
    -- filter=114 channel=4
    -27, -11, -18, -3, -18, -22, -8, -11, -17,
    -- filter=114 channel=5
    0, 3, 7, 9, 17, 14, 16, 1, 14,
    -- filter=114 channel=6
    0, 6, -5, -1, 8, 5, -8, 7, -2,
    -- filter=114 channel=7
    3, 8, -5, 6, -9, -8, 7, 3, -9,
    -- filter=114 channel=8
    -33, -25, -15, -5, -5, -21, -11, -20, -21,
    -- filter=114 channel=9
    10, 25, 30, 26, 45, 28, 14, 27, 32,
    -- filter=114 channel=10
    -2, 1, 0, 0, 3, -5, -10, 0, 5,
    -- filter=114 channel=11
    -24, -7, -10, 2, 3, 4, -6, 16, -1,
    -- filter=114 channel=12
    -3, -4, 0, -3, 5, -10, 3, -1, -2,
    -- filter=114 channel=13
    -24, -11, -17, -14, -6, -20, -2, -1, -5,
    -- filter=114 channel=14
    -6, -11, -2, -3, -11, -3, -8, -5, 1,
    -- filter=114 channel=15
    -31, -9, -16, -18, 0, -6, -21, -5, -23,
    -- filter=114 channel=16
    -13, 1, 3, 8, 21, 8, 9, 18, 10,
    -- filter=114 channel=17
    -8, -7, -25, -2, -15, -4, -8, -2, -14,
    -- filter=114 channel=18
    -21, -17, -20, -27, -31, -17, -21, -26, -19,
    -- filter=114 channel=19
    17, 31, 25, 27, 35, 28, 15, 26, 13,
    -- filter=114 channel=20
    6, 4, 0, -1, 14, 6, 3, 12, 7,
    -- filter=114 channel=21
    7, 5, 1, 2, 3, 7, -5, 6, 4,
    -- filter=114 channel=22
    9, -6, 3, -2, -10, 6, -7, -6, 9,
    -- filter=114 channel=23
    -12, -7, 7, -4, 3, 2, -5, 5, 6,
    -- filter=114 channel=24
    -25, -18, -7, -23, -6, -11, -19, -13, 0,
    -- filter=114 channel=25
    31, 61, 54, 31, 75, 50, 38, 56, 39,
    -- filter=114 channel=26
    14, 13, 0, 9, 20, 3, 17, 11, 4,
    -- filter=114 channel=27
    -2, 8, 21, 9, 17, 21, 5, 29, 13,
    -- filter=114 channel=28
    -8, -14, 0, 0, -4, 3, -3, 9, 2,
    -- filter=114 channel=29
    -18, 0, -7, 16, 8, -1, 14, 19, -9,
    -- filter=114 channel=30
    20, 13, 2, 20, 24, 21, 21, 7, 19,
    -- filter=114 channel=31
    8, -1, 8, 11, 6, 1, 8, -5, 3,
    -- filter=114 channel=32
    17, 34, 27, 17, 32, 22, 5, 22, 39,
    -- filter=114 channel=33
    -5, -9, 3, 5, 1, 3, -8, -3, 7,
    -- filter=114 channel=34
    -10, 7, 9, -3, 3, 1, -5, 14, -2,
    -- filter=114 channel=35
    -3, 35, 18, 0, 34, 20, -4, 32, 14,
    -- filter=114 channel=36
    9, 15, 0, 8, 7, 10, 8, 6, 8,
    -- filter=114 channel=37
    14, 6, 5, 16, 18, 23, 16, 30, 8,
    -- filter=114 channel=38
    -12, -7, 9, 2, 18, 14, 1, 28, 19,
    -- filter=114 channel=39
    2, 3, -8, 11, 3, 7, -6, 6, 3,
    -- filter=114 channel=40
    -7, 16, 10, -2, 9, 18, -7, -1, -1,
    -- filter=114 channel=41
    -17, -7, 1, 5, 17, -2, 6, 14, 3,
    -- filter=114 channel=42
    0, -4, -6, 1, 0, -4, 4, -10, 0,
    -- filter=114 channel=43
    -17, -9, 0, 2, -2, 4, 12, 25, 16,
    -- filter=114 channel=44
    28, 19, 21, 23, 25, 33, 13, 33, 21,
    -- filter=114 channel=45
    1, -8, -8, 0, 4, -3, -9, 7, 0,
    -- filter=114 channel=46
    2, 11, -1, -5, 10, 9, 14, 16, -5,
    -- filter=114 channel=47
    -2, -2, -6, 2, -3, 1, -1, 3, -3,
    -- filter=114 channel=48
    5, -6, -9, 10, 21, -2, 3, 0, -8,
    -- filter=114 channel=49
    -4, 3, 2, -16, -9, -1, -14, -3, -18,
    -- filter=114 channel=50
    4, -4, -4, -2, -4, -1, 11, 16, 13,
    -- filter=114 channel=51
    -18, -16, -26, -16, -36, -26, -28, -20, -21,
    -- filter=114 channel=52
    -8, 8, -2, 4, 9, -2, -1, -2, 2,
    -- filter=114 channel=53
    1, 27, 20, 12, 24, 32, 4, 28, 34,
    -- filter=114 channel=54
    15, 27, 28, 33, 44, 24, 17, 23, 23,
    -- filter=114 channel=55
    -2, 7, 0, -2, 8, -4, -2, 0, -4,
    -- filter=114 channel=56
    3, -3, -1, -5, -7, -9, 3, -7, -8,
    -- filter=114 channel=57
    -8, 0, 6, -4, -9, 4, 8, 5, -4,
    -- filter=114 channel=58
    0, 17, 2, 2, 6, 8, 18, 1, 5,
    -- filter=114 channel=59
    18, 21, 12, 18, 32, 27, 24, 16, 22,
    -- filter=114 channel=60
    -33, -38, -38, -10, -5, -10, -19, -11, -29,
    -- filter=114 channel=61
    -23, -30, -26, -27, -21, -14, -23, -20, -9,
    -- filter=114 channel=62
    11, 15, 19, 8, 34, 19, 11, 22, 11,
    -- filter=114 channel=63
    -5, -7, -5, 0, 5, 1, -4, -8, -3,
    -- filter=115 channel=0
    -1, 0, -8, 4, -3, -5, 6, -6, 0,
    -- filter=115 channel=1
    3, 0, 0, -6, -1, 3, -9, 4, 3,
    -- filter=115 channel=2
    7, -6, -9, -4, 9, 6, -7, 6, -1,
    -- filter=115 channel=3
    -1, -8, 6, 2, -6, 0, 5, -10, 0,
    -- filter=115 channel=4
    -6, -1, 5, -6, 8, -9, 4, -9, -1,
    -- filter=115 channel=5
    8, 9, -2, 3, -8, -4, -6, -7, -3,
    -- filter=115 channel=6
    10, 9, 4, -4, -9, -5, 7, -10, -6,
    -- filter=115 channel=7
    -6, -6, 3, -2, -2, 0, -9, 0, -4,
    -- filter=115 channel=8
    0, 7, 1, -8, -5, -6, -3, 7, 10,
    -- filter=115 channel=9
    -4, 7, -6, -2, -5, 8, -10, 8, 0,
    -- filter=115 channel=10
    3, -6, 4, 11, 2, 1, 10, 0, 9,
    -- filter=115 channel=11
    -6, 3, -3, 4, -6, 2, 6, -1, -6,
    -- filter=115 channel=12
    -1, 0, 2, 9, 7, 2, 1, -3, -10,
    -- filter=115 channel=13
    9, -7, -6, -8, -7, 7, 1, -7, 9,
    -- filter=115 channel=14
    5, -5, 6, 7, 0, -7, -2, 8, 5,
    -- filter=115 channel=15
    -7, 6, -8, -10, 10, 2, -6, 9, 7,
    -- filter=115 channel=16
    -6, -2, -8, 3, 5, 4, 7, 9, 6,
    -- filter=115 channel=17
    -7, -9, -5, -7, 2, 0, -2, -7, -7,
    -- filter=115 channel=18
    10, 7, -3, 9, 0, 7, -7, 4, 4,
    -- filter=115 channel=19
    -6, 2, 0, -8, 4, -3, -7, -6, 2,
    -- filter=115 channel=20
    6, 11, -2, 5, 5, 3, -5, 5, 6,
    -- filter=115 channel=21
    -9, 2, -5, 0, -8, 10, 2, 7, -3,
    -- filter=115 channel=22
    0, 0, -1, 2, 8, -2, 2, 1, 7,
    -- filter=115 channel=23
    -9, -7, -5, -1, 5, 5, 1, 9, -9,
    -- filter=115 channel=24
    6, 1, -8, -6, -7, -2, -7, -1, 0,
    -- filter=115 channel=25
    1, -9, 8, -9, 7, -3, 3, -3, 8,
    -- filter=115 channel=26
    8, 0, 2, 4, 7, 7, 8, 8, 0,
    -- filter=115 channel=27
    10, 0, 5, -8, -9, -5, -6, 5, 10,
    -- filter=115 channel=28
    -4, 0, -5, -5, -8, 4, -7, -10, -3,
    -- filter=115 channel=29
    -2, -1, 2, 7, 10, -5, -9, 2, 0,
    -- filter=115 channel=30
    7, 2, 11, -2, 4, -4, 0, 4, 7,
    -- filter=115 channel=31
    2, -7, -4, 8, 0, 1, -9, -10, -4,
    -- filter=115 channel=32
    -5, 0, -8, 10, -2, 0, -3, -7, 5,
    -- filter=115 channel=33
    -5, 8, -6, -1, -3, -1, 3, -4, -1,
    -- filter=115 channel=34
    -5, -8, -9, 5, 0, 1, -9, -1, -4,
    -- filter=115 channel=35
    -1, -7, -9, 1, 3, -9, 7, 5, -8,
    -- filter=115 channel=36
    1, 8, -2, 0, 10, 4, 5, -9, -1,
    -- filter=115 channel=37
    -8, 0, 9, -3, 0, -5, 3, 0, 2,
    -- filter=115 channel=38
    -5, -1, -6, -1, -4, -1, 8, 9, -7,
    -- filter=115 channel=39
    -10, 0, -4, 8, -1, -8, -5, 2, 9,
    -- filter=115 channel=40
    -1, -8, 10, 7, -7, -6, 2, 8, 6,
    -- filter=115 channel=41
    1, 11, 10, 0, 8, 8, -2, 9, -5,
    -- filter=115 channel=42
    7, -10, 5, 3, 3, -6, 7, -3, -1,
    -- filter=115 channel=43
    -2, -6, -10, -9, -2, 9, -5, 0, -4,
    -- filter=115 channel=44
    5, 0, 8, -2, -4, -7, 0, -3, -7,
    -- filter=115 channel=45
    9, -6, -2, -7, 0, -9, -1, 2, -1,
    -- filter=115 channel=46
    -7, 6, -6, 9, 2, -6, 4, 9, -6,
    -- filter=115 channel=47
    8, 8, 1, 5, -8, 0, -3, 7, -3,
    -- filter=115 channel=48
    5, -6, -5, 6, 1, -8, -6, 8, 10,
    -- filter=115 channel=49
    -8, 0, 1, 4, -5, 2, -9, 0, 1,
    -- filter=115 channel=50
    0, 4, 4, 6, 4, 1, 0, 0, 8,
    -- filter=115 channel=51
    -1, -8, 9, 0, 5, -2, 4, 8, 9,
    -- filter=115 channel=52
    3, -5, 4, 9, -1, -2, -4, 7, 9,
    -- filter=115 channel=53
    -10, 3, 0, -7, -9, -5, -6, -9, -8,
    -- filter=115 channel=54
    -2, 7, 6, -8, 8, -6, -1, 5, 8,
    -- filter=115 channel=55
    -1, -9, -9, -2, -4, 5, 6, 1, -6,
    -- filter=115 channel=56
    -10, 9, 0, 1, -5, -6, 7, -10, 5,
    -- filter=115 channel=57
    0, 2, 0, -5, -2, -2, 1, 8, -4,
    -- filter=115 channel=58
    4, -5, 1, 9, 0, -5, 11, 8, -9,
    -- filter=115 channel=59
    11, -2, 3, 3, -6, 4, -4, 9, -8,
    -- filter=115 channel=60
    1, -7, 0, -8, 4, -10, 1, 5, 4,
    -- filter=115 channel=61
    -1, 6, 7, -10, 8, 5, -4, 7, -9,
    -- filter=115 channel=62
    -8, -5, 0, 1, 5, -4, 7, 8, -4,
    -- filter=115 channel=63
    -3, -4, -8, 4, -7, 8, 0, -1, -5,
    -- filter=116 channel=0
    -7, -12, -3, 5, -4, -1, -3, 11, -7,
    -- filter=116 channel=1
    -3, -5, -16, -14, -1, 3, -7, -1, -9,
    -- filter=116 channel=2
    -15, -19, -7, 2, 6, -5, -10, -14, -11,
    -- filter=116 channel=3
    12, -4, -9, 22, 18, 14, 1, 16, 5,
    -- filter=116 channel=4
    -13, -4, -2, 11, 16, -2, 7, 13, 11,
    -- filter=116 channel=5
    15, -6, 0, 0, 2, -5, 10, -1, 10,
    -- filter=116 channel=6
    -12, -13, -15, 3, 12, 8, 7, 7, -1,
    -- filter=116 channel=7
    1, -4, -13, 0, 2, 7, 6, 4, -2,
    -- filter=116 channel=8
    -3, -17, -13, 17, 15, -2, 22, 10, -2,
    -- filter=116 channel=9
    -10, 2, -15, 12, 14, -6, 16, 22, -3,
    -- filter=116 channel=10
    -10, 0, -2, -10, -9, -6, 1, -11, 3,
    -- filter=116 channel=11
    -18, -8, -11, -7, 2, 0, 1, 2, 11,
    -- filter=116 channel=12
    -6, 10, 7, -3, 0, 5, -5, -9, -7,
    -- filter=116 channel=13
    -19, -15, -7, 11, 8, -2, 14, 22, 2,
    -- filter=116 channel=14
    5, 0, 8, -4, -7, 8, 6, 6, -3,
    -- filter=116 channel=15
    -11, -4, -15, 21, 15, -1, 14, 5, -5,
    -- filter=116 channel=16
    -12, -8, -33, 25, 2, 3, 25, 17, 0,
    -- filter=116 channel=17
    0, -4, -9, 18, 14, 15, 16, 8, 2,
    -- filter=116 channel=18
    3, -2, -9, 17, 10, 3, 13, 4, 6,
    -- filter=116 channel=19
    -2, -13, -15, -1, -1, 0, -3, 3, 7,
    -- filter=116 channel=20
    3, 4, 0, 0, 0, -11, -2, -3, -5,
    -- filter=116 channel=21
    0, -1, 1, 0, -9, 7, 5, 0, -9,
    -- filter=116 channel=22
    -3, -6, -3, 6, -7, 0, 0, 3, 7,
    -- filter=116 channel=23
    -1, -8, 4, 0, -5, -2, 3, -8, 0,
    -- filter=116 channel=24
    -2, -8, -10, 3, 16, 5, 7, 10, 14,
    -- filter=116 channel=25
    -3, -20, -18, -7, -1, 3, -2, -8, -3,
    -- filter=116 channel=26
    -9, -3, -4, -15, -5, -15, 0, 2, -13,
    -- filter=116 channel=27
    6, -13, -5, 8, 8, -4, -6, 17, 0,
    -- filter=116 channel=28
    -8, -9, -10, 19, 18, 7, -3, 3, 9,
    -- filter=116 channel=29
    -17, -15, -33, 25, 17, -6, 27, 23, -3,
    -- filter=116 channel=30
    -12, -8, -7, -1, -17, -19, 2, -4, -11,
    -- filter=116 channel=31
    7, 7, 13, 1, 0, -6, 6, -8, 3,
    -- filter=116 channel=32
    -9, 2, -8, -19, -16, 4, -16, -2, -1,
    -- filter=116 channel=33
    -2, 0, -9, -2, -6, 7, -6, 7, 0,
    -- filter=116 channel=34
    3, 0, -10, 1, -6, -6, 6, 10, 6,
    -- filter=116 channel=35
    -14, 3, 9, -12, -3, 10, -18, 0, -1,
    -- filter=116 channel=36
    13, 7, 9, 11, 0, 7, 7, -7, 0,
    -- filter=116 channel=37
    11, -7, -9, 7, 8, 6, 3, 18, 11,
    -- filter=116 channel=38
    -3, -13, -11, 0, 12, -1, 17, 18, 8,
    -- filter=116 channel=39
    8, 3, 7, -1, 0, 4, -7, 1, 8,
    -- filter=116 channel=40
    3, 10, -4, 6, -2, 6, 3, -4, 7,
    -- filter=116 channel=41
    6, -1, -21, 19, 21, 0, 11, 14, 1,
    -- filter=116 channel=42
    -6, -2, 8, 0, 6, 0, 6, 8, -1,
    -- filter=116 channel=43
    -29, -39, -17, -18, -40, -35, -7, -19, -15,
    -- filter=116 channel=44
    4, -9, -3, -11, -6, 3, -10, -4, 2,
    -- filter=116 channel=45
    -7, 1, 5, 1, 3, 1, 9, 5, -5,
    -- filter=116 channel=46
    2, 3, -12, 3, -7, -13, 6, -1, -10,
    -- filter=116 channel=47
    5, 8, 0, 7, -1, -4, -3, 10, 0,
    -- filter=116 channel=48
    -10, -14, -15, 3, 8, -2, 10, -2, -5,
    -- filter=116 channel=49
    -4, 15, 9, 6, 20, 20, -15, 2, 0,
    -- filter=116 channel=50
    -7, -14, -9, -17, -25, -25, -11, -2, -3,
    -- filter=116 channel=51
    9, 4, 5, -3, 5, -4, -11, 1, 10,
    -- filter=116 channel=52
    -5, -3, 10, -6, 9, 2, 3, 0, -4,
    -- filter=116 channel=53
    -8, -16, -10, -10, -19, -16, -4, -3, 7,
    -- filter=116 channel=54
    4, -6, -14, 4, 16, 3, 12, 19, 7,
    -- filter=116 channel=55
    5, 2, 10, -9, 4, 7, 0, 1, -4,
    -- filter=116 channel=56
    4, 6, 2, -10, -5, -7, -1, -7, -5,
    -- filter=116 channel=57
    -3, -6, 0, 0, -5, -3, -6, -5, -7,
    -- filter=116 channel=58
    0, 0, -2, 2, -11, -9, 3, -2, -5,
    -- filter=116 channel=59
    -9, -6, -9, 18, 8, -9, 8, 5, 11,
    -- filter=116 channel=60
    -8, -4, -17, 10, 19, 5, 36, 32, 18,
    -- filter=116 channel=61
    0, -1, -9, 15, 5, 10, 16, 22, 5,
    -- filter=116 channel=62
    -2, -4, -9, 13, 0, 6, 8, 16, 7,
    -- filter=116 channel=63
    -2, 10, -8, 4, 0, -1, 0, 0, -2,
    -- filter=117 channel=0
    -4, -1, 1, 7, 0, 4, 5, 0, -11,
    -- filter=117 channel=1
    -9, 0, -6, 6, 5, -6, 8, -3, 9,
    -- filter=117 channel=2
    11, -1, 0, 12, 10, 0, -8, 0, 8,
    -- filter=117 channel=3
    -15, 0, -10, 6, -2, 5, -12, -8, -5,
    -- filter=117 channel=4
    0, 7, 3, 12, 6, 7, 4, -1, -4,
    -- filter=117 channel=5
    3, -1, 7, 5, -3, -8, 2, 6, -8,
    -- filter=117 channel=6
    -6, -5, 2, 7, -6, -1, 11, -4, -8,
    -- filter=117 channel=7
    0, 5, -4, 4, -4, 10, 6, 5, -4,
    -- filter=117 channel=8
    2, -2, -12, 3, 0, -6, 4, 2, -3,
    -- filter=117 channel=9
    -7, -7, 6, -12, -10, 5, -11, 4, -9,
    -- filter=117 channel=10
    -5, 5, -10, -5, -1, 0, 10, 8, 7,
    -- filter=117 channel=11
    1, 4, -13, -6, -6, 2, 10, 11, -7,
    -- filter=117 channel=12
    -6, -5, -10, -1, 2, -8, 9, 3, -8,
    -- filter=117 channel=13
    -9, 5, -11, 12, -4, -6, 9, 9, 7,
    -- filter=117 channel=14
    -10, 6, -6, 7, -9, 0, 9, -7, -3,
    -- filter=117 channel=15
    -2, 1, 3, 18, 11, -1, -1, 8, -8,
    -- filter=117 channel=16
    -6, -9, -3, -2, 2, 11, 6, -1, 1,
    -- filter=117 channel=17
    3, -1, -8, -1, 6, 0, 1, 6, -4,
    -- filter=117 channel=18
    -1, 2, 13, 10, 11, -2, 11, 7, -2,
    -- filter=117 channel=19
    -4, 1, 10, 2, 9, 4, -8, -7, -2,
    -- filter=117 channel=20
    -2, 0, -9, 5, -11, -2, -4, -3, 7,
    -- filter=117 channel=21
    -2, -4, 3, 3, -5, 7, -10, -9, -3,
    -- filter=117 channel=22
    0, -3, -8, 0, 2, -2, -5, 9, 0,
    -- filter=117 channel=23
    3, -10, -7, -6, 1, -10, -5, -2, 11,
    -- filter=117 channel=24
    8, 8, 6, 0, 0, 4, -3, 12, 5,
    -- filter=117 channel=25
    0, -7, 0, 11, 6, 8, 3, -7, -8,
    -- filter=117 channel=26
    4, -1, -7, 2, -3, -5, 7, -10, 1,
    -- filter=117 channel=27
    -1, -9, -2, -1, 4, -3, -2, 0, -9,
    -- filter=117 channel=28
    13, 5, 8, 8, 12, 5, 4, 9, 2,
    -- filter=117 channel=29
    -7, 5, 0, 18, 13, 7, -5, 10, 8,
    -- filter=117 channel=30
    -10, -6, -9, 7, 0, 4, -5, 6, -5,
    -- filter=117 channel=31
    1, -1, 4, -10, 2, -7, -11, -8, 3,
    -- filter=117 channel=32
    0, -11, 2, -10, -12, -7, -2, -7, 6,
    -- filter=117 channel=33
    9, 7, 9, -3, -6, -4, -1, 10, 0,
    -- filter=117 channel=34
    -2, -6, 6, -3, -3, 7, 0, 10, -6,
    -- filter=117 channel=35
    -4, -12, 1, -8, -4, 9, 3, 2, 0,
    -- filter=117 channel=36
    -5, -6, 1, 8, 7, 2, -10, -7, -3,
    -- filter=117 channel=37
    1, 0, -12, -9, -4, 5, -10, -4, -3,
    -- filter=117 channel=38
    -6, -4, -1, 0, 0, -8, 11, 11, -6,
    -- filter=117 channel=39
    8, -1, -2, -6, -2, -2, 7, 4, 0,
    -- filter=117 channel=40
    5, -1, 0, 0, -2, 0, -1, -5, -6,
    -- filter=117 channel=41
    7, 1, -7, 11, 6, 1, 9, -2, -4,
    -- filter=117 channel=42
    0, -1, 10, 7, -2, -7, 9, 10, 3,
    -- filter=117 channel=43
    -4, -6, -8, 0, -13, 8, 0, 7, 4,
    -- filter=117 channel=44
    4, -4, -3, -3, 0, 4, -12, 4, 0,
    -- filter=117 channel=45
    0, 2, -7, -6, -4, -6, 7, 3, 4,
    -- filter=117 channel=46
    2, 0, 0, -9, -3, -3, -7, -1, 9,
    -- filter=117 channel=47
    -3, -4, 7, -1, 7, 9, -9, 3, 2,
    -- filter=117 channel=48
    -4, 3, -8, 9, 2, -7, 8, 9, -7,
    -- filter=117 channel=49
    0, -1, 3, -4, -4, 11, 2, -4, -8,
    -- filter=117 channel=50
    3, 0, -9, 8, 9, -4, -1, 12, 13,
    -- filter=117 channel=51
    -2, 4, 8, -5, 7, 8, 10, 0, 7,
    -- filter=117 channel=52
    0, -5, 6, 0, 3, 5, 6, -7, 6,
    -- filter=117 channel=53
    -6, 9, -3, -12, 5, 0, -11, 2, 8,
    -- filter=117 channel=54
    -9, -15, 2, 0, 4, 0, 0, -10, -7,
    -- filter=117 channel=55
    -1, -5, -6, 0, 6, 3, -2, 5, -10,
    -- filter=117 channel=56
    -2, -6, -4, -2, -2, 10, -7, -6, -1,
    -- filter=117 channel=57
    -7, 2, 7, 8, 2, 8, -4, -1, -9,
    -- filter=117 channel=58
    -7, 5, -2, -9, -1, 1, -7, 1, 11,
    -- filter=117 channel=59
    -12, -9, -17, -9, -9, -2, -8, -10, -13,
    -- filter=117 channel=60
    4, -6, -6, 16, 6, -2, 0, 6, 5,
    -- filter=117 channel=61
    0, -8, -9, 0, 4, 6, 0, 6, -4,
    -- filter=117 channel=62
    4, 2, -6, -7, 7, 5, -6, -13, 1,
    -- filter=117 channel=63
    5, 4, -10, -7, -6, 0, -6, -4, -6,
    -- filter=118 channel=0
    -6, -10, 1, -7, 0, -7, 0, -5, -6,
    -- filter=118 channel=1
    2, -9, 0, -2, 9, -1, 7, -6, -3,
    -- filter=118 channel=2
    4, 3, 3, -8, -6, 9, 7, 6, 4,
    -- filter=118 channel=3
    9, 1, -7, 1, 8, -3, -7, -2, 3,
    -- filter=118 channel=4
    -9, 0, 0, -4, 8, -7, 4, 7, -2,
    -- filter=118 channel=5
    -8, 0, 0, -2, 7, -8, 1, 8, -4,
    -- filter=118 channel=6
    -6, -4, 0, -5, 5, 7, 6, 8, 0,
    -- filter=118 channel=7
    9, -3, 4, 1, 4, 0, 8, 2, -3,
    -- filter=118 channel=8
    -3, -6, -9, 3, -7, -6, 2, 7, -6,
    -- filter=118 channel=9
    0, -5, 4, -1, -3, 0, 6, 0, 0,
    -- filter=118 channel=10
    4, -5, 10, 10, -1, 1, -8, 0, -9,
    -- filter=118 channel=11
    -4, 2, -1, -3, 5, -1, -6, -9, -5,
    -- filter=118 channel=12
    4, 0, 8, -1, -8, 8, 2, 2, -10,
    -- filter=118 channel=13
    -6, 2, -9, 6, -1, -9, 0, 1, 3,
    -- filter=118 channel=14
    7, -1, 6, 6, -5, -4, 7, 6, 1,
    -- filter=118 channel=15
    4, 2, 2, 7, -5, -1, -2, -5, 10,
    -- filter=118 channel=16
    4, 0, -9, 0, -10, 7, -7, -3, 10,
    -- filter=118 channel=17
    4, -10, -7, -9, 4, 8, 4, 4, 10,
    -- filter=118 channel=18
    -2, 6, 6, 6, 3, -2, 0, 6, 8,
    -- filter=118 channel=19
    -5, 8, 8, 5, 0, 3, 9, 6, -3,
    -- filter=118 channel=20
    8, -6, -1, -6, -1, 1, 8, 2, 3,
    -- filter=118 channel=21
    4, -1, -3, -1, -2, 8, 1, 6, 8,
    -- filter=118 channel=22
    -3, -10, 4, 5, 7, -3, 0, -7, -3,
    -- filter=118 channel=23
    -3, -5, 1, -7, -7, -4, 7, 5, -3,
    -- filter=118 channel=24
    -1, 9, -3, 6, -5, 7, 7, 8, -3,
    -- filter=118 channel=25
    -2, -5, 3, 1, 7, 6, -3, 9, -2,
    -- filter=118 channel=26
    10, -9, 5, 10, -4, -5, -7, 4, 3,
    -- filter=118 channel=27
    7, -4, -10, -3, -7, -6, 8, -5, -4,
    -- filter=118 channel=28
    8, 0, 6, 8, 5, -3, 1, 1, -5,
    -- filter=118 channel=29
    6, -8, -5, -2, -8, -2, -1, 0, 6,
    -- filter=118 channel=30
    -8, 0, -8, 3, 9, 0, 11, 0, 1,
    -- filter=118 channel=31
    -5, 7, -6, -2, 1, 11, 5, -4, 1,
    -- filter=118 channel=32
    -7, 3, -9, -6, 6, 8, 10, 0, 8,
    -- filter=118 channel=33
    -10, -5, 0, -9, 8, -2, 9, -1, 0,
    -- filter=118 channel=34
    0, 1, 7, 7, -5, 2, 8, 5, -2,
    -- filter=118 channel=35
    -5, 0, -3, -3, 9, -5, -8, 3, -8,
    -- filter=118 channel=36
    -1, -8, 6, -10, -6, 7, -7, 6, 3,
    -- filter=118 channel=37
    0, -2, 10, 6, 0, 6, 9, 2, -8,
    -- filter=118 channel=38
    4, -9, -7, -8, -9, 0, 8, -2, -6,
    -- filter=118 channel=39
    0, 7, -6, -5, 9, 7, 1, 4, 1,
    -- filter=118 channel=40
    0, 5, -2, 5, 7, 9, 4, 1, -2,
    -- filter=118 channel=41
    -10, -3, 2, 4, -7, 1, -3, -7, -4,
    -- filter=118 channel=42
    -4, -8, -2, 3, 4, -5, -10, -6, -6,
    -- filter=118 channel=43
    -6, -8, -7, -10, -5, -7, 0, 1, 4,
    -- filter=118 channel=44
    8, 1, 6, -4, -3, -9, 0, -9, 4,
    -- filter=118 channel=45
    0, -7, -1, -7, -5, 1, -9, 6, -5,
    -- filter=118 channel=46
    1, 0, -6, 1, -2, -9, -3, 10, 4,
    -- filter=118 channel=47
    -5, -6, -3, 3, -7, 0, -9, 9, 7,
    -- filter=118 channel=48
    -4, 8, 1, -4, -1, -6, 3, 9, -3,
    -- filter=118 channel=49
    5, 9, -6, -3, 0, 3, 11, -9, 3,
    -- filter=118 channel=50
    6, 3, 7, 7, 1, -4, 11, 0, -9,
    -- filter=118 channel=51
    10, 3, 9, -5, -5, -5, 0, -9, -8,
    -- filter=118 channel=52
    -9, -6, 8, 8, 5, 6, -4, -3, 3,
    -- filter=118 channel=53
    5, 9, -4, 10, -4, -1, 11, 4, 8,
    -- filter=118 channel=54
    -2, 2, -5, 11, 9, -5, 2, 7, 3,
    -- filter=118 channel=55
    4, 6, 2, -8, -4, -1, -6, 2, -4,
    -- filter=118 channel=56
    9, 6, 3, 0, 5, -9, 5, 1, 3,
    -- filter=118 channel=57
    -5, -10, 0, 5, -10, 0, 1, 7, -4,
    -- filter=118 channel=58
    3, 0, 7, -4, 10, -4, 7, -2, 4,
    -- filter=118 channel=59
    -7, 8, -10, -1, 0, -3, -2, -5, 3,
    -- filter=118 channel=60
    -8, -5, 6, -4, 6, -7, 6, 5, -5,
    -- filter=118 channel=61
    5, -10, 5, 2, 5, -1, 2, 0, -2,
    -- filter=118 channel=62
    8, 6, 0, -3, 0, 3, 7, 0, 2,
    -- filter=118 channel=63
    -6, 0, 10, 0, -3, -6, -9, -6, 2,
    -- filter=119 channel=0
    -13, 6, 14, -24, -8, 27, -10, -12, 23,
    -- filter=119 channel=1
    0, -12, 0, 12, -28, 7, 12, -22, -3,
    -- filter=119 channel=2
    -1, -25, 10, -11, -14, 22, -5, -19, 9,
    -- filter=119 channel=3
    -8, 0, 11, 0, 1, 18, -11, -1, 20,
    -- filter=119 channel=4
    -7, -5, 10, -3, -1, 12, -6, -4, 4,
    -- filter=119 channel=5
    17, 0, -5, 22, 4, -1, 17, 5, -3,
    -- filter=119 channel=6
    -16, -8, -1, -2, -4, 20, -5, -6, 17,
    -- filter=119 channel=7
    8, 18, 5, 6, 13, -1, 10, 5, 17,
    -- filter=119 channel=8
    11, -23, 17, -4, -32, 21, -2, -6, 23,
    -- filter=119 channel=9
    18, -4, 1, 10, -1, -15, 1, -6, -19,
    -- filter=119 channel=10
    0, 2, -3, -19, -6, -4, -8, -8, 8,
    -- filter=119 channel=11
    -2, -4, -8, 1, -12, 19, 1, -9, 10,
    -- filter=119 channel=12
    4, 1, -4, 4, -9, 1, -12, -9, 5,
    -- filter=119 channel=13
    -15, -3, -2, -3, -10, 17, -18, -2, 18,
    -- filter=119 channel=14
    9, 0, 3, 13, 6, 0, 10, 15, 6,
    -- filter=119 channel=15
    -13, -10, 33, -7, -23, 45, -9, -24, 23,
    -- filter=119 channel=16
    -8, -30, 13, 7, -26, 38, -3, -27, 22,
    -- filter=119 channel=17
    3, -10, 8, 11, -27, 3, 10, -20, 7,
    -- filter=119 channel=18
    -4, -3, -5, -6, 6, 16, -1, 11, 7,
    -- filter=119 channel=19
    24, -13, -8, 30, -3, -13, 16, -3, 1,
    -- filter=119 channel=20
    3, 0, 15, -7, 9, 20, -14, 14, 10,
    -- filter=119 channel=21
    -4, 4, 2, -1, 4, -3, -11, -10, 0,
    -- filter=119 channel=22
    10, 0, 0, -2, -7, -9, 0, -1, -10,
    -- filter=119 channel=23
    -7, -2, 2, -1, -11, 7, 0, -2, 17,
    -- filter=119 channel=24
    17, -7, -3, 6, -11, 2, 10, -6, 11,
    -- filter=119 channel=25
    -2, -12, 6, -25, -27, 20, -8, -23, 7,
    -- filter=119 channel=26
    4, 5, 19, 6, 18, 36, -10, 19, 15,
    -- filter=119 channel=27
    2, -25, 22, -5, -27, 19, 0, -27, 19,
    -- filter=119 channel=28
    1, -7, 1, 24, -25, 4, 4, -12, -9,
    -- filter=119 channel=29
    -1, -27, 25, -3, -33, 41, -6, -25, 34,
    -- filter=119 channel=30
    52, 32, 27, 69, 13, 23, 47, 24, 28,
    -- filter=119 channel=31
    -7, -7, 7, 2, -5, 2, -4, 0, 4,
    -- filter=119 channel=32
    9, -11, 8, 5, -2, -2, -6, 0, 9,
    -- filter=119 channel=33
    1, -2, 10, -5, -7, -7, 0, 5, 0,
    -- filter=119 channel=34
    2, -2, 16, 11, 14, 24, 12, 14, 14,
    -- filter=119 channel=35
    -12, -15, 16, -19, -15, 36, -16, -23, 15,
    -- filter=119 channel=36
    5, 9, -10, 9, -5, -4, -8, -9, 4,
    -- filter=119 channel=37
    12, -6, 9, 15, -9, 14, 7, -2, 14,
    -- filter=119 channel=38
    3, -29, 13, -8, -29, 29, 3, -20, 35,
    -- filter=119 channel=39
    -5, 4, -9, -4, -3, 5, 9, 3, 0,
    -- filter=119 channel=40
    -8, -11, 0, -10, -12, -1, -3, 0, -6,
    -- filter=119 channel=41
    -1, -34, 30, -11, -29, 34, -8, -27, 31,
    -- filter=119 channel=42
    1, 7, -8, 4, 8, -1, 0, -7, 0,
    -- filter=119 channel=43
    1, -4, -24, 0, -15, -16, -9, -10, -6,
    -- filter=119 channel=44
    0, 12, 0, 23, -8, -2, 6, -3, -4,
    -- filter=119 channel=45
    7, 0, 8, -5, 6, 5, -10, 7, 4,
    -- filter=119 channel=46
    -3, 4, 14, 3, 12, 21, -5, 11, 20,
    -- filter=119 channel=47
    0, -8, 3, 9, 5, 3, 2, -4, -5,
    -- filter=119 channel=48
    -17, -11, 12, -21, 1, 8, -2, -3, 7,
    -- filter=119 channel=49
    -8, -15, 24, -14, -1, 16, 2, -10, 11,
    -- filter=119 channel=50
    12, 21, 13, 39, 12, 14, 26, 20, 21,
    -- filter=119 channel=51
    -9, 1, 12, -11, 0, -1, 0, 3, -3,
    -- filter=119 channel=52
    -2, -4, 0, -10, 4, 9, 10, 1, 3,
    -- filter=119 channel=53
    21, 10, 19, 40, 21, 9, 31, 14, 22,
    -- filter=119 channel=54
    7, -12, -8, 20, -15, 3, 20, -6, -2,
    -- filter=119 channel=55
    -8, -10, -9, 6, 7, -1, 1, -2, 4,
    -- filter=119 channel=56
    -1, 3, 6, 2, 11, 12, 0, 3, 6,
    -- filter=119 channel=57
    -4, 0, -8, -7, 8, 0, 6, -4, 4,
    -- filter=119 channel=58
    0, 0, 4, -2, 10, -2, -17, -8, -10,
    -- filter=119 channel=59
    -4, -12, 16, -12, -25, 38, -8, -5, 30,
    -- filter=119 channel=60
    -4, -12, 21, -22, -28, 55, -19, -28, 52,
    -- filter=119 channel=61
    10, -17, 18, -1, -18, 24, 10, -16, 20,
    -- filter=119 channel=62
    16, -17, -3, 7, -18, 10, 11, 0, 9,
    -- filter=119 channel=63
    -7, 0, 9, 9, 0, 6, -7, -10, 10,
    -- filter=120 channel=0
    -15, -5, 7, -18, 7, 1, -11, -3, 4,
    -- filter=120 channel=1
    -9, -16, 0, -13, -9, 8, -7, -4, 10,
    -- filter=120 channel=2
    -18, -3, 23, -7, 9, 33, 1, -1, 5,
    -- filter=120 channel=3
    -3, 7, 24, 11, 19, 23, 6, 16, 21,
    -- filter=120 channel=4
    -14, -10, 6, -17, 5, 17, -1, 10, 14,
    -- filter=120 channel=5
    -11, 2, 1, -8, -3, 4, 1, 7, -5,
    -- filter=120 channel=6
    -2, 3, 13, -13, 9, 3, 4, -4, -2,
    -- filter=120 channel=7
    -2, 3, -2, -2, 4, -6, 4, -12, -11,
    -- filter=120 channel=8
    -35, -23, 10, -8, 11, 24, -18, -4, 17,
    -- filter=120 channel=9
    -15, 4, 10, -3, 22, 29, 15, 34, 26,
    -- filter=120 channel=10
    -4, -1, 2, -7, 0, -8, 0, 3, 5,
    -- filter=120 channel=11
    -9, -24, 1, -17, -13, 7, -12, 3, 23,
    -- filter=120 channel=12
    8, -5, -6, -4, 0, -1, -3, 7, -7,
    -- filter=120 channel=13
    -22, 0, -9, -6, 1, 9, 12, 4, 7,
    -- filter=120 channel=14
    -10, 7, -6, -8, 5, 6, -5, -12, 0,
    -- filter=120 channel=15
    -24, -2, 16, -15, 18, 38, 9, 9, 20,
    -- filter=120 channel=16
    -38, -10, 10, -14, -2, 45, 3, 15, 43,
    -- filter=120 channel=17
    -20, -8, 7, -15, -5, 9, -6, 7, 12,
    -- filter=120 channel=18
    -7, 8, -6, 9, -1, -1, -1, 4, -11,
    -- filter=120 channel=19
    1, -10, 4, -2, 5, 6, 0, 10, 15,
    -- filter=120 channel=20
    4, 3, -7, 5, 19, 5, 15, -2, -1,
    -- filter=120 channel=21
    3, -2, -3, 12, -7, 5, 7, 3, -10,
    -- filter=120 channel=22
    8, -5, 1, -3, -4, 6, -5, -5, -10,
    -- filter=120 channel=23
    6, -5, 4, -13, -3, -3, -11, -2, 1,
    -- filter=120 channel=24
    -20, -23, -11, -8, -12, 15, -17, 4, 10,
    -- filter=120 channel=25
    -21, 0, 26, -8, 10, 23, 6, 1, 21,
    -- filter=120 channel=26
    -6, 0, -6, -4, 11, 0, -5, 4, 10,
    -- filter=120 channel=27
    -21, -14, 23, -18, 2, 21, 1, 9, 21,
    -- filter=120 channel=28
    -18, -23, 7, -16, 1, 14, -12, 3, 5,
    -- filter=120 channel=29
    -19, -8, 10, -8, 19, 44, 5, 25, 35,
    -- filter=120 channel=30
    -3, -6, -18, -18, -24, -24, -13, -14, -19,
    -- filter=120 channel=31
    2, -1, 10, 0, -4, 3, 5, -1, 7,
    -- filter=120 channel=32
    -6, -7, 10, 2, -3, -1, -13, -8, -3,
    -- filter=120 channel=33
    2, -3, 5, 6, 0, -4, 9, 6, -6,
    -- filter=120 channel=34
    -7, -5, -1, 8, 2, 5, 2, 7, -3,
    -- filter=120 channel=35
    -11, 6, 9, -13, -2, 21, -13, -19, -2,
    -- filter=120 channel=36
    12, 7, 6, 12, 8, 1, 6, -2, -5,
    -- filter=120 channel=37
    -1, -2, -7, -9, 14, 13, -6, 7, 24,
    -- filter=120 channel=38
    -31, -10, 17, -27, 0, 31, -11, 7, 25,
    -- filter=120 channel=39
    10, -7, -1, -5, -4, 7, -6, -3, 10,
    -- filter=120 channel=40
    -9, -3, -2, -8, 2, 0, -3, -5, 1,
    -- filter=120 channel=41
    -28, -6, 9, 0, 18, 40, 5, 1, 31,
    -- filter=120 channel=42
    -1, -5, 10, 9, -4, 10, 10, 6, 6,
    -- filter=120 channel=43
    -9, -20, -40, -23, -17, -34, 1, -18, -12,
    -- filter=120 channel=44
    -10, -9, -1, -8, -2, 4, 2, -2, -6,
    -- filter=120 channel=45
    -1, 1, -6, 2, 2, 7, 0, -1, 1,
    -- filter=120 channel=46
    0, 1, 5, 16, 1, 0, 16, 9, 8,
    -- filter=120 channel=47
    1, 4, 1, -8, -7, -4, -8, -9, 4,
    -- filter=120 channel=48
    2, -2, 9, 1, 2, 6, 12, 18, 6,
    -- filter=120 channel=49
    -1, -2, 0, -10, 7, 0, -3, -10, -7,
    -- filter=120 channel=50
    0, -13, -25, -11, -22, -20, 0, -14, -14,
    -- filter=120 channel=51
    0, 7, -2, -3, -11, -2, 4, -3, -3,
    -- filter=120 channel=52
    11, -2, 1, -1, 2, -8, 8, 0, 9,
    -- filter=120 channel=53
    -4, -18, -6, -20, -12, -7, -23, -6, -3,
    -- filter=120 channel=54
    -22, 5, 0, 10, 20, 30, 5, 21, 22,
    -- filter=120 channel=55
    -4, 0, 5, 8, 10, -3, 7, -4, 2,
    -- filter=120 channel=56
    -7, -2, -5, 3, -1, 3, -6, -7, -9,
    -- filter=120 channel=57
    -8, 2, 1, -7, -3, 3, -1, -2, 0,
    -- filter=120 channel=58
    2, 1, 5, 17, 3, -11, 3, -1, -8,
    -- filter=120 channel=59
    -2, 1, 14, 6, 15, 22, 0, 21, 28,
    -- filter=120 channel=60
    -26, -27, 13, -8, 12, 37, 5, 15, 43,
    -- filter=120 channel=61
    -17, -25, -1, -28, -12, 9, -16, 10, 29,
    -- filter=120 channel=62
    -18, -6, 13, -7, -2, 24, 0, 10, 12,
    -- filter=120 channel=63
    -1, -4, 9, 0, 2, -7, 0, -10, 0,
    -- filter=121 channel=0
    0, 9, 10, 10, 5, 13, 9, 10, -3,
    -- filter=121 channel=1
    -13, 0, -11, 2, -10, -2, -3, -2, -16,
    -- filter=121 channel=2
    0, 7, -6, 0, -12, 0, -9, -18, -7,
    -- filter=121 channel=3
    -4, -1, 1, 12, 0, 0, -5, -2, 4,
    -- filter=121 channel=4
    0, 9, -4, 6, -1, 0, -1, -6, -3,
    -- filter=121 channel=5
    0, 7, 3, 0, -2, 12, 6, 16, 3,
    -- filter=121 channel=6
    11, 4, -7, -10, -4, -9, -8, -5, 8,
    -- filter=121 channel=7
    14, 14, 14, 4, 1, -2, 15, 8, 4,
    -- filter=121 channel=8
    6, 21, 2, 7, 2, 1, -2, 7, 2,
    -- filter=121 channel=9
    -1, 6, -16, 7, -5, -12, -5, -2, -16,
    -- filter=121 channel=10
    -8, 1, -1, 4, 1, 0, -3, -2, -4,
    -- filter=121 channel=11
    -5, 13, 0, -3, 7, 0, 3, -8, 4,
    -- filter=121 channel=12
    -8, -1, 4, -4, -9, -1, -4, -8, 0,
    -- filter=121 channel=13
    -2, 2, 1, 8, 2, -5, -7, -4, -2,
    -- filter=121 channel=14
    -1, 9, -1, 11, 15, 1, 14, 15, 8,
    -- filter=121 channel=15
    17, 13, -2, -3, -3, 0, -9, 3, 7,
    -- filter=121 channel=16
    9, 6, -10, 4, 0, -14, -5, -1, -19,
    -- filter=121 channel=17
    -4, 5, -6, 0, 12, 11, 7, 4, 4,
    -- filter=121 channel=18
    -5, -1, 0, 8, 6, 1, -2, 1, 8,
    -- filter=121 channel=19
    -5, 7, -13, -3, 10, -13, -2, -2, 2,
    -- filter=121 channel=20
    2, 9, -2, 5, 5, 15, 7, 7, 5,
    -- filter=121 channel=21
    8, 3, 0, 1, -1, 5, -9, -9, -10,
    -- filter=121 channel=22
    3, -10, -5, 7, -9, 1, -8, -2, 8,
    -- filter=121 channel=23
    3, -2, 3, -3, 8, 11, 7, -2, 0,
    -- filter=121 channel=24
    -6, 16, 12, 5, 9, -1, -3, 14, -8,
    -- filter=121 channel=25
    -13, -8, -17, -2, -5, -7, -14, -20, -12,
    -- filter=121 channel=26
    7, 13, 0, 8, 14, 19, 0, 10, 12,
    -- filter=121 channel=27
    -6, 7, 6, -9, 1, -5, -9, 0, -9,
    -- filter=121 channel=28
    2, 2, 1, 2, 0, -3, 8, 0, -14,
    -- filter=121 channel=29
    18, -1, -8, 1, -8, -12, 1, 1, 1,
    -- filter=121 channel=30
    8, 20, 6, 13, 37, 18, 27, 24, 22,
    -- filter=121 channel=31
    8, 0, -8, -2, 0, -9, -1, 2, 3,
    -- filter=121 channel=32
    -2, -10, 5, -7, 7, 3, -10, -4, -6,
    -- filter=121 channel=33
    -3, 8, 7, 8, -10, 9, -1, 9, -10,
    -- filter=121 channel=34
    6, 13, -3, 12, 2, 13, 6, 2, -2,
    -- filter=121 channel=35
    -3, -3, 2, -4, -5, -13, -11, -5, -12,
    -- filter=121 channel=36
    -5, 5, 7, -2, 6, -1, 7, 3, -4,
    -- filter=121 channel=37
    1, 6, -1, 3, 9, -7, 5, 0, -3,
    -- filter=121 channel=38
    -8, 1, -9, 5, -1, -8, 3, -7, -2,
    -- filter=121 channel=39
    -4, 2, 5, -6, 9, -9, -6, -1, -5,
    -- filter=121 channel=40
    0, -4, 9, -8, 10, -10, -7, 8, 0,
    -- filter=121 channel=41
    14, 16, -5, 13, 6, -7, 5, -11, -4,
    -- filter=121 channel=42
    3, 4, 7, 2, -8, -9, 1, 2, 3,
    -- filter=121 channel=43
    -4, 8, 0, 0, -4, 10, -10, 6, -7,
    -- filter=121 channel=44
    -7, 11, 5, -4, -8, -9, -8, -2, -3,
    -- filter=121 channel=45
    9, 2, -1, 6, -10, -5, 7, 7, 1,
    -- filter=121 channel=46
    13, 18, 12, 0, 4, 1, 0, 18, 1,
    -- filter=121 channel=47
    -3, 3, -2, -5, -6, 5, 8, 9, -6,
    -- filter=121 channel=48
    4, 6, -4, 10, 2, 2, 5, 4, 0,
    -- filter=121 channel=49
    -9, 2, 9, 1, 0, -6, 0, -3, 3,
    -- filter=121 channel=50
    14, 21, 14, 14, 10, 6, 16, 10, 13,
    -- filter=121 channel=51
    7, -6, 7, 4, 2, 12, 0, 10, 5,
    -- filter=121 channel=52
    0, 7, 1, 3, -2, -7, -5, -6, -1,
    -- filter=121 channel=53
    16, 19, 13, 14, 14, 1, 11, 13, 8,
    -- filter=121 channel=54
    -3, 11, -7, 6, 2, -1, 4, -3, -14,
    -- filter=121 channel=55
    0, 0, -9, -6, 4, -8, -1, 7, -3,
    -- filter=121 channel=56
    8, 2, 6, 9, 7, 9, 0, 3, 9,
    -- filter=121 channel=57
    9, -6, -5, 9, -9, 0, 8, 0, 1,
    -- filter=121 channel=58
    9, 0, 5, 0, 4, -7, 2, -3, 7,
    -- filter=121 channel=59
    6, 1, 9, -5, -1, -15, -3, -16, -8,
    -- filter=121 channel=60
    16, 21, 5, 21, 14, 1, -6, 1, 4,
    -- filter=121 channel=61
    6, 17, -4, 13, 19, 10, -5, 8, -4,
    -- filter=121 channel=62
    0, 11, 3, -8, 12, -12, -8, -7, -10,
    -- filter=121 channel=63
    1, 7, -1, 3, -1, 6, -2, -5, 5,
    -- filter=122 channel=0
    13, 18, 12, 15, 35, 19, 21, 21, 23,
    -- filter=122 channel=1
    -26, -15, -14, -22, -11, -18, -6, -9, -12,
    -- filter=122 channel=2
    -13, -15, -13, -18, -28, -6, -14, -14, -17,
    -- filter=122 channel=3
    -25, -14, -3, -22, -17, -10, -12, -14, -7,
    -- filter=122 channel=4
    9, 27, -1, 27, 24, 6, 18, 27, 21,
    -- filter=122 channel=5
    -18, -10, -8, -3, -17, 3, -12, -16, 0,
    -- filter=122 channel=6
    3, 15, 11, 15, 14, 1, 12, 8, 6,
    -- filter=122 channel=7
    -1, 3, 9, 7, -5, 14, -6, 7, 0,
    -- filter=122 channel=8
    3, 18, 0, 31, 36, 13, 4, 11, 4,
    -- filter=122 channel=9
    -37, -49, -69, -49, -69, -78, -39, -71, -66,
    -- filter=122 channel=10
    14, 11, 25, 19, 40, 20, 20, 32, 18,
    -- filter=122 channel=11
    6, 4, 11, 14, 17, 6, -6, 1, 14,
    -- filter=122 channel=12
    -6, -5, 11, 9, 9, -6, -8, -2, 10,
    -- filter=122 channel=13
    5, 8, -4, 8, 9, 9, 17, 9, 0,
    -- filter=122 channel=14
    -8, 11, 3, 7, 2, 13, 0, -6, 11,
    -- filter=122 channel=15
    19, 2, 15, 14, 21, 11, 4, 4, 11,
    -- filter=122 channel=16
    -11, -12, -9, -1, -3, 0, -17, -16, -22,
    -- filter=122 channel=17
    8, 8, 7, 16, 19, 15, 0, 9, 18,
    -- filter=122 channel=18
    35, 33, 26, 40, 39, 21, 21, 33, 18,
    -- filter=122 channel=19
    -19, -26, -16, -31, -24, -18, -14, -37, -20,
    -- filter=122 channel=20
    -10, -19, -8, -9, -14, 0, -10, -9, 3,
    -- filter=122 channel=21
    12, 11, 5, 1, 6, 10, -3, 7, 4,
    -- filter=122 channel=22
    8, -9, 4, -3, 9, -8, -1, -7, -4,
    -- filter=122 channel=23
    11, 21, 31, 25, 32, 32, 7, 26, 28,
    -- filter=122 channel=24
    5, 16, 9, 17, 26, 5, 11, 7, 3,
    -- filter=122 channel=25
    -25, -36, -18, -18, -38, -21, -32, -25, -18,
    -- filter=122 channel=26
    -3, 0, 2, -9, 0, 9, -6, -5, 17,
    -- filter=122 channel=27
    -13, -6, 3, -12, 0, 1, -9, -7, 9,
    -- filter=122 channel=28
    1, -3, 5, -1, 6, -9, -1, -6, -6,
    -- filter=122 channel=29
    -1, -18, -14, 6, -20, -3, -14, -13, -15,
    -- filter=122 channel=30
    -16, 2, 24, -10, 0, 10, -9, -4, 12,
    -- filter=122 channel=31
    3, 0, -1, 0, -2, 11, 2, 3, 7,
    -- filter=122 channel=32
    -16, -10, 1, -16, -18, 5, -16, -11, 2,
    -- filter=122 channel=33
    0, 4, -8, -7, -6, -8, -5, -3, 9,
    -- filter=122 channel=34
    -3, -4, 3, -3, -5, 3, 0, -4, 6,
    -- filter=122 channel=35
    -3, 23, 14, -3, 29, 27, -1, 8, 21,
    -- filter=122 channel=36
    1, 1, 13, 0, 2, -5, 3, -4, 12,
    -- filter=122 channel=37
    -19, -17, -31, -24, -33, -17, -24, -28, -24,
    -- filter=122 channel=38
    2, 1, -13, -2, 15, 6, -10, 2, -6,
    -- filter=122 channel=39
    4, 9, -4, -3, -1, 1, -4, -2, -10,
    -- filter=122 channel=40
    -6, 2, -4, 6, 0, -2, 0, 0, -4,
    -- filter=122 channel=41
    0, 0, 6, 0, 20, 5, -6, 16, 16,
    -- filter=122 channel=42
    -6, -8, -6, -6, 6, 8, 0, 8, 3,
    -- filter=122 channel=43
    -12, -13, 12, -11, -3, 9, 9, 8, 9,
    -- filter=122 channel=44
    -16, -5, -9, -8, -14, -7, -6, -17, -5,
    -- filter=122 channel=45
    7, 3, -9, -7, 8, -2, 8, -8, 8,
    -- filter=122 channel=46
    5, -13, 6, 3, -4, 8, 0, -6, 6,
    -- filter=122 channel=47
    1, 6, 1, 5, 4, -6, 9, -9, 0,
    -- filter=122 channel=48
    0, -13, -2, -2, -8, -6, 0, 0, -3,
    -- filter=122 channel=49
    22, 40, 22, 30, 44, 42, 4, 36, 22,
    -- filter=122 channel=50
    1, 1, 9, -2, -12, 17, 4, -7, 6,
    -- filter=122 channel=51
    30, 37, 38, 40, 56, 43, 32, 46, 31,
    -- filter=122 channel=52
    -7, 5, 8, 9, 3, 0, 5, 0, 3,
    -- filter=122 channel=53
    -14, -15, 17, -11, -14, 4, -7, -2, 16,
    -- filter=122 channel=54
    -28, -53, -60, -43, -52, -54, -33, -44, -45,
    -- filter=122 channel=55
    9, 4, -4, -2, -6, 8, -6, -4, -5,
    -- filter=122 channel=56
    -2, -4, -2, 12, 13, 15, 8, 8, 0,
    -- filter=122 channel=57
    1, 7, -5, 3, -9, -5, 0, -6, 9,
    -- filter=122 channel=58
    -1, 13, 19, 12, 1, 0, 7, 5, 14,
    -- filter=122 channel=59
    -11, -16, 3, -20, -13, -2, -20, 1, -9,
    -- filter=122 channel=60
    22, 21, -3, 29, 33, 27, 16, 36, 21,
    -- filter=122 channel=61
    10, 24, 14, 12, 32, 32, 12, 34, 25,
    -- filter=122 channel=62
    -9, -7, -16, -15, -4, -7, -14, -11, -17,
    -- filter=122 channel=63
    3, 0, -1, -5, 3, -7, 2, 8, -2,
    -- filter=123 channel=0
    -5, -3, 16, -3, -7, 15, -11, -1, 21,
    -- filter=123 channel=1
    -5, 4, -2, -9, -6, 8, 3, -13, 1,
    -- filter=123 channel=2
    4, -10, -8, 2, -3, 3, -2, -16, -2,
    -- filter=123 channel=3
    8, -8, 10, -3, 0, 0, -5, -6, 12,
    -- filter=123 channel=4
    -10, 6, 10, 4, -2, 14, 6, 3, -1,
    -- filter=123 channel=5
    1, -1, 0, 9, 7, 11, 8, 0, 7,
    -- filter=123 channel=6
    6, 1, 3, -5, -5, -1, -14, -10, 10,
    -- filter=123 channel=7
    7, 13, 4, 2, 15, 13, -1, 11, -4,
    -- filter=123 channel=8
    1, 8, 19, -7, -14, 18, 10, 2, 14,
    -- filter=123 channel=9
    9, -1, -17, 7, 6, -10, -4, -11, 0,
    -- filter=123 channel=10
    -5, 1, -4, -5, -1, 8, -14, -7, 2,
    -- filter=123 channel=11
    -11, 0, 9, 6, -4, -6, 0, -8, 10,
    -- filter=123 channel=12
    -1, -3, -10, -7, -5, -6, -2, 5, -2,
    -- filter=123 channel=13
    4, 3, 4, -12, -4, 8, -7, 4, 6,
    -- filter=123 channel=14
    15, 3, 14, -3, -4, 11, 0, 12, 7,
    -- filter=123 channel=15
    -1, 15, 22, -9, -4, 25, -10, -14, 10,
    -- filter=123 channel=16
    -11, 0, -1, -10, 0, 5, -7, -7, 0,
    -- filter=123 channel=17
    -2, 4, 15, -6, -15, -3, 11, -7, 3,
    -- filter=123 channel=18
    -1, -3, 5, -8, 2, 7, 2, -4, 11,
    -- filter=123 channel=19
    -4, 1, -3, 11, 2, 2, 10, -4, -14,
    -- filter=123 channel=20
    -4, 8, -5, 7, 10, 10, 4, 0, -2,
    -- filter=123 channel=21
    0, -5, 1, -7, 8, -6, -6, 4, -8,
    -- filter=123 channel=22
    6, -3, -1, -5, 3, -5, 4, -9, 7,
    -- filter=123 channel=23
    3, -5, 5, -3, 5, -6, 0, 2, 7,
    -- filter=123 channel=24
    -7, 2, 10, 4, -7, 12, 0, -9, 6,
    -- filter=123 channel=25
    2, -3, 7, -9, -4, -5, 0, -17, 6,
    -- filter=123 channel=26
    8, 10, 2, 3, 20, 16, -9, -1, 14,
    -- filter=123 channel=27
    -11, -11, 16, -2, -1, 8, -10, -22, 14,
    -- filter=123 channel=28
    1, 0, 6, 2, -5, -1, 14, -4, 4,
    -- filter=123 channel=29
    -11, 3, 14, -20, -8, 8, 0, -8, 16,
    -- filter=123 channel=30
    11, 18, 24, 22, 21, 28, 27, 26, 8,
    -- filter=123 channel=31
    -4, 5, -5, -4, 7, 0, 4, 10, 6,
    -- filter=123 channel=32
    10, -1, 10, 6, -3, -6, 0, 2, 3,
    -- filter=123 channel=33
    7, 7, 7, -5, -5, -6, -6, -4, -7,
    -- filter=123 channel=34
    -2, 0, 8, 7, 4, 1, 9, 8, 1,
    -- filter=123 channel=35
    -12, -7, 2, -16, -17, 11, 2, -15, 8,
    -- filter=123 channel=36
    -10, -4, 1, -6, 2, 5, -11, 0, 1,
    -- filter=123 channel=37
    2, 10, -7, 0, 3, -6, -6, 0, 1,
    -- filter=123 channel=38
    4, 4, -2, -16, -11, 0, -14, -19, 6,
    -- filter=123 channel=39
    -4, -1, -9, 7, 0, -5, -4, 0, 1,
    -- filter=123 channel=40
    5, 2, -5, -7, -2, 10, -7, 3, -10,
    -- filter=123 channel=41
    -4, 11, 22, -19, -10, 14, -4, -15, 20,
    -- filter=123 channel=42
    -7, -8, 5, 5, 0, 2, 8, 9, -7,
    -- filter=123 channel=43
    13, 10, 0, 14, 0, 6, 0, -3, 4,
    -- filter=123 channel=44
    11, -8, 9, 4, -5, 9, 10, -3, 8,
    -- filter=123 channel=45
    -8, 10, -4, -1, 3, 3, -6, 0, 0,
    -- filter=123 channel=46
    -3, 14, 2, 10, 10, 6, -4, 12, 2,
    -- filter=123 channel=47
    -1, -1, -10, 1, 7, -4, -7, -5, 5,
    -- filter=123 channel=48
    3, -6, 5, -1, -1, 10, 6, 1, 16,
    -- filter=123 channel=49
    -14, -1, 9, -2, -12, 7, -9, -5, -2,
    -- filter=123 channel=50
    7, 12, 17, 17, 8, 14, 0, 13, 3,
    -- filter=123 channel=51
    -7, 7, 7, 7, 0, -3, -14, 0, 0,
    -- filter=123 channel=52
    3, 9, -7, 1, 4, -9, 3, -3, 8,
    -- filter=123 channel=53
    13, 19, 24, 4, 10, 10, 16, 13, 6,
    -- filter=123 channel=54
    -7, 4, -2, -2, 2, -6, 3, 4, 0,
    -- filter=123 channel=55
    -3, 6, 4, -5, 6, 1, 7, 9, -1,
    -- filter=123 channel=56
    0, 6, 9, 7, -4, 3, 6, -4, 0,
    -- filter=123 channel=57
    2, -2, 0, -7, -4, 7, -9, 7, 0,
    -- filter=123 channel=58
    4, 0, -11, 5, 10, 2, -3, 6, -5,
    -- filter=123 channel=59
    -1, -10, 1, -5, -12, 18, -6, -4, 6,
    -- filter=123 channel=60
    -13, 5, 21, -14, 2, 19, -8, -20, 20,
    -- filter=123 channel=61
    8, 11, 8, 2, -3, 14, -10, -15, 7,
    -- filter=123 channel=62
    -1, -2, 4, 5, -6, 3, 3, -8, 0,
    -- filter=123 channel=63
    6, -5, -3, 4, 8, 9, 8, -1, -2,
    -- filter=124 channel=0
    -2, 2, 1, 5, -1, -13, -10, 2, -2,
    -- filter=124 channel=1
    0, -7, 3, 6, -5, -5, 9, -6, -6,
    -- filter=124 channel=2
    -7, 4, 6, 2, 1, 2, -3, 2, -7,
    -- filter=124 channel=3
    2, 0, -2, 9, 0, 10, -3, 0, 13,
    -- filter=124 channel=4
    8, 8, 0, -2, -3, -11, -4, 1, -9,
    -- filter=124 channel=5
    -2, 5, 9, -1, -5, 11, 1, 2, 8,
    -- filter=124 channel=6
    9, 1, -9, -5, 2, 5, -8, 7, -1,
    -- filter=124 channel=7
    0, -1, 6, 1, -6, -8, 6, -1, 5,
    -- filter=124 channel=8
    -6, 9, -6, 0, 0, -5, -3, -3, 4,
    -- filter=124 channel=9
    2, 28, 24, 23, 38, 39, 18, 34, 23,
    -- filter=124 channel=10
    -4, -5, -7, 2, -6, 0, 11, -1, -3,
    -- filter=124 channel=11
    -8, 0, -12, 8, 1, -4, -4, 6, -10,
    -- filter=124 channel=12
    7, -6, -1, 8, 7, 0, -2, 5, 12,
    -- filter=124 channel=13
    11, -4, 0, -2, 2, 0, 6, 0, 1,
    -- filter=124 channel=14
    -6, -1, 9, 10, 10, -6, 0, 9, 8,
    -- filter=124 channel=15
    5, 5, -2, 0, 5, 6, 0, 0, -10,
    -- filter=124 channel=16
    1, 12, -8, -11, 0, 7, -14, 0, -1,
    -- filter=124 channel=17
    -4, -2, 0, -2, -7, 4, 1, -12, 6,
    -- filter=124 channel=18
    13, 0, -6, 5, 5, 10, 15, 11, -3,
    -- filter=124 channel=19
    -4, 8, 13, 14, 2, 0, 15, 17, 7,
    -- filter=124 channel=20
    10, 6, 3, 3, 9, 7, 13, 16, 0,
    -- filter=124 channel=21
    2, 2, 13, 7, 12, -1, 8, -4, -3,
    -- filter=124 channel=22
    -8, 0, 10, -2, -1, 0, -5, -10, 5,
    -- filter=124 channel=23
    4, -3, -7, -12, 0, -14, -4, -11, -8,
    -- filter=124 channel=24
    -2, 9, 1, 6, 7, -7, -7, -5, -3,
    -- filter=124 channel=25
    -11, -6, -2, 0, 6, -9, -14, -13, 0,
    -- filter=124 channel=26
    1, 9, -8, 2, 1, -2, 1, -1, 2,
    -- filter=124 channel=27
    6, -10, 4, -7, -7, -10, -9, -6, -10,
    -- filter=124 channel=28
    -9, 14, 0, 9, 6, 15, 5, -5, 6,
    -- filter=124 channel=29
    -3, 16, 3, 7, 5, 1, -3, 13, 5,
    -- filter=124 channel=30
    -10, -2, 3, 4, -6, 6, -4, 1, 6,
    -- filter=124 channel=31
    1, 5, -1, 11, 6, 2, -4, 0, 10,
    -- filter=124 channel=32
    6, 8, 0, -8, 2, -10, 7, 0, -6,
    -- filter=124 channel=33
    -2, -3, -9, 10, -9, 1, 10, -8, -3,
    -- filter=124 channel=34
    -7, -3, 7, 3, -2, 8, -3, -7, 7,
    -- filter=124 channel=35
    -6, -5, -6, 0, -17, -13, -8, -9, -4,
    -- filter=124 channel=36
    4, -3, 8, -6, -3, -2, 9, -8, 11,
    -- filter=124 channel=37
    4, 8, 8, 2, 8, 8, 0, -1, 1,
    -- filter=124 channel=38
    -9, -6, -5, -11, -7, -8, -3, -10, -13,
    -- filter=124 channel=39
    0, -9, -2, 7, 6, -3, 3, -10, 10,
    -- filter=124 channel=40
    -3, -2, 2, 6, -4, -11, 2, -7, -5,
    -- filter=124 channel=41
    -8, -8, 8, -6, 6, 3, 2, -3, -15,
    -- filter=124 channel=42
    -5, 8, 5, 4, -6, -2, 7, 8, 8,
    -- filter=124 channel=43
    6, 4, 3, 5, -1, 1, -1, -5, 3,
    -- filter=124 channel=44
    7, 2, 2, -9, -2, 9, 1, -4, -5,
    -- filter=124 channel=45
    10, -10, -7, -1, -3, 7, 1, 10, 0,
    -- filter=124 channel=46
    -5, 10, -9, 3, 4, -6, -8, -7, -1,
    -- filter=124 channel=47
    -6, 9, 6, -10, -3, 7, -3, -5, 6,
    -- filter=124 channel=48
    2, 5, 4, 10, 12, 11, -3, 7, 12,
    -- filter=124 channel=49
    0, 4, -1, 2, -9, -6, 4, -13, -7,
    -- filter=124 channel=50
    1, -4, 0, 1, -9, 10, -3, 7, 0,
    -- filter=124 channel=51
    0, 5, 0, -3, 1, -4, -8, -1, -12,
    -- filter=124 channel=52
    6, -6, -4, 8, 2, -7, -5, -1, 4,
    -- filter=124 channel=53
    5, -12, -8, -12, -8, 0, -2, 3, 0,
    -- filter=124 channel=54
    14, 18, 6, 9, 20, 12, -1, 24, 23,
    -- filter=124 channel=55
    4, -9, 10, 0, -1, 0, -5, 0, -8,
    -- filter=124 channel=56
    -8, -9, 0, -9, -5, 0, 3, 7, 5,
    -- filter=124 channel=57
    -9, -5, -4, -7, 8, -7, 3, -10, -1,
    -- filter=124 channel=58
    9, 0, 0, 12, 4, 4, 3, -3, -2,
    -- filter=124 channel=59
    0, 12, 0, 7, 7, 10, 5, -9, 8,
    -- filter=124 channel=60
    2, -4, -6, 5, -5, -10, -14, -13, -11,
    -- filter=124 channel=61
    -3, -9, -4, -8, -7, -4, -14, -1, -2,
    -- filter=124 channel=62
    -5, 10, 10, 0, -4, 1, 8, 7, -5,
    -- filter=124 channel=63
    -1, 8, 2, -6, -1, -7, 8, 0, 10,
    -- filter=125 channel=0
    7, 12, 2, 7, 14, 9, 10, 4, 7,
    -- filter=125 channel=1
    -26, -16, -15, -24, -9, -6, -14, -13, 3,
    -- filter=125 channel=2
    -13, -15, -9, -15, -19, -21, -19, -9, -14,
    -- filter=125 channel=3
    3, -7, -3, 1, 0, 2, -7, 1, 10,
    -- filter=125 channel=4
    -9, 13, 6, -1, 10, 5, 4, 1, 9,
    -- filter=125 channel=5
    10, 5, 8, -3, 0, 7, -6, 9, 3,
    -- filter=125 channel=6
    -6, -3, 5, -9, -1, 6, 1, 3, -1,
    -- filter=125 channel=7
    -6, -1, 2, -10, 4, 2, 4, -7, 2,
    -- filter=125 channel=8
    0, 16, -8, 13, 12, 3, 10, 18, 10,
    -- filter=125 channel=9
    0, -8, -14, 1, -1, -2, -4, -9, 2,
    -- filter=125 channel=10
    4, -4, 1, -11, 7, 1, 2, 6, -1,
    -- filter=125 channel=11
    -15, 5, 2, -16, 3, 13, -8, 13, 12,
    -- filter=125 channel=12
    10, 9, 1, 11, -3, -6, 7, 9, 6,
    -- filter=125 channel=13
    3, 3, -14, 13, 12, -8, 8, 5, -1,
    -- filter=125 channel=14
    2, 9, 9, -10, -1, 0, -2, 2, 13,
    -- filter=125 channel=15
    -5, 7, -9, 15, 29, 4, 11, 21, 10,
    -- filter=125 channel=16
    -13, -2, -24, 4, 6, -12, 6, 15, 5,
    -- filter=125 channel=17
    -12, 0, 6, 0, 23, 12, 7, 24, 20,
    -- filter=125 channel=18
    -2, 4, 10, 15, 25, 4, 5, 6, -6,
    -- filter=125 channel=19
    -15, -20, -8, -9, -12, -15, -14, -10, -14,
    -- filter=125 channel=20
    -12, -5, -14, -10, -5, -4, -6, -13, -14,
    -- filter=125 channel=21
    0, 1, -5, 2, -5, -1, -5, 4, 5,
    -- filter=125 channel=22
    -4, 3, -9, -2, 7, 0, -3, -2, 3,
    -- filter=125 channel=23
    -6, -6, -4, -5, -4, 1, 2, 11, 6,
    -- filter=125 channel=24
    -6, -1, -1, 4, 17, 4, 7, 13, 15,
    -- filter=125 channel=25
    -9, -19, -16, -24, -8, -22, -5, -6, -12,
    -- filter=125 channel=26
    3, 3, -9, -10, 2, -16, -6, 1, -4,
    -- filter=125 channel=27
    -2, 3, -12, 0, 1, 4, -12, 9, 4,
    -- filter=125 channel=28
    1, 9, -6, -8, 5, 11, -3, 7, 9,
    -- filter=125 channel=29
    -10, 8, -6, 7, 14, 0, 17, 19, 0,
    -- filter=125 channel=30
    -9, -16, -4, -20, -6, -7, -5, -15, 8,
    -- filter=125 channel=31
    -3, -4, 0, 6, 9, 6, 4, -6, 2,
    -- filter=125 channel=32
    -12, -11, -1, -26, -14, -12, -18, -18, 2,
    -- filter=125 channel=33
    -8, 7, 6, 6, -4, 0, -2, 9, 3,
    -- filter=125 channel=34
    7, 1, -2, 7, 5, -3, -3, -1, -2,
    -- filter=125 channel=35
    -17, -5, 0, -22, -13, 2, -14, -5, 8,
    -- filter=125 channel=36
    8, 10, 12, 4, -8, 4, 8, 3, -3,
    -- filter=125 channel=37
    -7, -15, -10, -10, 3, 0, 0, 9, 7,
    -- filter=125 channel=38
    -5, 5, -12, 0, -2, -10, 0, 5, 13,
    -- filter=125 channel=39
    -9, -3, -3, -8, 2, -5, 6, 10, -7,
    -- filter=125 channel=40
    -10, -4, -9, 3, -11, -2, -8, 4, -4,
    -- filter=125 channel=41
    -4, 14, 3, -4, 9, 2, -2, 14, 8,
    -- filter=125 channel=42
    -7, -6, -8, -8, -1, 6, -3, 1, 6,
    -- filter=125 channel=43
    -33, -49, -24, -32, -36, -25, -22, -23, -22,
    -- filter=125 channel=44
    -11, -5, 0, -16, -5, -3, -23, -17, -7,
    -- filter=125 channel=45
    8, -7, 6, 0, -3, -7, 1, 10, -5,
    -- filter=125 channel=46
    0, 6, -2, 0, 2, -11, 12, 10, -11,
    -- filter=125 channel=47
    -2, -6, 4, -7, 9, 10, 0, -4, -7,
    -- filter=125 channel=48
    3, 0, 4, 14, 4, -8, 4, -6, 6,
    -- filter=125 channel=49
    -1, 22, 4, 11, 7, 17, 4, 9, 16,
    -- filter=125 channel=50
    -3, -6, -15, -16, -13, -11, -14, -13, -8,
    -- filter=125 channel=51
    2, 15, 10, 5, 5, 4, -3, 16, 6,
    -- filter=125 channel=52
    -8, -6, -2, -9, 5, -1, 7, 2, 2,
    -- filter=125 channel=53
    -19, -11, -3, -8, -25, 1, -19, -11, -3,
    -- filter=125 channel=54
    -15, -8, 0, -6, 7, 0, 5, -4, 4,
    -- filter=125 channel=55
    1, 9, 5, -1, -7, -5, 0, 0, 9,
    -- filter=125 channel=56
    5, -3, 5, -5, -9, -3, -5, 11, 5,
    -- filter=125 channel=57
    7, 9, -8, 8, 5, -7, -5, 0, 9,
    -- filter=125 channel=58
    1, -1, -3, 0, -7, 8, 6, 0, 3,
    -- filter=125 channel=59
    -5, -9, -14, 10, -3, 3, 0, 12, 11,
    -- filter=125 channel=60
    -2, 8, -8, 8, 39, 2, 20, 31, 4,
    -- filter=125 channel=61
    -14, -2, 1, 11, 15, 15, 2, 30, 14,
    -- filter=125 channel=62
    -7, 3, -1, -5, 7, 1, -12, -4, -4,
    -- filter=125 channel=63
    6, 9, -2, -9, 2, 0, -3, -1, 0,
    -- filter=126 channel=0
    10, -5, 3, 3, 3, -8, 5, -5, -10,
    -- filter=126 channel=1
    4, 3, 6, -2, 16, 1, 4, 11, -4,
    -- filter=126 channel=2
    16, -1, 3, 0, -12, -18, 3, -14, -14,
    -- filter=126 channel=3
    26, 2, 0, 12, 13, -7, -1, 2, -12,
    -- filter=126 channel=4
    -2, 15, 5, -5, -6, -11, 8, -11, -7,
    -- filter=126 channel=5
    17, 0, -1, 10, 11, -9, -1, -2, -11,
    -- filter=126 channel=6
    -3, 3, 0, 5, -5, -11, 5, -4, -15,
    -- filter=126 channel=7
    -6, 3, -9, 5, -4, -10, 1, 12, 10,
    -- filter=126 channel=8
    19, 24, 1, 5, 1, -1, -6, -15, -20,
    -- filter=126 channel=9
    23, 8, -2, 9, 15, -6, -7, 6, -4,
    -- filter=126 channel=10
    -15, -12, 6, 6, -10, 6, 1, 4, 13,
    -- filter=126 channel=11
    11, 18, 4, 13, 15, -6, -4, -2, -3,
    -- filter=126 channel=12
    -4, -2, -7, 11, -7, 3, -2, 2, -3,
    -- filter=126 channel=13
    11, 3, 2, 11, 3, -7, 2, -16, -23,
    -- filter=126 channel=14
    6, -3, 2, -1, 4, 4, 4, -2, 7,
    -- filter=126 channel=15
    21, 8, 2, 9, -1, -11, -6, -13, -20,
    -- filter=126 channel=16
    21, 7, 7, 6, -8, -18, -6, -13, -39,
    -- filter=126 channel=17
    22, 6, 2, 3, 11, 0, 7, 10, -10,
    -- filter=126 channel=18
    -2, 5, -4, -2, 0, -8, 4, -2, 0,
    -- filter=126 channel=19
    11, 18, -8, 1, 16, -14, 6, 3, 0,
    -- filter=126 channel=20
    5, 0, -11, 2, 0, 0, -10, 2, -10,
    -- filter=126 channel=21
    3, -10, 9, -6, -7, -2, 11, 7, -6,
    -- filter=126 channel=22
    -8, -4, 1, 10, 5, -9, 3, 8, 3,
    -- filter=126 channel=23
    -6, 4, 7, -11, 2, 0, -8, 3, 10,
    -- filter=126 channel=24
    19, 2, 11, 2, 9, -1, -2, 5, -5,
    -- filter=126 channel=25
    18, 2, -12, 5, 4, -8, -4, 0, -15,
    -- filter=126 channel=26
    9, -11, -4, 7, -5, 1, 6, 3, 4,
    -- filter=126 channel=27
    8, 17, 6, 13, 12, -13, 12, -3, -15,
    -- filter=126 channel=28
    21, 0, -2, 6, 0, -15, -11, 1, -18,
    -- filter=126 channel=29
    23, 0, -9, 22, -5, -17, -7, -19, -44,
    -- filter=126 channel=30
    14, 9, -4, 10, 10, 0, 0, 13, 10,
    -- filter=126 channel=31
    0, 0, -3, 1, -7, 1, -5, 9, 6,
    -- filter=126 channel=32
    2, 10, -2, 0, 10, 16, 9, 11, 9,
    -- filter=126 channel=33
    3, 3, 3, -5, 5, -9, -8, -1, -10,
    -- filter=126 channel=34
    6, -6, 4, 1, -2, -2, -9, 5, 4,
    -- filter=126 channel=35
    1, 9, -2, -3, 4, 0, -8, 5, 3,
    -- filter=126 channel=36
    2, -7, -5, -1, 0, 11, 0, 3, 1,
    -- filter=126 channel=37
    10, 15, 2, 20, 1, 6, 4, 2, 3,
    -- filter=126 channel=38
    9, 13, -2, 21, 0, -12, 10, -12, -9,
    -- filter=126 channel=39
    -7, -1, 1, -5, 4, 9, 0, -9, 6,
    -- filter=126 channel=40
    11, 7, -6, 9, -4, 0, 0, -5, -8,
    -- filter=126 channel=41
    36, 10, -7, 14, 2, -24, -10, -4, -29,
    -- filter=126 channel=42
    4, 7, 8, -10, -3, -8, -9, 0, 8,
    -- filter=126 channel=43
    -2, -15, -6, -4, -2, -4, -6, 3, -5,
    -- filter=126 channel=44
    8, 7, -4, 2, 0, 8, -2, -2, -3,
    -- filter=126 channel=45
    5, 3, 3, -5, 2, 4, 0, 8, 0,
    -- filter=126 channel=46
    9, -10, -4, -5, -5, -2, 8, -10, 3,
    -- filter=126 channel=47
    0, -6, 0, -5, -7, -4, 10, 1, -1,
    -- filter=126 channel=48
    17, -7, -3, -1, 0, -9, 4, -1, -7,
    -- filter=126 channel=49
    -1, 0, -8, -3, -7, 2, 6, -1, 1,
    -- filter=126 channel=50
    -2, 8, -8, 14, 0, 1, 8, 0, 1,
    -- filter=126 channel=51
    -9, -10, 0, -5, -5, 8, 1, -5, 11,
    -- filter=126 channel=52
    8, 7, -6, 5, 5, -7, 9, -1, -2,
    -- filter=126 channel=53
    11, 1, -4, 5, 16, 15, 14, 2, 13,
    -- filter=126 channel=54
    16, 21, 10, 3, 19, -8, 13, -4, -16,
    -- filter=126 channel=55
    9, 6, -6, -9, -2, 9, -4, -3, -5,
    -- filter=126 channel=56
    1, 5, 4, 10, -4, 6, 12, -8, -9,
    -- filter=126 channel=57
    -10, -7, -7, 0, -3, 7, 7, -5, 6,
    -- filter=126 channel=58
    -3, -13, 0, 5, 0, -8, -11, -11, -4,
    -- filter=126 channel=59
    31, 18, 2, 19, 8, 2, 1, -8, -19,
    -- filter=126 channel=60
    37, 17, 1, 19, 0, -8, 10, -4, -17,
    -- filter=126 channel=61
    11, 17, 0, 19, 20, -13, -8, -7, -11,
    -- filter=126 channel=62
    24, 14, 4, 1, 1, -8, -4, 12, -2,
    -- filter=126 channel=63
    0, 4, -4, 10, 9, 3, -2, -6, 7,
    -- filter=127 channel=0
    -4, -5, 6, -4, -1, -3, 0, -11, -1,
    -- filter=127 channel=1
    3, 6, -11, -8, 0, 1, -9, -7, -10,
    -- filter=127 channel=2
    -7, -6, 9, 9, -9, -10, 2, -7, 7,
    -- filter=127 channel=3
    -4, -2, -6, 5, -1, -9, -5, 0, -6,
    -- filter=127 channel=4
    -9, -2, 0, 6, 8, -2, -7, 5, -9,
    -- filter=127 channel=5
    -5, 1, -12, -6, 15, 6, 6, 0, -6,
    -- filter=127 channel=6
    7, -1, 6, 12, -5, 5, 11, -2, -10,
    -- filter=127 channel=7
    8, 8, -9, 0, 8, -4, 10, 0, 6,
    -- filter=127 channel=8
    -4, -2, -10, 8, 6, -16, 6, -1, -13,
    -- filter=127 channel=9
    -5, 3, 0, 10, -8, -1, 2, -9, 11,
    -- filter=127 channel=10
    0, -1, -3, 3, 5, 10, -2, 4, 5,
    -- filter=127 channel=11
    10, 14, -6, -3, 7, -11, 11, -3, -14,
    -- filter=127 channel=12
    7, 10, 0, 0, 6, -6, -10, 2, 2,
    -- filter=127 channel=13
    -5, 2, -8, -5, 2, 9, 7, 3, -4,
    -- filter=127 channel=14
    12, 4, 9, 1, 10, 3, 6, -1, 0,
    -- filter=127 channel=15
    13, 5, 7, 3, -14, 8, 17, -2, 6,
    -- filter=127 channel=16
    2, -4, -6, 15, -5, -7, 12, 2, -5,
    -- filter=127 channel=17
    -6, 4, -10, -7, 9, 3, 6, 0, -15,
    -- filter=127 channel=18
    -4, 6, -6, -2, 5, 8, -8, -3, -4,
    -- filter=127 channel=19
    -1, 0, 3, -8, 7, -2, 4, -3, -9,
    -- filter=127 channel=20
    0, 0, 4, 13, -6, -3, 12, -9, -3,
    -- filter=127 channel=21
    2, 6, 4, 0, -7, 6, -4, 5, 0,
    -- filter=127 channel=22
    -7, -7, 0, -4, 4, 5, -1, 6, 6,
    -- filter=127 channel=23
    -7, 8, 2, 4, -1, -12, 2, 11, 2,
    -- filter=127 channel=24
    3, -3, 2, -8, -3, -2, 2, -4, -10,
    -- filter=127 channel=25
    -5, 2, 2, -1, -13, 0, 8, -11, 6,
    -- filter=127 channel=26
    5, -1, -3, 12, -2, -4, 10, 9, 0,
    -- filter=127 channel=27
    -4, 8, -8, -6, 2, -10, -3, -9, -8,
    -- filter=127 channel=28
    -4, -6, 2, 6, -8, -12, 0, -6, -8,
    -- filter=127 channel=29
    -1, -6, 0, 12, -7, -4, 14, -9, 2,
    -- filter=127 channel=30
    13, 16, 0, 12, 13, 0, 10, 28, -2,
    -- filter=127 channel=31
    -10, 7, -4, -2, 9, 2, -2, 6, 8,
    -- filter=127 channel=32
    0, -7, -5, -7, 13, 0, 0, 2, -9,
    -- filter=127 channel=33
    1, -1, -2, 7, -3, 9, -9, 2, 5,
    -- filter=127 channel=34
    4, 5, 10, 0, -2, 6, 5, -4, -5,
    -- filter=127 channel=35
    2, -9, -5, 3, 6, 7, 12, -2, 6,
    -- filter=127 channel=36
    1, -4, 6, -6, 4, 6, 0, -3, -10,
    -- filter=127 channel=37
    -4, -1, 9, -7, 10, 8, 6, 3, -5,
    -- filter=127 channel=38
    -1, 11, -8, 14, -2, -11, 10, -6, -4,
    -- filter=127 channel=39
    8, -10, -8, -5, 1, -7, 10, -8, 5,
    -- filter=127 channel=40
    7, 4, -9, 0, 6, -4, 10, 0, -1,
    -- filter=127 channel=41
    12, 9, -4, 15, -8, -5, 4, 4, -3,
    -- filter=127 channel=42
    4, 1, 3, -9, -6, 8, -8, 6, -5,
    -- filter=127 channel=43
    -9, -4, 2, -12, -2, 9, -2, -4, -1,
    -- filter=127 channel=44
    -3, 9, 3, -3, 11, -13, -4, 9, -1,
    -- filter=127 channel=45
    -2, 7, -2, 0, -7, 0, -9, -2, -7,
    -- filter=127 channel=46
    16, -6, 0, 2, -8, 0, 1, 10, 5,
    -- filter=127 channel=47
    0, -6, 8, -8, 5, 8, -6, -7, -10,
    -- filter=127 channel=48
    2, 1, -1, -5, -6, 5, -5, -4, -6,
    -- filter=127 channel=49
    0, 6, 4, -1, 1, -2, -7, -8, 4,
    -- filter=127 channel=50
    7, 10, -9, -5, 13, -3, -3, 1, 3,
    -- filter=127 channel=51
    -8, -3, 2, -8, 6, -2, -10, 6, 8,
    -- filter=127 channel=52
    5, 3, -4, -8, 2, -5, -3, -2, 5,
    -- filter=127 channel=53
    -1, 11, 4, 3, 12, 7, -7, 15, -5,
    -- filter=127 channel=54
    4, 12, -5, -3, -6, 6, 0, 5, 3,
    -- filter=127 channel=55
    9, 5, -1, -10, 4, -4, 1, 3, 7,
    -- filter=127 channel=56
    3, 10, 6, -8, 7, -6, 1, -7, -2,
    -- filter=127 channel=57
    -3, -3, -8, 1, 0, -6, 0, -9, 1,
    -- filter=127 channel=58
    9, 1, -7, 2, -12, -8, 2, -12, 7,
    -- filter=127 channel=59
    5, -4, 5, 16, -9, -8, 0, -8, 5,
    -- filter=127 channel=60
    14, -5, 0, 18, -5, -3, 14, -7, 1,
    -- filter=127 channel=61
    5, 3, -6, -6, 0, -2, 14, -1, -12,
    -- filter=127 channel=62
    -2, 11, 5, 8, 5, -10, -6, 12, -7,
    -- filter=127 channel=63
    -1, -6, 5, -9, -2, -7, 7, -9, 6,

    -- ifmap
    -- channel=0
    234, 234, 239, 238, 237, 225, 247, 258, 240, 209, 183, 193, 199, 202, 201, 
    236, 241, 247, 244, 249, 228, 206, 211, 169, 130, 76, 82, 128, 190, 202, 
    164, 236, 247, 248, 255, 246, 143, 100, 86, 124, 74, 72, 51, 114, 191, 
    33, 157, 235, 251, 204, 182, 120, 68, 69, 156, 82, 88, 54, 40, 179, 
    41, 137, 193, 260, 170, 123, 88, 55, 50, 137, 105, 52, 75, 36, 91, 
    48, 135, 181, 178, 199, 139, 106, 78, 25, 196, 93, 51, 92, 58, 34, 
    48, 84, 170, 172, 182, 171, 152, 95, 47, 191, 73, 47, 69, 86, 67, 
    65, 87, 74, 148, 168, 210, 90, 109, 79, 187, 99, 48, 86, 103, 132, 
    72, 110, 11, 130, 106, 124, 98, 86, 119, 116, 128, 51, 79, 138, 195, 
    127, 117, 24, 107, 70, 85, 126, 94, 69, 121, 52, 40, 92, 196, 201, 
    151, 117, 34, 188, 50, 49, 120, 101, 30, 18, 4, 3, 12, 63, 48, 
    74, 117, 91, 219, 63, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 54, 139, 141, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 102, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    47, 65, 51, 50, 40, 60, 57, 51, 43, 53, 67, 69, 64, 54, 45, 
    39, 64, 51, 53, 43, 50, 49, 73, 83, 44, 35, 43, 55, 55, 48, 
    82, 62, 48, 52, 41, 88, 78, 51, 35, 35, 68, 52, 43, 35, 61, 
    68, 0, 49, 45, 60, 32, 58, 43, 40, 46, 88, 67, 66, 40, 38, 
    65, 27, 50, 3, 84, 48, 106, 74, 65, 1, 64, 62, 46, 46, 17, 
    62, 86, 75, 56, 156, 118, 112, 63, 62, 0, 98, 83, 50, 45, 30, 
    53, 107, 78, 93, 64, 57, 123, 74, 88, 22, 100, 60, 33, 38, 48, 
    73, 110, 15, 67, 11, 101, 120, 90, 86, 42, 89, 71, 47, 70, 53, 
    93, 96, 76, 70, 42, 85, 76, 56, 32, 40, 93, 95, 51, 44, 35, 
    108, 84, 109, 32, 100, 44, 37, 78, 41, 106, 86, 47, 34, 39, 55, 
    92, 88, 110, 11, 64, 32, 66, 136, 102, 38, 12, 9, 10, 18, 21, 
    65, 97, 80, 43, 170, 103, 68, 69, 52, 28, 25, 27, 28, 22, 35, 
    9, 48, 41, 136, 120, 39, 42, 35, 24, 16, 12, 17, 34, 33, 14, 
    26, 22, 32, 177, 49, 27, 30, 35, 35, 31, 24, 36, 24, 12, 59, 
    36, 32, 27, 78, 27, 35, 45, 37, 25, 23, 29, 16, 0, 29, 36, 
    
    -- channel=2
    132, 151, 150, 146, 139, 154, 149, 142, 135, 114, 106, 120, 140, 133, 117, 
    134, 163, 156, 147, 153, 241, 155, 139, 103, 132, 140, 112, 96, 104, 120, 
    95, 99, 145, 146, 141, 142, 110, 80, 101, 198, 166, 149, 111, 61, 127, 
    112, 140, 138, 151, 152, 152, 185, 126, 110, 156, 171, 124, 97, 52, 104, 
    182, 234, 152, 197, 335, 292, 210, 142, 88, 168, 212, 146, 129, 91, 69, 
    178, 224, 167, 161, 213, 237, 255, 167, 113, 246, 212, 116, 124, 120, 108, 
    206, 219, 116, 137, 180, 258, 237, 204, 124, 251, 181, 131, 123, 147, 123, 
    247, 259, 147, 154, 167, 267, 193, 146, 119, 216, 178, 116, 122, 137, 121, 
    273, 275, 159, 190, 164, 139, 138, 153, 145, 159, 106, 69, 90, 133, 157, 
    257, 261, 178, 227, 150, 148, 201, 245, 146, 107, 70, 59, 119, 171, 135, 
    250, 265, 176, 327, 341, 224, 251, 215, 138, 112, 95, 131, 129, 104, 85, 
    119, 228, 232, 381, 197, 68, 96, 95, 80, 90, 96, 109, 121, 121, 113, 
    92, 119, 245, 302, 86, 119, 112, 105, 95, 99, 114, 128, 122, 121, 155, 
    92, 103, 174, 177, 95, 123, 118, 106, 111, 119, 111, 98, 103, 132, 96, 
    110, 111, 109, 66, 60, 73, 84, 111, 140, 145, 110, 107, 175, 168, 81, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 67, 0, 0, 96, 40, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 89, 0, 0, 111, 29, 42, 0, 0, 89, 19, 0, 0, 0, 0, 
    0, 77, 0, 0, 17, 73, 78, 0, 0, 112, 0, 0, 0, 0, 0, 
    45, 60, 0, 0, 0, 136, 0, 0, 0, 69, 0, 0, 0, 0, 0, 
    82, 109, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    97, 107, 0, 50, 0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 
    125, 97, 0, 167, 91, 10, 92, 55, 0, 0, 0, 0, 0, 0, 0, 
    49, 91, 34, 259, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 30, 92, 194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 87, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 20, 0, 
    
    -- channel=4
    123, 115, 120, 123, 123, 114, 126, 126, 119, 111, 97, 96, 100, 106, 103, 
    120, 117, 120, 126, 122, 137, 130, 113, 85, 73, 84, 79, 76, 95, 108, 
    101, 97, 130, 124, 131, 112, 98, 59, 63, 84, 101, 75, 79, 72, 94, 
    85, 93, 135, 122, 122, 93, 107, 82, 77, 82, 104, 82, 64, 60, 67, 
    100, 131, 142, 98, 145, 132, 108, 82, 65, 64, 108, 94, 70, 60, 61, 
    122, 134, 145, 132, 93, 109, 128, 88, 75, 93, 141, 82, 69, 68, 59, 
    117, 140, 110, 106, 79, 129, 139, 119, 78, 105, 121, 87, 72, 79, 89, 
    137, 115, 107, 111, 97, 138, 127, 95, 84, 111, 114, 84, 65, 94, 88, 
    146, 132, 128, 96, 132, 78, 89, 95, 82, 112, 91, 60, 54, 80, 118, 
    141, 140, 118, 86, 104, 84, 82, 121, 109, 84, 58, 28, 59, 114, 115, 
    126, 143, 115, 117, 171, 126, 129, 117, 90, 57, 48, 59, 71, 89, 92, 
    88, 118, 121, 185, 173, 74, 60, 56, 56, 58, 63, 61, 65, 72, 68, 
    82, 85, 114, 198, 77, 60, 59, 57, 58, 60, 60, 71, 74, 66, 75, 
    69, 64, 97, 136, 76, 63, 66, 58, 53, 59, 66, 67, 62, 74, 91, 
    76, 56, 76, 54, 64, 57, 59, 60, 65, 71, 70, 58, 75, 97, 63, 
    
    -- channel=5
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 0, 2, 0, 29, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 27, 14, 0, 0, 41, 24, 44, 0, 0, 
    122, 0, 0, 0, 0, 0, 27, 35, 9, 0, 63, 7, 35, 16, 0, 
    147, 0, 20, 0, 51, 41, 72, 50, 18, 0, 43, 77, 1, 47, 0, 
    111, 0, 40, 0, 0, 34, 73, 59, 71, 0, 92, 82, 0, 34, 28, 
    112, 56, 0, 32, 0, 0, 50, 63, 90, 0, 112, 62, 0, 0, 34, 
    96, 76, 58, 34, 0, 0, 96, 10, 46, 0, 61, 65, 0, 0, 0, 
    106, 33, 135, 0, 27, 0, 36, 16, 0, 19, 0, 54, 0, 0, 0, 
    43, 31, 148, 0, 86, 2, 0, 63, 23, 5, 53, 7, 0, 0, 0, 
    0, 40, 137, 0, 179, 94, 0, 55, 113, 57, 25, 20, 13, 3, 41, 
    0, 0, 86, 0, 172, 97, 21, 22, 50, 30, 31, 29, 36, 38, 56, 
    69, 0, 0, 52, 179, 39, 43, 33, 38, 34, 35, 39, 46, 45, 43, 
    84, 38, 0, 114, 78, 31, 57, 39, 31, 35, 40, 40, 53, 25, 61, 
    90, 42, 23, 31, 45, 9, 25, 37, 31, 45, 61, 35, 11, 84, 112, 
    
    -- channel=6
    134, 134, 137, 136, 137, 139, 138, 139, 135, 123, 114, 119, 126, 124, 118, 
    133, 143, 141, 138, 143, 162, 138, 130, 109, 114, 108, 104, 108, 117, 122, 
    103, 131, 142, 139, 142, 136, 98, 98, 95, 129, 91, 88, 79, 96, 119, 
    77, 142, 139, 144, 131, 140, 119, 86, 82, 121, 90, 88, 66, 59, 119, 
    90, 149, 131, 171, 172, 161, 108, 79, 66, 132, 122, 85, 88, 63, 94, 
    99, 126, 124, 130, 125, 122, 115, 96, 67, 168, 109, 70, 91, 79, 78, 
    106, 108, 114, 104, 135, 150, 124, 112, 67, 168, 93, 80, 92, 98, 83, 
    119, 115, 113, 124, 137, 151, 97, 92, 76, 143, 93, 74, 89, 95, 90, 
    123, 136, 77, 114, 118, 106, 93, 96, 111, 130, 88, 52, 83, 102, 128, 
    122, 130, 70, 141, 83, 103, 131, 121, 103, 72, 57, 61, 98, 135, 124, 
    143, 137, 81, 184, 128, 116, 136, 100, 66, 81, 76, 82, 90, 112, 101, 
    97, 124, 114, 206, 85, 43, 70, 66, 50, 62, 58, 64, 63, 61, 53, 
    50, 93, 146, 145, 34, 59, 56, 56, 53, 55, 61, 64, 59, 61, 74, 
    38, 58, 128, 67, 51, 66, 58, 55, 56, 58, 57, 49, 50, 63, 45, 
    40, 47, 64, 54, 48, 49, 47, 55, 67, 68, 51, 55, 84, 66, 28, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 0, 3, 10, 5, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 30, 5, 22, 0, 7, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 31, 15, 5, 0, 22, 3, 27, 0, 0, 
    89, 0, 0, 0, 6, 0, 10, 33, 0, 0, 29, 9, 23, 21, 0, 
    93, 0, 32, 0, 0, 19, 38, 33, 9, 0, 9, 60, 0, 30, 0, 
    89, 0, 42, 18, 0, 26, 19, 35, 39, 0, 56, 61, 0, 17, 18, 
    87, 0, 1, 44, 0, 0, 9, 26, 60, 0, 69, 41, 0, 0, 23, 
    65, 0, 42, 11, 0, 0, 58, 0, 30, 0, 32, 45, 0, 0, 0, 
    52, 0, 101, 0, 34, 0, 16, 0, 0, 0, 0, 43, 0, 0, 0, 
    0, 0, 89, 0, 67, 4, 0, 5, 19, 16, 35, 5, 0, 0, 6, 
    0, 0, 75, 0, 75, 62, 0, 6, 66, 19, 0, 0, 0, 0, 12, 
    0, 0, 34, 0, 113, 53, 0, 0, 14, 0, 0, 0, 0, 0, 4, 
    10, 0, 0, 0, 123, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 20, 37, 0, 7, 1, 0, 0, 0, 0, 0, 0, 8, 
    25, 0, 0, 0, 11, 0, 0, 0, 0, 0, 11, 0, 0, 9, 44, 
    
    -- channel=8
    293, 295, 297, 305, 299, 293, 309, 307, 294, 276, 246, 244, 255, 259, 242, 
    291, 298, 304, 313, 307, 386, 331, 291, 219, 209, 231, 197, 187, 233, 258, 
    250, 246, 309, 306, 306, 314, 249, 162, 155, 250, 286, 234, 201, 158, 236, 
    242, 216, 319, 310, 307, 257, 305, 210, 189, 239, 299, 211, 167, 119, 175, 
    339, 378, 348, 319, 510, 393, 338, 221, 155, 178, 342, 251, 193, 157, 111, 
    342, 414, 370, 247, 341, 358, 402, 274, 195, 268, 402, 233, 202, 194, 147, 
    349, 403, 299, 267, 248, 371, 456, 341, 245, 311, 363, 231, 185, 222, 226, 
    401, 413, 299, 312, 261, 445, 379, 273, 236, 296, 332, 226, 185, 239, 226, 
    453, 442, 318, 309, 294, 234, 260, 253, 255, 272, 240, 158, 119, 214, 287, 
    441, 436, 358, 282, 327, 210, 271, 385, 263, 239, 160, 80, 174, 291, 302, 
    406, 438, 352, 398, 547, 380, 381, 399, 292, 164, 134, 165, 198, 253, 245, 
    272, 386, 413, 560, 495, 210, 169, 164, 166, 159, 171, 172, 190, 202, 196, 
    204, 232, 369, 569, 265, 178, 171, 159, 156, 161, 178, 206, 216, 204, 241, 
    198, 175, 270, 439, 211, 187, 186, 164, 159, 177, 182, 190, 179, 214, 229, 
    209, 166, 178, 200, 149, 143, 170, 178, 194, 211, 191, 169, 238, 289, 186, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 20, 136, 181, 156, 94, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 93, 134, 123, 71, 84, 118, 90, 0, 
    182, 106, 0, 0, 0, 0, 49, 94, 128, 100, 75, 75, 119, 114, 0, 
    261, 192, 0, 0, 99, 19, 45, 60, 107, 180, 114, 102, 135, 142, 109, 
    249, 212, 0, 0, 0, 33, 94, 80, 110, 202, 128, 130, 142, 160, 96, 
    249, 239, 76, 0, 0, 148, 126, 105, 75, 76, 105, 122, 165, 106, 0, 
    298, 311, 231, 133, 0, 57, 33, 100, 95, 0, 63, 85, 113, 0, 0, 
    249, 294, 241, 253, 159, 82, 91, 146, 139, 58, 98, 147, 105, 0, 0, 
    311, 240, 221, 318, 260, 270, 336, 313, 269, 207, 338, 412, 437, 334, 303, 
    612, 405, 257, 269, 331, 463, 488, 496, 537, 556, 613, 641, 678, 678, 683, 
    765, 580, 360, 298, 440, 593, 593, 578, 594, 636, 689, 713, 705, 717, 762, 
    811, 712, 571, 422, 525, 614, 607, 600, 624, 670, 725, 750, 749, 827, 793, 
    789, 774, 666, 544, 577, 629, 635, 614, 627, 666, 692, 700, 742, 806, 757, 
    
    -- channel=10
    242, 243, 248, 246, 248, 237, 252, 268, 262, 233, 210, 212, 216, 224, 231, 
    247, 253, 255, 251, 252, 193, 220, 235, 216, 149, 93, 110, 153, 203, 220, 
    201, 230, 254, 259, 264, 221, 183, 150, 129, 84, 53, 60, 73, 142, 190, 
    71, 130, 231, 259, 225, 191, 109, 93, 81, 114, 71, 102, 85, 94, 171, 
    30, 47, 188, 237, 75, 89, 69, 79, 79, 123, 68, 75, 80, 71, 135, 
    45, 34, 171, 241, 120, 118, 60, 74, 52, 116, 57, 77, 84, 71, 73, 
    42, 12, 159, 210, 143, 120, 67, 71, 56, 88, 51, 67, 78, 78, 73, 
    42, 0, 73, 134, 157, 95, 52, 90, 83, 114, 78, 67, 86, 87, 130, 
    14, 9, 30, 73, 125, 114, 97, 85, 86, 115, 130, 92, 104, 122, 188, 
    42, 23, 6, 45, 54, 107, 94, 33, 71, 126, 87, 92, 84, 168, 209, 
    33, 36, 10, 51, 0, 16, 41, 22, 23, 47, 28, 11, 3, 30, 45, 
    0, 12, 16, 37, 8, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 41, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    168, 178, 169, 175, 174, 163, 181, 185, 174, 165, 149, 142, 143, 150, 146, 
    164, 171, 177, 183, 171, 173, 185, 173, 161, 87, 89, 86, 93, 124, 144, 
    164, 139, 173, 180, 176, 230, 162, 91, 47, 91, 137, 109, 115, 73, 126, 
    134, 43, 172, 177, 178, 112, 136, 95, 89, 104, 168, 117, 96, 60, 83, 
    155, 133, 193, 132, 203, 171, 184, 110, 96, 34, 151, 127, 83, 81, 52, 
    153, 181, 196, 164, 191, 190, 203, 137, 110, 36, 218, 134, 91, 94, 52, 
    131, 229, 146, 181, 142, 139, 249, 162, 145, 108, 198, 108, 76, 79, 100, 
    159, 203, 123, 147, 118, 201, 238, 169, 118, 142, 185, 122, 79, 120, 123, 
    204, 198, 152, 131, 121, 154, 134, 118, 88, 170, 119, 129, 54, 98, 147, 
    212, 201, 192, 107, 152, 96, 100, 172, 113, 150, 132, 40, 51, 141, 175, 
    162, 194, 198, 76, 229, 124, 159, 224, 155, 81, 11, 22, 57, 91, 85, 
    117, 165, 175, 226, 336, 114, 79, 73, 54, 44, 46, 47, 44, 58, 53, 
    56, 88, 104, 305, 162, 51, 57, 49, 42, 33, 36, 42, 71, 62, 44, 
    55, 41, 70, 283, 79, 53, 54, 47, 44, 45, 51, 58, 51, 27, 106, 
    69, 39, 55, 111, 53, 41, 62, 54, 51, 56, 57, 38, 34, 96, 66, 
    
    -- channel=12
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    77, 71, 70, 67, 66, 68, 70, 65, 58, 76, 89, 90, 73, 59, 51, 
    65, 58, 68, 67, 72, 82, 49, 70, 79, 84, 66, 66, 93, 92, 63, 
    83, 140, 70, 62, 71, 137, 75, 61, 65, 142, 114, 109, 70, 96, 95, 
    10, 117, 70, 70, 58, 86, 72, 78, 99, 182, 107, 108, 83, 60, 128, 
    77, 147, 69, 117, 108, 97, 97, 74, 88, 152, 102, 59, 93, 52, 90, 
    136, 208, 80, 80, 250, 163, 111, 76, 41, 213, 141, 89, 120, 84, 50, 
    123, 165, 125, 27, 170, 166, 179, 119, 64, 236, 120, 75, 102, 107, 84, 
    146, 153, 99, 68, 118, 235, 168, 158, 96, 195, 135, 77, 124, 135, 96, 
    170, 210, 93, 167, 88, 164, 99, 91, 136, 87, 127, 99, 110, 107, 79, 
    213, 212, 98, 175, 101, 124, 148, 101, 113, 145, 105, 72, 115, 116, 87, 
    250, 195, 111, 243, 102, 86, 224, 227, 135, 80, 78, 101, 142, 168, 134, 
    290, 272, 164, 284, 209, 172, 170, 164, 146, 146, 160, 166, 168, 173, 164, 
    175, 256, 266, 247, 144, 152, 148, 149, 145, 150, 164, 171, 188, 192, 191, 
    176, 172, 299, 243, 151, 165, 142, 143, 157, 165, 180, 192, 179, 198, 222, 
    171, 176, 182, 193, 150, 178, 188, 166, 161, 160, 155, 169, 191, 183, 147, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 8, 10, 6, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 23, 8, 24, 0, 6, 0, 0, 0, 0, 
    28, 0, 0, 0, 0, 0, 51, 12, 0, 0, 8, 3, 26, 0, 0, 
    84, 0, 0, 0, 21, 0, 5, 20, 0, 0, 42, 0, 29, 14, 0, 
    84, 0, 26, 0, 0, 0, 34, 34, 13, 0, 0, 47, 0, 31, 0, 
    57, 0, 37, 4, 0, 10, 37, 26, 48, 0, 53, 62, 0, 16, 10, 
    52, 8, 0, 53, 0, 0, 6, 31, 57, 0, 68, 35, 0, 0, 11, 
    38, 13, 17, 16, 0, 0, 73, 1, 29, 0, 42, 40, 0, 0, 0, 
    43, 0, 92, 0, 17, 0, 12, 2, 0, 3, 0, 55, 0, 0, 0, 
    2, 0, 98, 0, 35, 0, 0, 4, 0, 14, 52, 0, 0, 0, 11, 
    0, 0, 82, 0, 94, 20, 0, 12, 72, 31, 0, 0, 0, 0, 15, 
    0, 0, 18, 0, 114, 60, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 133, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 0, 0, 72, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    
    -- channel=15
    205, 218, 219, 220, 213, 218, 218, 217, 211, 187, 164, 178, 193, 179, 171, 
    215, 220, 224, 221, 235, 365, 195, 196, 131, 207, 192, 135, 135, 183, 185, 
    144, 205, 224, 220, 223, 232, 164, 101, 137, 288, 222, 200, 132, 107, 208, 
    118, 246, 218, 235, 215, 230, 254, 152, 159, 255, 218, 160, 132, 74, 185, 
    236, 358, 197, 307, 454, 281, 229, 157, 110, 256, 283, 153, 180, 115, 71, 
    203, 379, 212, 160, 383, 277, 333, 201, 124, 413, 255, 135, 189, 157, 111, 
    230, 316, 202, 164, 277, 387, 362, 259, 154, 406, 235, 161, 171, 228, 161, 
    292, 355, 178, 226, 249, 434, 211, 209, 179, 328, 261, 146, 188, 193, 177, 
    347, 391, 169, 327, 193, 185, 207, 227, 249, 172, 213, 70, 123, 218, 227, 
    395, 382, 230, 323, 209, 143, 282, 340, 161, 176, 80, 79, 196, 259, 208, 
    452, 369, 222, 529, 444, 280, 356, 312, 184, 117, 149, 189, 193, 217, 188, 
    270, 385, 336, 586, 273, 145, 160, 155, 162, 165, 183, 188, 214, 214, 201, 
    185, 237, 411, 449, 124, 190, 170, 169, 171, 185, 210, 227, 216, 218, 277, 
    192, 186, 302, 332, 189, 201, 186, 168, 180, 197, 196, 204, 197, 263, 186, 
    186, 197, 183, 182, 137, 167, 183, 191, 220, 230, 186, 196, 309, 271, 154, 
    
    -- channel=16
    216, 226, 225, 224, 214, 228, 229, 212, 203, 199, 187, 192, 201, 188, 160, 
    205, 220, 229, 228, 234, 345, 251, 217, 177, 209, 232, 179, 158, 180, 177, 
    180, 194, 221, 219, 221, 282, 223, 136, 152, 317, 339, 278, 202, 131, 195, 
    195, 199, 235, 228, 229, 232, 305, 224, 209, 319, 336, 248, 190, 106, 165, 
    387, 420, 281, 320, 544, 453, 387, 247, 166, 265, 393, 264, 214, 150, 95, 
    438, 507, 324, 248, 490, 479, 468, 299, 179, 391, 464, 261, 237, 215, 149, 
    458, 485, 287, 191, 303, 467, 533, 392, 253, 438, 425, 257, 219, 270, 234, 
    531, 520, 324, 265, 291, 559, 441, 339, 255, 383, 402, 249, 237, 278, 223, 
    594, 591, 377, 389, 306, 315, 299, 281, 293, 267, 276, 169, 150, 230, 250, 
    582, 585, 420, 407, 370, 250, 351, 443, 297, 273, 165, 95, 192, 268, 241, 
    552, 570, 417, 578, 648, 433, 510, 524, 349, 185, 170, 228, 273, 299, 272, 
    425, 555, 524, 742, 621, 328, 291, 286, 269, 253, 276, 293, 321, 336, 326, 
    326, 381, 553, 710, 359, 296, 284, 268, 260, 271, 304, 337, 352, 351, 394, 
    337, 306, 463, 549, 307, 309, 298, 275, 283, 307, 320, 334, 322, 373, 376, 
    348, 318, 320, 301, 236, 260, 292, 296, 324, 344, 316, 304, 406, 442, 305, 
    
    -- channel=17
    186, 201, 194, 205, 197, 191, 201, 204, 203, 194, 170, 158, 167, 169, 165, 
    189, 196, 199, 211, 200, 262, 221, 208, 160, 122, 141, 106, 93, 139, 171, 
    196, 137, 199, 204, 197, 202, 182, 85, 81, 127, 193, 153, 139, 68, 141, 
    195, 67, 195, 203, 222, 146, 208, 144, 121, 107, 221, 132, 119, 77, 63, 
    253, 207, 228, 173, 362, 245, 237, 160, 108, 39, 214, 182, 119, 120, 29, 
    223, 253, 248, 163, 198, 232, 293, 185, 153, 87, 290, 173, 115, 134, 88, 
    219, 279, 169, 218, 127, 219, 324, 234, 194, 126, 260, 157, 96, 126, 147, 
    261, 279, 170, 203, 136, 285, 289, 178, 167, 145, 238, 155, 99, 143, 139, 
    311, 272, 235, 181, 187, 118, 157, 170, 133, 150, 146, 129, 47, 112, 178, 
    297, 269, 283, 119, 231, 126, 137, 263, 150, 186, 134, 42, 80, 170, 207, 
    229, 269, 261, 174, 415, 258, 246, 290, 236, 105, 62, 93, 105, 128, 137, 
    114, 225, 270, 311, 384, 135, 68, 67, 93, 85, 92, 87, 95, 102, 111, 
    113, 85, 172, 393, 217, 99, 96, 83, 82, 82, 89, 108, 125, 115, 125, 
    119, 83, 82, 352, 148, 96, 106, 87, 85, 94, 95, 102, 94, 110, 141, 
    131, 87, 77, 100, 80, 68, 99, 104, 107, 114, 107, 79, 112, 180, 123, 
    
    -- channel=18
    84, 67, 76, 80, 82, 67, 75, 75, 78, 83, 76, 72, 70, 82, 88, 
    85, 64, 78, 77, 79, 65, 76, 60, 55, 68, 89, 88, 82, 82, 88, 
    78, 76, 75, 73, 83, 71, 48, 70, 94, 102, 104, 105, 115, 111, 79, 
    95, 127, 78, 73, 63, 66, 85, 111, 116, 111, 74, 96, 92, 121, 103, 
    80, 129, 81, 75, 57, 75, 57, 86, 109, 96, 79, 95, 111, 118, 125, 
    75, 86, 63, 57, 21, 22, 48, 92, 111, 119, 69, 76, 113, 111, 115, 
    66, 81, 62, 56, 97, 56, 63, 68, 96, 114, 57, 91, 108, 105, 120, 
    50, 56, 107, 68, 114, 88, 65, 76, 87, 113, 64, 88, 109, 107, 101, 
    49, 61, 75, 78, 82, 62, 67, 93, 109, 80, 80, 83, 106, 103, 102, 
    50, 72, 66, 87, 81, 97, 74, 81, 116, 82, 93, 107, 131, 108, 85, 
    63, 56, 63, 99, 69, 120, 105, 61, 86, 100, 126, 134, 133, 103, 90, 
    131, 59, 76, 96, 36, 53, 86, 86, 111, 132, 142, 139, 138, 147, 140, 
    168, 128, 67, 57, 56, 129, 134, 136, 145, 151, 153, 154, 151, 140, 147, 
    157, 145, 125, 53, 118, 141, 137, 139, 138, 143, 151, 148, 144, 158, 153, 
    153, 147, 136, 117, 145, 145, 144, 139, 143, 143, 151, 152, 153, 158, 154, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 35, 21, 70, 51, 3, 0, 0, 
    29, 0, 0, 0, 0, 3, 50, 51, 26, 25, 114, 93, 109, 0, 0, 
    174, 0, 0, 0, 0, 0, 75, 85, 74, 0, 132, 76, 108, 67, 0, 
    184, 20, 0, 0, 95, 87, 148, 115, 103, 0, 98, 128, 71, 110, 0, 
    148, 67, 19, 0, 30, 82, 142, 116, 150, 0, 154, 138, 58, 101, 79, 
    130, 165, 0, 58, 0, 0, 133, 113, 166, 0, 168, 118, 61, 55, 80, 
    130, 179, 64, 54, 0, 26, 181, 91, 100, 0, 123, 131, 49, 61, 23, 
    170, 128, 178, 40, 50, 68, 85, 87, 14, 82, 42, 136, 36, 0, 0, 
    126, 115, 223, 47, 135, 51, 26, 144, 72, 76, 139, 79, 11, 0, 0, 
    59, 112, 218, 0, 223, 130, 75, 169, 182, 137, 93, 99, 101, 76, 96, 
    85, 90, 136, 14, 295, 186, 143, 143, 148, 139, 143, 153, 158, 159, 174, 
    183, 72, 0, 178, 268, 155, 165, 151, 151, 147, 153, 157, 172, 172, 159, 
    209, 159, 0, 269, 167, 148, 169, 157, 155, 161, 171, 172, 182, 151, 214, 
    222, 180, 144, 173, 153, 130, 147, 153, 150, 167, 184, 156, 127, 224, 234, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 66, 0, 0, 0, 8, 0, 
    0, 73, 0, 0, 0, 0, 0, 0, 5, 89, 0, 0, 0, 0, 24, 
    0, 44, 0, 0, 0, 0, 0, 0, 0, 106, 0, 0, 5, 0, 52, 
    0, 0, 0, 0, 19, 0, 0, 0, 0, 218, 0, 0, 21, 0, 0, 
    0, 0, 0, 0, 54, 23, 0, 0, 0, 182, 0, 0, 21, 24, 0, 
    0, 0, 0, 0, 32, 69, 0, 0, 0, 97, 0, 0, 42, 9, 0, 
    0, 5, 0, 10, 0, 0, 0, 0, 14, 0, 5, 0, 40, 0, 0, 
    0, 3, 0, 88, 0, 17, 16, 0, 17, 0, 0, 13, 53, 0, 0, 
    68, 0, 0, 185, 0, 6, 109, 0, 0, 0, 65, 97, 101, 64, 27, 
    170, 51, 0, 133, 0, 0, 69, 66, 55, 95, 107, 116, 116, 116, 101, 
    114, 172, 98, 0, 0, 90, 90, 94, 96, 114, 126, 131, 116, 119, 130, 
    97, 127, 249, 0, 29, 106, 80, 99, 110, 119, 128, 124, 111, 173, 114, 
    88, 131, 132, 42, 83, 125, 104, 91, 113, 107, 100, 120, 161, 106, 52, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 26, 29, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 9, 16, 17, 14, 16, 6, 11, 
    19, 0, 0, 0, 0, 14, 13, 14, 18, 21, 19, 14, 3, 7, 11, 
    21, 18, 0, 0, 10, 7, 17, 14, 16, 14, 13, 7, 19, 14, 0, 
    19, 21, 7, 0, 15, 9, 5, 14, 13, 13, 14, 17, 9, 0, 28, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 7, 0, 0, 10, 10, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 11, 2, 0, 0, 0, 12, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 12, 14, 7, 0, 0, 5, 0, 0, 5, 0, 
    4, 11, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    9, 12, 5, 0, 5, 0, 0, 0, 0, 7, 6, 0, 0, 0, 0, 
    10, 6, 8, 0, 0, 0, 15, 27, 16, 0, 0, 0, 0, 0, 0, 
    33, 25, 17, 4, 43, 18, 8, 9, 9, 7, 11, 11, 11, 13, 14, 
    20, 23, 9, 21, 14, 8, 12, 9, 8, 7, 9, 8, 20, 20, 8, 
    22, 15, 20, 36, 12, 9, 8, 9, 12, 11, 16, 21, 18, 9, 40, 
    22, 17, 21, 20, 12, 15, 22, 14, 11, 7, 15, 13, 7, 16, 25, 
    
    -- channel=23
    295, 309, 307, 309, 306, 294, 317, 338, 315, 267, 241, 249, 262, 276, 277, 
    304, 320, 315, 318, 306, 279, 273, 285, 234, 143, 93, 106, 156, 230, 269, 
    241, 257, 319, 326, 321, 262, 210, 129, 103, 77, 70, 69, 84, 127, 233, 
    107, 135, 290, 314, 284, 194, 140, 94, 82, 84, 114, 99, 86, 91, 168, 
    49, 87, 250, 215, 160, 119, 111, 97, 86, 71, 88, 94, 83, 82, 111, 
    25, 80, 246, 255, 132, 126, 128, 92, 87, 71, 100, 88, 76, 71, 72, 
    21, 72, 184, 274, 146, 131, 116, 105, 86, 64, 81, 74, 66, 66, 93, 
    39, 43, 63, 176, 136, 116, 106, 98, 111, 119, 107, 76, 66, 103, 170, 
    32, 19, 49, 87, 131, 95, 105, 97, 81, 132, 120, 103, 88, 146, 235, 
    69, 35, 52, 16, 67, 97, 77, 78, 72, 135, 97, 56, 84, 209, 252, 
    35, 47, 48, 18, 45, 18, 37, 41, 42, 25, 0, 0, 0, 0, 0, 
    0, 0, 31, 54, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 64, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    159, 158, 156, 162, 163, 151, 165, 169, 168, 162, 146, 135, 134, 141, 139, 
    158, 151, 157, 169, 155, 159, 187, 167, 152, 105, 117, 118, 115, 120, 138, 
    176, 118, 163, 167, 169, 209, 188, 128, 74, 83, 154, 113, 126, 94, 110, 
    165, 61, 168, 161, 183, 119, 147, 113, 106, 91, 184, 134, 120, 91, 64, 
    176, 129, 194, 101, 168, 164, 199, 140, 118, 39, 166, 151, 96, 93, 72, 
    214, 194, 206, 194, 190, 194, 213, 148, 135, 20, 244, 167, 98, 104, 72, 
    191, 246, 170, 174, 112, 154, 239, 183, 158, 83, 233, 149, 103, 99, 121, 
    217, 208, 160, 160, 100, 169, 251, 178, 141, 123, 207, 165, 90, 131, 123, 
    246, 212, 225, 127, 178, 165, 168, 149, 94, 192, 156, 150, 78, 91, 132, 
    239, 222, 236, 112, 184, 114, 106, 175, 161, 151, 137, 53, 44, 123, 174, 
    175, 223, 243, 75, 240, 151, 145, 215, 172, 109, 56, 48, 87, 134, 145, 
    148, 177, 185, 207, 394, 208, 147, 140, 115, 90, 90, 94, 95, 112, 114, 
    126, 130, 131, 335, 244, 95, 96, 92, 92, 85, 86, 95, 115, 108, 99, 
    124, 96, 109, 306, 136, 96, 106, 92, 84, 90, 108, 114, 108, 94, 163, 
    133, 91, 117, 156, 117, 94, 101, 90, 86, 104, 115, 90, 77, 154, 126, 
    
    -- channel=25
    132, 159, 154, 146, 135, 161, 157, 148, 135, 119, 116, 132, 145, 133, 112, 
    137, 172, 164, 149, 156, 222, 146, 152, 113, 118, 103, 82, 88, 118, 118, 
    97, 127, 146, 150, 139, 131, 90, 55, 86, 158, 112, 100, 61, 60, 137, 
    58, 122, 137, 158, 140, 136, 150, 85, 65, 149, 108, 92, 51, 28, 124, 
    117, 196, 124, 215, 310, 229, 155, 91, 44, 149, 161, 93, 87, 52, 53, 
    93, 180, 139, 114, 225, 211, 194, 117, 48, 241, 133, 63, 94, 73, 70, 
    123, 142, 125, 118, 173, 223, 201, 136, 79, 220, 109, 73, 73, 108, 77, 
    168, 182, 101, 127, 152, 264, 99, 101, 84, 171, 118, 56, 97, 100, 91, 
    179, 205, 65, 174, 102, 104, 99, 98, 129, 76, 106, 21, 59, 117, 148, 
    179, 182, 93, 170, 129, 98, 161, 181, 83, 100, 27, 45, 120, 159, 124, 
    207, 189, 86, 285, 222, 166, 208, 165, 94, 40, 47, 79, 65, 50, 30, 
    68, 171, 176, 301, 82, 0, 20, 20, 15, 15, 15, 19, 26, 19, 16, 
    0, 57, 196, 196, 0, 37, 32, 22, 7, 9, 17, 28, 26, 26, 46, 
    0, 11, 131, 76, 12, 32, 21, 25, 31, 28, 4, 1, 0, 27, 0, 
    0, 12, 12, 0, 0, 0, 10, 27, 50, 38, 6, 6, 72, 30, 0, 
    
    -- channel=26
    14, 15, 18, 7, 9, 20, 17, 12, 10, 13, 12, 26, 15, 4, 0, 
    17, 21, 26, 6, 25, 28, 0, 13, 4, 32, 0, 0, 34, 35, 1, 
    0, 71, 14, 8, 23, 66, 0, 0, 16, 86, 0, 0, 0, 41, 42, 
    0, 117, 9, 30, 0, 35, 0, 0, 0, 131, 0, 4, 0, 0, 119, 
    0, 71, 0, 121, 0, 0, 0, 0, 0, 143, 0, 0, 0, 0, 57, 
    0, 30, 0, 16, 146, 0, 0, 0, 0, 258, 0, 0, 28, 0, 0, 
    0, 0, 6, 0, 146, 76, 0, 0, 0, 231, 0, 0, 10, 24, 0, 
    0, 0, 0, 0, 91, 132, 0, 0, 0, 147, 0, 0, 45, 9, 0, 
    0, 18, 0, 63, 0, 39, 0, 0, 47, 0, 49, 0, 34, 36, 28, 
    0, 9, 0, 113, 0, 0, 54, 0, 0, 0, 0, 7, 73, 72, 1, 
    114, 1, 0, 214, 0, 0, 82, 0, 0, 0, 4, 15, 30, 40, 0, 
    135, 58, 0, 179, 0, 0, 17, 10, 0, 0, 0, 2, 0, 0, 0, 
    0, 113, 110, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 200, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 
    0, 0, 11, 7, 0, 18, 1, 0, 1, 0, 0, 0, 39, 0, 0, 
    
    -- channel=27
    324, 349, 346, 348, 336, 339, 358, 365, 338, 295, 265, 276, 300, 298, 281, 
    329, 363, 359, 358, 355, 419, 341, 324, 256, 200, 175, 141, 163, 251, 287, 
    243, 290, 354, 359, 348, 328, 244, 133, 124, 216, 201, 176, 134, 111, 267, 
    174, 170, 337, 360, 326, 273, 270, 156, 128, 195, 244, 158, 120, 54, 188, 
    255, 288, 331, 356, 498, 356, 283, 168, 97, 158, 274, 186, 144, 108, 64, 
    206, 307, 351, 257, 320, 339, 357, 220, 129, 236, 304, 167, 148, 141, 97, 
    226, 283, 261, 315, 252, 334, 380, 280, 181, 260, 267, 152, 119, 161, 156, 
    280, 324, 183, 293, 244, 385, 295, 210, 188, 253, 263, 142, 130, 181, 211, 
    324, 325, 181, 255, 217, 194, 200, 184, 196, 218, 172, 114, 82, 197, 290, 
    342, 312, 239, 208, 222, 164, 238, 314, 148, 202, 123, 49, 141, 292, 311, 
    310, 323, 236, 320, 431, 245, 287, 305, 199, 94, 31, 63, 57, 99, 92, 
    74, 273, 312, 446, 307, 46, 17, 12, 8, 6, 3, 2, 10, 7, 6, 
    0, 45, 261, 402, 104, 25, 17, 6, 0, 0, 0, 9, 22, 19, 36, 
    0, 0, 93, 286, 58, 22, 18, 1, 6, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 0, 0, 4, 24, 38, 32, 0, 0, 50, 50, 0, 
    
    -- channel=28
    43, 53, 46, 53, 48, 54, 44, 32, 41, 62, 69, 59, 64, 50, 43, 
    45, 41, 43, 53, 50, 147, 87, 67, 69, 109, 165, 112, 64, 56, 57, 
    79, 44, 40, 43, 30, 65, 110, 74, 86, 164, 216, 201, 170, 54, 69, 
    208, 66, 58, 44, 84, 92, 187, 156, 154, 114, 232, 135, 155, 98, 37, 
    316, 231, 122, 76, 343, 236, 240, 176, 136, 82, 232, 196, 154, 161, 26, 
    259, 280, 153, 15, 170, 211, 294, 205, 192, 104, 284, 197, 147, 178, 139, 
    268, 306, 117, 99, 99, 194, 304, 250, 223, 154, 283, 187, 140, 165, 168, 
    291, 348, 192, 177, 100, 242, 292, 183, 183, 123, 245, 181, 134, 153, 117, 
    351, 331, 267, 215, 147, 132, 167, 177, 165, 144, 104, 149, 79, 106, 81, 
    318, 310, 333, 203, 242, 132, 178, 300, 156, 153, 167, 101, 127, 100, 96, 
    285, 299, 316, 228, 490, 300, 276, 333, 296, 194, 170, 211, 217, 222, 217, 
    235, 310, 334, 323, 392, 243, 196, 198, 231, 230, 251, 256, 279, 277, 285, 
    310, 204, 254, 381, 319, 257, 253, 241, 241, 250, 276, 291, 298, 298, 330, 
    329, 275, 172, 425, 270, 260, 272, 244, 250, 268, 280, 286, 296, 306, 321, 
    335, 290, 248, 250, 224, 217, 251, 266, 273, 294, 284, 269, 309, 376, 334, 
    
    -- channel=29
    175, 188, 182, 181, 169, 194, 181, 160, 153, 168, 165, 171, 174, 146, 121, 
    161, 180, 187, 183, 200, 344, 187, 177, 150, 220, 240, 171, 150, 166, 149, 
    146, 197, 178, 169, 178, 290, 163, 111, 160, 403, 364, 303, 205, 136, 194, 
    164, 247, 191, 190, 181, 237, 321, 232, 236, 407, 328, 263, 191, 94, 204, 
    380, 499, 218, 346, 602, 467, 376, 233, 177, 335, 412, 246, 247, 154, 104, 
    421, 564, 250, 206, 562, 462, 463, 300, 173, 544, 453, 231, 283, 237, 150, 
    431, 518, 247, 137, 388, 508, 576, 393, 246, 598, 400, 245, 248, 315, 238, 
    517, 561, 298, 257, 345, 676, 426, 353, 252, 481, 396, 232, 285, 314, 205, 
    603, 659, 326, 445, 286, 334, 285, 300, 337, 262, 298, 146, 182, 246, 234, 
    627, 642, 392, 502, 362, 256, 395, 492, 298, 283, 164, 119, 257, 293, 210, 
    675, 616, 398, 738, 654, 467, 625, 586, 352, 205, 223, 308, 346, 367, 311, 
    575, 656, 559, 905, 611, 321, 347, 338, 320, 338, 372, 395, 429, 439, 421, 
    421, 506, 645, 780, 326, 380, 369, 352, 347, 370, 416, 451, 463, 465, 520, 
    433, 407, 609, 602, 362, 407, 377, 360, 380, 411, 429, 446, 426, 509, 488, 
    440, 429, 408, 392, 312, 358, 392, 390, 429, 447, 409, 410, 550, 562, 379, 
    
    -- channel=30
    0, 4, 0, 2, 0, 0, 0, 3, 13, 24, 21, 0, 0, 13, 29, 
    0, 0, 0, 13, 0, 0, 78, 31, 89, 0, 36, 19, 0, 0, 10, 
    91, 0, 0, 8, 0, 3, 135, 65, 0, 0, 57, 27, 123, 0, 0, 
    343, 0, 0, 0, 64, 0, 54, 45, 8, 0, 166, 5, 103, 48, 0, 
    265, 0, 99, 0, 43, 0, 174, 115, 81, 0, 43, 166, 0, 126, 0, 
    116, 0, 127, 0, 0, 0, 168, 119, 226, 0, 187, 194, 0, 66, 40, 
    72, 147, 0, 213, 0, 0, 96, 106, 249, 0, 241, 121, 0, 0, 58, 
    38, 140, 20, 121, 0, 0, 262, 32, 118, 0, 130, 162, 0, 0, 12, 
    105, 0, 245, 0, 5, 0, 71, 31, 0, 109, 0, 201, 0, 0, 0, 
    10, 0, 340, 0, 141, 0, 0, 109, 0, 28, 200, 5, 0, 0, 37, 
    0, 0, 325, 0, 291, 46, 0, 79, 218, 120, 0, 0, 0, 0, 19, 
    0, 0, 64, 0, 426, 160, 0, 0, 14, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 81, 387, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 0, 0, 345, 74, 0, 12, 0, 0, 0, 0, 0, 0, 0, 41, 
    74, 0, 0, 49, 16, 0, 0, 0, 0, 0, 7, 0, 0, 36, 146, 
    
    -- channel=31
    28, 22, 24, 22, 24, 19, 29, 30, 21, 22, 24, 26, 23, 28, 29, 
    27, 25, 26, 23, 21, 0, 14, 18, 22, 0, 0, 9, 26, 34, 28, 
    17, 47, 26, 24, 26, 8, 0, 10, 9, 0, 0, 0, 0, 37, 31, 
    0, 30, 29, 21, 5, 0, 0, 0, 0, 0, 0, 0, 0, 18, 51, 
    0, 0, 11, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 42, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 11, 5, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 12, 21, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 19, 27, 19, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    187, 199, 195, 196, 195, 189, 204, 220, 206, 171, 152, 156, 167, 176, 178, 
    186, 211, 204, 203, 197, 144, 193, 187, 168, 85, 40, 63, 95, 133, 165, 
    148, 147, 204, 211, 204, 190, 150, 113, 59, 12, 23, 21, 27, 59, 125, 
    77, 17, 181, 205, 184, 134, 75, 41, 13, 18, 62, 49, 42, 19, 73, 
    36, 0, 165, 151, 75, 86, 88, 55, 31, 10, 54, 56, 24, 22, 44, 
    36, 0, 163, 179, 65, 112, 73, 65, 35, 0, 68, 67, 21, 25, 18, 
    39, 2, 111, 205, 65, 51, 61, 60, 52, 0, 66, 41, 16, 8, 27, 
    31, 24, 30, 115, 71, 21, 88, 56, 57, 28, 55, 51, 11, 33, 88, 
    21, 0, 32, 1, 79, 80, 72, 36, 12, 102, 61, 76, 29, 53, 120, 
    28, 1, 29, 0, 40, 57, 42, 26, 27, 70, 57, 23, 0, 93, 162, 
    0, 23, 42, 0, 0, 0, 0, 12, 7, 15, 0, 0, 0, 0, 0, 
    0, 0, 10, 0, 50, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 12, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=34
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 33, 0, 0, 0, 4, 0, 0, 0, 3, 0, 
    0, 12, 0, 0, 0, 31, 0, 0, 0, 37, 0, 0, 0, 0, 20, 
    0, 35, 0, 0, 1, 0, 8, 0, 0, 31, 0, 0, 0, 0, 33, 
    0, 51, 0, 0, 25, 0, 0, 0, 0, 16, 0, 0, 4, 0, 0, 
    0, 30, 0, 0, 62, 0, 1, 0, 0, 79, 0, 0, 7, 0, 0, 
    0, 41, 0, 0, 65, 17, 22, 0, 0, 96, 0, 0, 0, 7, 0, 
    0, 11, 0, 0, 14, 61, 0, 0, 0, 63, 0, 0, 7, 5, 0, 
    0, 10, 0, 39, 0, 0, 0, 12, 1, 3, 15, 0, 2, 13, 5, 
    0, 1, 0, 43, 0, 0, 0, 28, 0, 0, 0, 0, 30, 36, 0, 
    72, 0, 0, 61, 0, 0, 33, 2, 0, 0, 0, 5, 9, 6, 0, 
    43, 19, 0, 94, 0, 0, 0, 0, 0, 0, 1, 2, 2, 5, 0, 
    0, 28, 0, 46, 0, 0, 0, 0, 0, 1, 5, 3, 5, 0, 1, 
    0, 1, 25, 23, 0, 0, 0, 0, 1, 2, 1, 4, 0, 8, 5, 
    0, 5, 6, 17, 0, 5, 2, 0, 6, 3, 0, 0, 17, 4, 0, 
    
    -- channel=35
    395, 419, 419, 418, 411, 404, 436, 456, 421, 346, 299, 325, 353, 369, 364, 
    409, 449, 436, 429, 423, 445, 378, 382, 275, 206, 136, 152, 210, 304, 356, 
    288, 335, 434, 442, 433, 368, 245, 166, 137, 157, 91, 87, 83, 148, 321, 
    125, 231, 402, 437, 387, 285, 222, 97, 77, 138, 133, 111, 75, 65, 246, 
    48, 197, 330, 348, 330, 212, 166, 112, 75, 134, 166, 104, 113, 75, 123, 
    0, 145, 316, 296, 228, 174, 211, 138, 95, 203, 117, 69, 103, 74, 76, 
    1, 114, 239, 360, 243, 234, 191, 136, 96, 185, 86, 80, 81, 101, 103, 
    41, 118, 72, 267, 205, 232, 91, 111, 119, 218, 116, 77, 85, 121, 203, 
    51, 90, 0, 155, 155, 114, 141, 141, 129, 187, 162, 61, 92, 207, 331, 
    111, 81, 36, 94, 88, 97, 144, 169, 78, 134, 53, 43, 123, 313, 331, 
    126, 104, 41, 179, 100, 60, 75, 52, 0, 13, 0, 0, 0, 0, 0, 
    0, 23, 62, 212, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 39, 133, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=36
    37, 37, 37, 37, 37, 34, 38, 42, 42, 41, 38, 38, 33, 39, 44, 
    37, 38, 37, 37, 34, 1, 32, 42, 35, 14, 2, 19, 30, 35, 42, 
    47, 28, 37, 38, 37, 12, 18, 23, 29, 0, 0, 0, 9, 34, 30, 
    16, 11, 34, 36, 36, 14, 2, 16, 7, 0, 0, 7, 9, 34, 26, 
    0, 0, 20, 12, 0, 0, 0, 9, 17, 0, 0, 5, 9, 22, 40, 
    0, 0, 11, 23, 0, 0, 0, 0, 13, 0, 0, 0, 5, 6, 19, 
    0, 0, 8, 42, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 6, 1, 0, 0, 0, 1, 0, 0, 0, 6, 0, 15, 
    0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 17, 18, 13, 8, 25, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 22, 13, 29, 13, 12, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 67, 40, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 8, 0, 0, 30, 63, 11, 8, 0, 0, 
    93, 61, 0, 0, 108, 26, 81, 16, 6, 0, 62, 12, 5, 0, 0, 
    88, 148, 0, 0, 154, 80, 106, 33, 13, 0, 111, 39, 21, 13, 0, 
    76, 161, 0, 0, 21, 38, 166, 64, 59, 62, 110, 21, 0, 16, 4, 
    103, 183, 3, 0, 0, 147, 138, 69, 38, 33, 82, 32, 16, 34, 0, 
    165, 188, 71, 79, 0, 48, 31, 20, 22, 0, 31, 27, 0, 0, 0, 
    178, 169, 138, 74, 95, 0, 28, 109, 13, 48, 32, 0, 0, 0, 0, 
    183, 151, 143, 102, 175, 76, 135, 213, 127, 17, 11, 33, 61, 75, 54, 
    202, 201, 155, 181, 262, 144, 115, 111, 109, 94, 114, 125, 140, 142, 146, 
    153, 149, 130, 251, 181, 120, 119, 107, 103, 108, 130, 145, 165, 163, 175, 
    181, 138, 134, 307, 120, 124, 118, 111, 119, 134, 147, 168, 156, 170, 212, 
    182, 160, 121, 182, 99, 115, 139, 128, 124, 140, 142, 134, 153, 212, 173, 
    
    -- channel=38
    315, 331, 324, 326, 316, 321, 341, 344, 314, 281, 256, 271, 280, 277, 258, 
    307, 339, 336, 335, 332, 372, 316, 306, 243, 200, 161, 161, 199, 250, 266, 
    252, 297, 334, 336, 335, 412, 243, 168, 118, 236, 223, 180, 129, 148, 264, 
    146, 198, 332, 337, 309, 261, 251, 140, 132, 263, 246, 190, 129, 60, 223, 
    203, 308, 315, 333, 415, 319, 300, 168, 124, 186, 289, 166, 154, 83, 105, 
    231, 372, 331, 270, 454, 355, 345, 218, 120, 281, 324, 175, 180, 132, 72, 
    228, 347, 295, 276, 315, 346, 422, 270, 180, 343, 287, 161, 146, 173, 156, 
    285, 363, 190, 277, 244, 448, 331, 269, 194, 342, 277, 174, 164, 222, 219, 
    343, 391, 182, 285, 218, 279, 242, 207, 213, 261, 255, 144, 129, 215, 277, 
    400, 384, 239, 272, 246, 170, 254, 308, 198, 233, 132, 54, 139, 294, 300, 
    399, 384, 265, 384, 324, 207, 307, 358, 184, 92, 41, 43, 90, 164, 133, 
    258, 355, 315, 530, 418, 151, 144, 135, 74, 58, 59, 69, 74, 86, 74, 
    36, 204, 330, 519, 173, 76, 69, 64, 51, 44, 54, 73, 93, 85, 100, 
    40, 46, 261, 390, 91, 86, 65, 60, 60, 67, 64, 77, 52, 72, 105, 
    54, 45, 67, 180, 48, 62, 79, 72, 80, 88, 63, 55, 108, 126, 20, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=40
    40, 47, 50, 51, 51, 48, 50, 55, 59, 46, 31, 30, 37, 39, 38, 
    51, 55, 55, 54, 53, 83, 60, 57, 23, 12, 12, 3, 1, 17, 37, 
    39, 11, 51, 53, 53, 23, 19, 0, 0, 6, 0, 0, 0, 0, 15, 
    13, 11, 39, 59, 65, 30, 34, 6, 0, 0, 10, 0, 0, 0, 0, 
    12, 27, 41, 54, 92, 66, 20, 5, 0, 0, 19, 12, 0, 0, 0, 
    2, 4, 38, 46, 0, 15, 36, 11, 0, 18, 27, 0, 0, 0, 0, 
    7, 7, 0, 44, 7, 41, 27, 21, 0, 10, 3, 0, 0, 0, 0, 
    26, 7, 12, 29, 17, 32, 11, 0, 0, 5, 4, 0, 0, 0, 0, 
    27, 11, 7, 0, 33, 0, 0, 10, 0, 14, 0, 0, 0, 0, 32, 
    11, 6, 3, 0, 0, 14, 8, 28, 6, 0, 0, 0, 0, 39, 48, 
    0, 17, 0, 25, 69, 42, 30, 1, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 2, 54, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=41
    286, 306, 310, 311, 301, 303, 316, 313, 302, 269, 229, 241, 263, 251, 233, 
    294, 316, 319, 318, 325, 476, 313, 299, 202, 221, 217, 153, 147, 220, 251, 
    226, 243, 315, 313, 314, 307, 219, 97, 128, 299, 264, 214, 154, 93, 246, 
    169, 231, 309, 329, 322, 274, 323, 181, 160, 257, 281, 180, 123, 47, 173, 
    300, 418, 310, 380, 624, 432, 323, 193, 104, 218, 345, 207, 180, 111, 52, 
    274, 438, 329, 259, 405, 372, 439, 245, 143, 407, 376, 166, 184, 164, 102, 
    296, 408, 244, 264, 295, 460, 484, 341, 191, 425, 314, 183, 156, 223, 180, 
    390, 434, 231, 297, 285, 545, 330, 248, 190, 361, 319, 160, 172, 214, 190, 
    463, 477, 244, 349, 274, 193, 219, 255, 247, 230, 216, 76, 79, 207, 296, 
    480, 461, 307, 325, 275, 188, 300, 424, 205, 221, 92, 29, 171, 325, 294, 
    489, 463, 290, 551, 612, 379, 459, 414, 246, 117, 97, 165, 179, 211, 188, 
    231, 424, 408, 718, 422, 100, 96, 90, 97, 108, 123, 127, 147, 154, 143, 
    123, 189, 424, 619, 130, 138, 121, 109, 102, 113, 137, 169, 172, 164, 218, 
    118, 116, 279, 415, 155, 146, 135, 109, 120, 138, 130, 131, 120, 191, 145, 
    133, 118, 121, 103, 65, 84, 117, 136, 173, 179, 127, 114, 245, 249, 87, 
    
    -- channel=42
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    25, 26, 0, 0, 0, 5, 8, 12, 0, 46, 83, 65, 9, 0, 1, 
    0, 0, 0, 2, 0, 0, 0, 39, 150, 0, 0, 0, 67, 46, 0, 
    114, 130, 1, 1, 16, 227, 82, 78, 0, 0, 0, 0, 0, 75, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 97, 0, 64, 23, 1, 67, 
    0, 0, 0, 0, 0, 0, 0, 0, 44, 0, 0, 0, 0, 0, 59, 
    19, 0, 0, 146, 288, 97, 0, 0, 0, 0, 0, 35, 8, 0, 0, 
    0, 0, 80, 5, 104, 0, 28, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 46, 105, 131, 9, 46, 19, 5, 23, 51, 0, 
    0, 0, 0, 0, 0, 214, 29, 0, 0, 2, 164, 153, 85, 0, 0, 
    24, 0, 0, 0, 0, 18, 0, 0, 0, 171, 122, 35, 0, 0, 6, 
    10, 0, 0, 0, 0, 0, 0, 116, 0, 0, 0, 0, 0, 11, 11, 
    241, 85, 0, 0, 266, 232, 162, 154, 45, 0, 0, 0, 0, 0, 0, 
    0, 185, 0, 69, 182, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 189, 179, 11, 0, 0, 0, 0, 0, 0, 25, 0, 0, 105, 
    0, 0, 16, 184, 48, 72, 65, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=44
    99, 107, 105, 110, 109, 105, 110, 119, 115, 93, 84, 78, 91, 106, 99, 
    104, 115, 108, 115, 100, 80, 149, 110, 86, 31, 52, 58, 45, 56, 89, 
    90, 28, 108, 116, 101, 41, 107, 66, 40, 0, 46, 42, 62, 28, 43, 
    123, 0, 102, 107, 115, 58, 61, 65, 25, 0, 85, 37, 45, 51, 0, 
    121, 0, 145, 53, 81, 126, 104, 81, 35, 0, 61, 106, 19, 59, 30, 
    119, 0, 163, 105, 0, 101, 91, 83, 76, 0, 113, 102, 0, 46, 65, 
    139, 29, 81, 132, 0, 16, 37, 90, 83, 0, 110, 78, 17, 2, 62, 
    123, 41, 113, 78, 15, 0, 120, 33, 61, 0, 70, 76, 0, 16, 73, 
    99, 5, 147, 0, 97, 21, 58, 28, 7, 72, 0, 78, 0, 15, 73, 
    24, 15, 118, 0, 82, 77, 21, 38, 73, 34, 62, 15, 0, 35, 102, 
    0, 37, 103, 0, 144, 84, 0, 17, 87, 49, 0, 0, 0, 0, 0, 
    0, 0, 63, 0, 90, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 100, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=45
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=46
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 0, 7, 35, 0, 0, 0, 12, 0, 0, 0, 5, 0, 
    0, 34, 0, 0, 3, 18, 0, 0, 0, 89, 0, 0, 0, 10, 22, 
    0, 121, 0, 6, 0, 18, 0, 0, 0, 113, 0, 0, 0, 0, 89, 
    0, 83, 0, 99, 0, 0, 0, 0, 0, 141, 0, 0, 0, 0, 38, 
    0, 30, 0, 0, 96, 0, 0, 0, 0, 268, 0, 0, 19, 0, 0, 
    0, 0, 0, 0, 121, 75, 0, 0, 0, 228, 0, 0, 7, 22, 0, 
    0, 0, 0, 0, 83, 113, 0, 0, 0, 147, 0, 0, 35, 2, 0, 
    0, 9, 0, 53, 0, 3, 0, 0, 43, 0, 8, 0, 23, 39, 23, 
    0, 11, 0, 108, 0, 0, 52, 0, 0, 0, 0, 0, 68, 59, 0, 
    96, 0, 0, 239, 0, 0, 83, 0, 0, 0, 0, 25, 34, 12, 0, 
    95, 47, 0, 193, 0, 0, 0, 0, 0, 0, 4, 10, 9, 13, 0, 
    0, 91, 115, 0, 0, 0, 0, 0, 0, 8, 19, 17, 4, 6, 25, 
    0, 8, 180, 0, 0, 12, 0, 0, 9, 10, 6, 3, 0, 42, 0, 
    0, 9, 17, 0, 0, 18, 4, 0, 20, 6, 0, 11, 72, 0, 0, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    15, 15, 16, 12, 8, 22, 11, 3, 0, 7, 16, 27, 25, 8, 0, 
    14, 13, 14, 7, 21, 82, 1, 7, 0, 70, 63, 46, 49, 40, 10, 
    0, 61, 13, 7, 7, 42, 11, 29, 54, 138, 81, 89, 30, 48, 52, 
    0, 124, 18, 19, 4, 67, 64, 42, 58, 140, 61, 56, 42, 20, 90, 
    72, 158, 11, 109, 145, 88, 66, 43, 35, 159, 106, 29, 73, 28, 41, 
    85, 179, 26, 0, 195, 115, 100, 64, 16, 237, 74, 39, 90, 58, 43, 
    108, 109, 77, 0, 122, 161, 124, 86, 32, 222, 72, 51, 80, 101, 54, 
    125, 150, 78, 49, 87, 187, 64, 85, 60, 152, 83, 43, 96, 80, 56, 
    143, 190, 43, 155, 42, 94, 76, 70, 130, 34, 79, 15, 70, 91, 42, 
    168, 178, 61, 183, 74, 67, 149, 111, 68, 56, 17, 46, 106, 75, 22, 
    231, 167, 68, 303, 133, 102, 167, 144, 73, 53, 94, 109, 123, 132, 96, 
    214, 224, 154, 269, 64, 102, 128, 127, 119, 118, 133, 141, 155, 152, 142, 
    140, 192, 261, 159, 66, 135, 123, 125, 123, 134, 155, 163, 153, 161, 199, 
    148, 152, 244, 130, 108, 147, 127, 125, 134, 146, 148, 157, 152, 193, 138, 
    136, 158, 142, 144, 102, 135, 138, 139, 148, 155, 132, 154, 211, 167, 119, 
    
    -- channel=49
    255, 266, 273, 278, 275, 255, 279, 294, 278, 223, 182, 195, 228, 244, 248, 
    278, 283, 284, 282, 284, 317, 256, 227, 155, 149, 134, 104, 110, 196, 241, 
    153, 195, 280, 287, 280, 171, 156, 94, 116, 133, 105, 118, 111, 94, 210, 
    140, 173, 264, 284, 244, 198, 187, 118, 99, 89, 126, 84, 88, 83, 151, 
    148, 187, 243, 258, 295, 182, 121, 106, 67, 114, 155, 125, 115, 120, 73, 
    39, 119, 234, 140, 58, 111, 182, 145, 118, 151, 102, 81, 97, 111, 116, 
    74, 89, 149, 239, 126, 171, 140, 137, 118, 112, 98, 97, 88, 118, 126, 
    78, 126, 110, 203, 174, 143, 66, 68, 118, 125, 117, 81, 83, 90, 175, 
    83, 82, 55, 137, 116, 43, 112, 123, 137, 117, 76, 44, 59, 173, 244, 
    94, 83, 95, 83, 96, 76, 128, 180, 63, 84, 54, 64, 128, 221, 226, 
    80, 87, 73, 158, 247, 148, 77, 41, 62, 59, 55, 64, 20, 9, 14, 
    0, 24, 128, 156, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 58, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 13, 0, 0, 2, 11, 
    0, 0, 0, 0, 0, 0, 32, 0, 63, 0, 0, 0, 0, 0, 0, 
    35, 0, 0, 0, 0, 30, 80, 54, 0, 0, 28, 11, 43, 0, 0, 
    132, 0, 0, 0, 0, 0, 0, 28, 0, 0, 73, 24, 62, 28, 0, 
    125, 0, 51, 0, 0, 0, 80, 54, 43, 0, 0, 77, 0, 42, 0, 
    135, 0, 72, 28, 0, 60, 26, 53, 70, 0, 106, 130, 0, 26, 0, 
    110, 19, 14, 86, 0, 0, 26, 41, 114, 0, 141, 61, 0, 0, 24, 
    58, 29, 31, 8, 0, 0, 177, 49, 69, 0, 77, 95, 0, 0, 32, 
    62, 0, 150, 0, 8, 58, 54, 0, 0, 45, 0, 151, 0, 0, 0, 
    13, 0, 158, 0, 80, 5, 0, 0, 17, 52, 127, 16, 0, 0, 11, 
    0, 0, 167, 0, 29, 0, 0, 48, 113, 42, 0, 0, 0, 0, 0, 
    0, 0, 41, 0, 272, 166, 32, 34, 27, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 295, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 0, 152, 61, 0, 2, 0, 0, 0, 0, 0, 3, 0, 49, 
    49, 0, 0, 62, 37, 0, 0, 0, 0, 0, 13, 0, 0, 0, 84, 
    
    -- channel=51
    269, 260, 270, 273, 275, 250, 277, 296, 283, 246, 222, 228, 235, 247, 259, 
    276, 269, 273, 276, 275, 218, 241, 240, 210, 162, 110, 129, 173, 228, 251, 
    208, 259, 282, 284, 288, 230, 200, 169, 140, 93, 71, 89, 95, 161, 218, 
    107, 164, 265, 279, 242, 209, 125, 107, 104, 105, 100, 105, 112, 116, 188, 
    59, 69, 226, 226, 86, 73, 81, 100, 103, 118, 85, 92, 107, 103, 142, 
    45, 60, 212, 204, 95, 94, 80, 99, 93, 91, 71, 103, 104, 97, 97, 
    47, 27, 187, 238, 129, 110, 72, 94, 88, 69, 75, 92, 99, 95, 106, 
    28, 31, 85, 179, 145, 70, 84, 102, 121, 111, 93, 96, 95, 105, 176, 
    10, 12, 48, 85, 130, 112, 121, 103, 112, 138, 128, 124, 120, 155, 207, 
    51, 25, 40, 39, 66, 110, 106, 56, 80, 132, 116, 107, 101, 189, 233, 
    39, 36, 45, 42, 0, 18, 12, 25, 44, 77, 53, 21, 8, 53, 68, 
    0, 19, 38, 14, 0, 31, 9, 11, 4, 3, 0, 0, 0, 0, 0, 
    0, 0, 41, 3, 35, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 17, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 13, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=53
    51, 60, 52, 63, 60, 48, 58, 74, 68, 49, 48, 34, 53, 65, 71, 
    53, 56, 48, 68, 44, 0, 97, 47, 86, 2, 21, 6, 0, 20, 53, 
    44, 3, 53, 75, 41, 0, 145, 79, 0, 0, 16, 36, 54, 0, 1, 
    184, 0, 52, 42, 60, 20, 14, 36, 0, 0, 115, 0, 84, 37, 0, 
    208, 0, 119, 0, 0, 0, 104, 83, 30, 0, 27, 106, 0, 77, 0, 
    121, 0, 165, 0, 0, 90, 108, 84, 102, 0, 109, 164, 0, 45, 42, 
    143, 0, 73, 162, 0, 0, 14, 95, 139, 0, 177, 87, 0, 0, 44, 
    82, 70, 50, 91, 0, 0, 173, 24, 113, 0, 110, 106, 0, 0, 83, 
    82, 0, 177, 0, 12, 18, 87, 0, 0, 38, 0, 153, 0, 0, 0, 
    18, 0, 210, 0, 84, 0, 0, 16, 0, 30, 130, 21, 0, 0, 64, 
    0, 0, 199, 0, 180, 0, 0, 14, 146, 63, 0, 0, 0, 0, 0, 
    0, 0, 84, 0, 176, 146, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 298, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 130, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 35, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 83, 63, 40, 0, 0, 
    36, 0, 0, 0, 0, 0, 0, 12, 40, 0, 31, 0, 32, 0, 0, 
    145, 48, 0, 0, 20, 0, 19, 27, 35, 0, 24, 30, 30, 52, 0, 
    122, 101, 0, 0, 0, 0, 44, 11, 75, 0, 66, 34, 22, 57, 32, 
    109, 159, 0, 0, 0, 0, 61, 35, 73, 24, 80, 53, 29, 47, 20, 
    125, 180, 5, 0, 0, 34, 69, 4, 9, 0, 39, 44, 29, 0, 0, 
    190, 190, 144, 47, 0, 0, 0, 32, 0, 0, 0, 3, 0, 0, 0, 
    131, 153, 197, 100, 90, 0, 0, 122, 21, 0, 34, 31, 8, 0, 0, 
    171, 123, 169, 101, 285, 196, 189, 206, 195, 126, 192, 257, 267, 211, 197, 
    327, 225, 161, 126, 251, 260, 260, 268, 322, 340, 383, 397, 429, 422, 433, 
    506, 293, 139, 215, 287, 368, 369, 353, 363, 393, 435, 455, 451, 455, 497, 
    540, 454, 234, 347, 327, 375, 388, 368, 382, 418, 455, 470, 479, 526, 519, 
    529, 493, 404, 328, 343, 361, 380, 380, 392, 428, 441, 429, 463, 554, 521, 
    
    -- channel=55
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    3, 0, 0, 0, 0, 0, 2, 0, 0, 0, 3, 2, 0, 1, 0, 
    3, 0, 0, 0, 0, 0, 14, 2, 0, 0, 0, 8, 8, 0, 0, 
    10, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 2, 17, 0, 
    0, 12, 4, 0, 0, 0, 0, 9, 5, 0, 3, 2, 0, 23, 0, 
    0, 0, 25, 0, 0, 17, 0, 10, 3, 0, 0, 11, 0, 0, 31, 
    44, 0, 37, 33, 0, 14, 0, 0, 0, 0, 21, 15, 0, 0, 14, 
    48, 0, 27, 0, 0, 0, 0, 10, 0, 0, 6, 9, 0, 0, 12, 
    49, 0, 49, 0, 0, 0, 24, 0, 0, 0, 0, 2, 0, 3, 9, 
    20, 0, 58, 0, 45, 0, 0, 0, 0, 0, 0, 12, 0, 0, 3, 
    0, 0, 7, 0, 5, 44, 0, 0, 43, 4, 4, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 11, 7, 0, 21, 0, 0, 0, 9, 0, 3, 
    0, 0, 0, 0, 4, 22, 0, 0, 2, 0, 0, 0, 0, 0, 1, 
    22, 9, 18, 0, 15, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 
    7, 11, 27, 0, 5, 0, 2, 0, 0, 0, 1, 0, 0, 0, 13, 
    12, 0, 23, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    
    -- channel=57
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=58
    36, 36, 37, 34, 37, 38, 29, 30, 37, 41, 50, 52, 50, 43, 50, 
    37, 34, 36, 31, 40, 26, 16, 32, 59, 78, 63, 57, 60, 57, 47, 
    32, 65, 32, 32, 32, 27, 40, 68, 83, 81, 41, 70, 64, 72, 60, 
    37, 78, 23, 37, 26, 70, 39, 68, 75, 79, 33, 58, 72, 78, 86, 
    41, 33, 11, 81, 10, 28, 16, 50, 68, 111, 30, 42, 74, 78, 86, 
    25, 15, 1, 37, 33, 28, 4, 45, 52, 104, 0, 46, 75, 77, 84, 
    32, 0, 24, 30, 73, 39, 0, 32, 42, 80, 10, 47, 76, 74, 54, 
    12, 15, 39, 29, 82, 23, 7, 42, 50, 60, 29, 41, 82, 53, 60, 
    1, 11, 11, 56, 27, 58, 41, 47, 73, 34, 40, 63, 89, 73, 43, 
    11, 13, 5, 74, 13, 70, 77, 23, 33, 52, 73, 106, 92, 48, 34, 
    34, 8, 5, 72, 0, 25, 47, 20, 42, 82, 98, 102, 91, 70, 68, 
    59, 43, 28, 8, 0, 48, 69, 70, 81, 94, 93, 93, 89, 83, 81, 
    77, 67, 66, 0, 31, 88, 87, 90, 93, 96, 97, 86, 79, 90, 85, 
    82, 89, 72, 0, 77, 89, 83, 87, 97, 92, 89, 84, 93, 88, 60, 
    74, 95, 81, 63, 87, 93, 92, 93, 92, 83, 79, 97, 97, 57, 79, 
    
    -- channel=59
    193, 207, 207, 204, 193, 209, 212, 206, 187, 160, 140, 159, 171, 159, 133, 
    189, 214, 214, 207, 217, 323, 199, 188, 106, 142, 121, 95, 111, 146, 148, 
    127, 180, 211, 206, 208, 240, 133, 64, 77, 228, 178, 141, 57, 68, 164, 
    40, 186, 205, 219, 193, 191, 196, 93, 83, 228, 179, 122, 55, 0, 143, 
    168, 308, 201, 298, 419, 315, 229, 113, 44, 209, 250, 108, 106, 17, 40, 
    220, 354, 230, 185, 395, 327, 303, 156, 36, 364, 270, 100, 127, 80, 35, 
    250, 282, 207, 128, 245, 372, 350, 234, 85, 370, 219, 109, 106, 150, 102, 
    322, 319, 171, 177, 201, 434, 245, 196, 120, 311, 224, 97, 126, 159, 133, 
    365, 394, 158, 265, 190, 188, 165, 157, 191, 154, 172, 31, 68, 157, 200, 
    387, 384, 183, 281, 189, 148, 253, 269, 165, 147, 21, 0, 109, 223, 185, 
    404, 382, 189, 499, 371, 236, 344, 313, 139, 41, 37, 73, 106, 148, 108, 
    241, 373, 309, 591, 302, 99, 107, 101, 66, 59, 70, 83, 101, 106, 92, 
    65, 208, 409, 475, 95, 90, 72, 66, 53, 61, 84, 112, 113, 111, 161, 
    62, 78, 322, 281, 84, 102, 78, 67, 73, 89, 85, 92, 74, 141, 97, 
    72, 77, 93, 94, 26, 61, 76, 85, 111, 120, 75, 79, 185, 161, 21, 
    
    -- channel=60
    392, 402, 402, 403, 393, 387, 416, 414, 383, 354, 324, 339, 346, 332, 311, 
    388, 395, 409, 413, 415, 521, 372, 374, 291, 280, 242, 201, 241, 328, 336, 
    316, 404, 415, 409, 416, 461, 314, 170, 165, 359, 320, 272, 194, 194, 352, 
    169, 319, 409, 415, 385, 339, 346, 213, 224, 370, 350, 254, 191, 107, 295, 
    309, 473, 395, 436, 602, 416, 369, 231, 176, 297, 382, 226, 231, 140, 130, 
    330, 567, 422, 331, 604, 462, 483, 276, 166, 478, 447, 234, 259, 206, 121, 
    329, 503, 384, 314, 409, 526, 578, 397, 230, 531, 391, 225, 220, 275, 234, 
    425, 498, 273, 357, 340, 648, 446, 368, 276, 479, 411, 221, 246, 315, 295, 
    511, 562, 284, 446, 316, 336, 308, 301, 331, 306, 327, 180, 180, 312, 373, 
    594, 561, 355, 399, 327, 245, 369, 440, 266, 332, 188, 79, 237, 404, 379, 
    621, 545, 360, 612, 566, 334, 518, 528, 307, 144, 107, 159, 212, 307, 265, 
    412, 573, 474, 808, 561, 247, 213, 200, 180, 170, 190, 194, 212, 223, 205, 
    194, 343, 553, 738, 242, 195, 176, 172, 162, 168, 191, 218, 242, 235, 273, 
    190, 182, 428, 593, 230, 208, 183, 162, 177, 194, 202, 221, 195, 248, 266, 
    197, 183, 208, 256, 154, 182, 216, 205, 218, 226, 185, 184, 289, 294, 147, 
    
    -- channel=61
    338, 348, 340, 351, 345, 333, 357, 368, 351, 325, 288, 279, 286, 294, 288, 
    333, 346, 350, 365, 349, 366, 355, 339, 285, 199, 180, 168, 192, 260, 292, 
    305, 294, 357, 363, 362, 399, 301, 188, 123, 169, 223, 170, 161, 151, 254, 
    226, 140, 354, 357, 348, 256, 262, 159, 143, 185, 266, 188, 152, 95, 170, 
    264, 252, 357, 298, 395, 278, 298, 181, 137, 94, 273, 202, 142, 117, 83, 
    263, 329, 370, 291, 360, 325, 347, 225, 159, 127, 349, 215, 156, 144, 82, 
    243, 345, 308, 328, 235, 292, 416, 279, 221, 198, 328, 186, 132, 156, 170, 
    290, 331, 212, 303, 216, 368, 354, 260, 218, 236, 307, 203, 135, 200, 213, 
    347, 335, 249, 243, 244, 242, 248, 215, 183, 265, 252, 178, 99, 187, 281, 
    374, 339, 304, 179, 277, 148, 193, 298, 190, 248, 171, 57, 101, 262, 332, 
    317, 342, 312, 211, 376, 228, 251, 337, 231, 107, 38, 35, 77, 181, 190, 
    179, 289, 308, 394, 501, 195, 117, 110, 87, 59, 53, 50, 53, 64, 65, 
    51, 129, 230, 499, 253, 58, 55, 46, 42, 32, 34, 48, 75, 68, 63, 
    53, 32, 130, 427, 127, 58, 59, 45, 38, 42, 46, 63, 45, 40, 110, 
    61, 22, 50, 159, 64, 45, 69, 56, 52, 62, 58, 31, 51, 114, 53, 
    
    -- channel=62
    52, 66, 56, 62, 52, 63, 67, 59, 45, 42, 38, 38, 47, 44, 26, 
    48, 65, 58, 68, 56, 120, 91, 62, 32, 19, 51, 31, 13, 25, 37, 
    48, 22, 61, 62, 52, 89, 63, 4, 0, 57, 117, 75, 50, 0, 36, 
    94, 0, 77, 55, 70, 33, 105, 44, 33, 44, 138, 56, 37, 0, 0, 
    168, 145, 116, 34, 248, 171, 173, 76, 28, 0, 149, 96, 36, 25, 0, 
    162, 200, 152, 36, 156, 173, 216, 108, 67, 12, 211, 94, 39, 45, 10, 
    165, 223, 100, 79, 48, 131, 238, 156, 109, 70, 195, 82, 29, 50, 68, 
    204, 236, 99, 113, 30, 189, 211, 110, 89, 76, 156, 87, 26, 77, 57, 
    251, 236, 163, 113, 91, 81, 99, 78, 60, 93, 64, 47, 0, 37, 60, 
    231, 225, 212, 93, 161, 39, 75, 191, 87, 73, 42, 0, 12, 65, 73, 
    185, 225, 209, 125, 318, 164, 154, 220, 145, 32, 0, 12, 28, 56, 51, 
    101, 190, 215, 256, 324, 104, 59, 55, 47, 28, 42, 47, 64, 72, 74, 
    76, 74, 139, 331, 160, 57, 56, 44, 36, 36, 48, 69, 84, 73, 94, 
    84, 57, 67, 286, 73, 58, 66, 49, 43, 55, 59, 69, 63, 69, 116, 
    100, 60, 57, 88, 30, 24, 47, 57, 62, 80, 73, 49, 79, 148, 90, 
    
    -- channel=63
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end inmem_package;
