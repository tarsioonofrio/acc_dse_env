library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    -898, -1227, -985, -3082, -1917, -140, -404, 325, -529, 623, -473, -667, -119, -615, -262, -735, -597, -555, -770, -135, -1357, -196, 182, -311, 914, -1203, -353, -521, -693, 207, -2759, -624, -388, -400, -1066, -4, -691, -726, 294, -551, -311, 110, -1235, 161, -727, -701, -618, -375, -127, -369, -360, -818, -146, -411, -348, -229, 103, -1965, -148, -301, -772, -736, -558, -257, -682, -1326, 110, -308, -6, -1106, -253, 647, -797, -1722, 673, -171, -127, -1102, -754, -182, -796, -740, -538, -755, -273, -100, -342, -608, -2835, -256, -424, -513, -778, -567, -990, -854, -613, -1185, -43, -378, -2143, -212, -551, -244, -931, 111, 41, -660, -763, 246, 38, -476, -1111, -844, -303, 118, 81, -568, -1116, -377, 362, -202, -274, -585, -1348, -861, 125, -781, -552, -1424, 446, -1400, -538, -845, -476, -41, -664, -231, -812, -610, -726, -956, -906, 371, -320, -344, -398, -247, -597, -504, -841, -645, -269, -882, 71, 806, -515, -1032, -370, 15, -478, -1024, 321, -325, -924, 1077, -328, -1286, -117, -703, -1465, -337, -1156, -1311, -233, -138, -1302, -795, -363, -1443, -629, -465, -1248, -790, -982, 1483, 376, -1141, -1282, -270, -685, -1533, -209, -666, 358, 84, -572, -2147, -145, -1267, -673, -425, -241, -664, -714, -40, -707, -422, -119, -1051, -1835, -310, -521, -1033, -1276, 334, -935, -1285, -1432, 789, -365, 983, -1823, -650, -538, -355, -1540, -114, 607, -506, -655, -1397, -589, -695, -606, -1389, -226, -1566, -1349, 161, -1319, -1602, -667, 451, -1236, 210, -1450, -2008, -1173, -166, -642, -527, 482, -160, -158, 159, -249, -950, -1360, -1570, -252, 747, -421, 13, -254, -578, -866, -45, 1471, -746, 430, -939, -58, -853, -265, -903, -439, -173, -137, -1207, -268, -269, -743, 308, -360, -288, -814, -577, -1078, 384, -981, 67, -1103, -284, 386, -437, -292, -1054, -318, 511, -532, -590, 181, -353, -758, -1088, -1395, -210, -726, -1122, -170, -1608, -561, -353, -1281, -818, -205, 152, -644, -994, -700, -379, -704, -174, 4, 273, -413, -253, -164, -546, -167, -599, 18, -399, -1126, -717, 55, 104, 307, -198, 340, 72, -370, -519, -343, -1141, -593, -739, -1177, -243, -181, 335, 64, -2166, -308, -721, -706, -323, -674, -1127, -707, -233, -488, -493, -416, -146, -86, -227, -1000, -332, -716, -1266, -1228, -57, -392, -292, -487, -307, -137, 814, -518, 206, -1523, -476, -1143, -664, -710, 576, -222, -445, -452, 611, -184, -309, -850, -277, -1331, -1852, -670, -2055, 107, 414, -1017, -2371, 69, -529, -119, -716, -30, 163, -978, -699, -910, -1571, -132, -764, -228, -1475, -143, -880, -685, -1064, -219, -242, -885, -791, 202, 211, -623, -426, 35, -726, -220, -218, -2848, -727, -363, -787, -1180, -508, 186, -1212, -397, -693, -1285, -711, -438, -1132, -404, 1000, 155, -1103, 475, -372, 64, -887, -731, -317, -94, -830, -120, -119, -628, 748, 205, -947, -528, -160, -1697, -1787, -247, -887, 630, -345, -465, -1292, -496, 835, 409, -323, -48, -189, -1340, -1078, -1244, -1918, -815, -384, -820, -206, -1499, -545, -282, -161, 352, -104, -424, -954, -683, -412, -672, -18, -1454, -491, -204, -725, 1197, 181, -19, -523, -246, -884, -555, -320, -303, -673, -1741, 404, -1181, -704, -409, -2167, -1779, -660, -816, 77, -404, -552, -287, -312, 17, -915, -15, -444, -214, 180, -108, -903, -1209, 703, 1131, -407, -1431, 128, -477, 107, -672, -215, -74, 281, -1196, -228, -1427, -792, -1595, -1587, -539, -407, 441, -1213, 365, -851, -225, -1287, -406, -677, -674, -699, -897, -64, -90, 625, -599, -355, -494, -763, -487, -1301, -172, -160, 342, -1912, 528, -590, -949, -949, -525, -238, -1216, -646, -298, -373, -1266, 427, -1454, -654, -765, 868, -184, -536, -464, -404, -325, -132, -245, -1130, -454, -418, -511, -559, -407, 135, -623, -669, -100, -742, -319, -730, -229, -152, -154, -429, -364, -799, -167, -71, -67, -335, -85, -718, 2, -1075, -1238, -331, -227, -1673, -522, -625, 342, -860, -31, 29, -285, -188, -1015, -606, -578, 268, -752, -486, -741, -520, -233, -973, -813, -1085, -691, -1639, -1649, -1328, -1190, 972, 47, -961, -501, -584, 191, -466, -888, -535, -200, -779, 264, -889, -1204, -1093, -84, -117, -1133, -982, -872, -387, -364, 438, -1050, 25, 613, -503, -575, 0, -676, -1089, -810, -1524, -1670, 170, -282, -1645, -480, -501, -537, -55, -822, -406, -18, -1851, -502, -1481, -961, -632, -498, -517, -200, -1827, -404, 1440, 222, -526, 289, -285, -1073, -526, -910, 419, -185, -994, -574, -811, -47, -335, -638, -333, -320, 546, 292, -854, -831, -407, 652, 539, -123, -525, -173, 223, -485, -843, -1187, -805, -498, -887, -842, -147, -103, -1012, -1425, -2178, -833, -162, -621, -771, 449, -1120, -1165, -202, -1407, -501, -852, -483, -674, -476, -861, -818, 435, -352, -466, -7, -96, -444, -132, -38, -662, 317, -496, -163, -663, -889, -518, -1520, -1403, 132, -852, -602, 436, -370, -1230, -486, -1531, -740, -1568, -700, 254, 279, 55, -604, -409, -407, -1113, -203, -1093, -1343, -837, -278, -140, -205, 271, -1506, -178, -569, -176, -985, 557, -310, -284, -338, -899, -118, -717, -597, -1026, 284, -686, -306, -907, -1391, -917, -1759, -578, -1133, -970, 193, 507, -402, -1341, -300, -1172, -829, 378, 191, -589, -785, 58, -295, -1107, -1049, -460, -640, 157, -717, -871, -163, -98, -197, -454, -980, -910, -2351, -870, 183, -883, -359, -1305, -196, -817, -329, -145, -415, -1496, -463, -744, -297, -687, -871, -1589, -666, -1110, -929, -15, -196, -1060, 593, -537, -376, -322, 65, -223, -624, -1009, -1174, -1062, -270, -1450, -321, 440, -171, -604, -574, 427, -383, -156, -1192, -1409, -129, -1373, 84, -545, -762, 55, -1596, 25, -364, -511, -360, -2009, -40, -1217, 871, -683, -1130, 283, -599, -715, 1011, -1694, 224, 698, -714, -324, -318, 194, -980, -199, -175, -1069, -427, -328, -1024, 517, -296, -1542, -782, -1000, -1098, 142, -548, -164, -914, -197, -320, -383, 128, -747, -522, -807, -338, -295, -1258, -784, -627, 107, -321, -108, -535, 179, -188, -636, 593, 341, -468, -709, -84, -512, -301, -216, -1507, 118, -557, -562, -479, -395, -187, -471, -276, -323, 4, 40, -1244, -1988, -1093, -563, 325, 9, -1819, 379, 434, -540, -770, -791, 226, -1144, -1513, -332, 177, -623, -691, -836, -917, -1345, -117, -740, -277, -18, -1975, -104, -473, -498, -454, -2181, -1046, 252, -627, -1061, 287, -908, -260, -202, -659, -875, -113, -223, -20, -64, -53, -505, -1303, -423, -781, -695, -1282, -529, -423, -695, -1053, -1564, -866, 234, 102, -1280, -1191, -544, -1603, -227, -595, -2035, -732, -541, -320, -1069, -766, -860, -101, -122, -144, -897, -551, 380, 48, -73, -300, -268, -481, 1519, -508, -215, -865, 149, -317, 108, -359, 553, -693, -1820, -213, -1060, -349, 34, -799, -518, 1, -212, 383, -310, -1092, -76, -796, 299, 22, 142, 46, -353, 85, -1119, -688, 96, -1015, -872, -572, -343, -1341, 254, -560, -676, -122, 74, -378, -27, 563, -781, -385, -928, -216, -818, -403, -540, -239, -526, -407, -943, -401, -1819, 357, -1726, -922, 122, -737, -943, -1427, -1597, -256, -540, -794, -1251, -492, -321, -159, -6, -880, -1045, 27, -37, 191, -1090, -587, -1053, -829, -1463, -311, -1461, -704, -661, -288, -215, -1686, -122, -619, -1551, -75, -401, -156, -1168, 5, 255, -597, -447, -619, -716, -640, -934, -64, 340, -2587, -1428, -312, -521, -40, -623, -597, -831, -740, -817, -764, -636, -186, -1093, -149, 336, -809, -730, -982, -1186, -568, -447, -306, 403, -25, -579, -609, -466, 269, -1659, -1327, -2632, 280, -40, -475, -2427, -535, -521, -510, 462, -53, -534, -743, -766, -367, -554, -147, -1262, 338, -785, -484, 313, -823, -449, 67, -121, -20, -999, -393, -1314, -497, -385, 1, 172, -202, -348, -663, 154, -884, -472, -651, -589, -451, -36, -519, -801, -1205, -287, -681, -1409, -231, -112, 5, -361, 496, -519, -701, -926, -609, -822, 155, -975, -857, 323, -67, -59, -1190, -136, -1839, -715, -838, -1235, -599, -65, -724, -71, -244, -244, -1957, -206, -256, -446, -71, 593, -650, -1054, -728, -1433, -688, -650, -766, -333, -371, -329, 259, -849, -1186, -937, -1765, -990, -1138, -786, -1109, -97, -943, -1839, 275, -766, -1040, 120, -999, -518, -866, 596, -616, -409, -2325, -1681, -667, -504, -972, -1203, 141, -1623, 38, -801, -906, -447, -77, 398, 300, -1751, -965, 60, -250, -514, -335, -297, -589, -995, 89, -680, -406, -1293, 477, -492, -470, -271, -580, 365, -1216, 430, -557, -1690, -990, -3, -767, -851, -232, -575, -84, -237, 217, -325, -748, -792, -901, 82, -241, -689, -118, -362, 206, -647, -781, 76, -1650, -368, -213, -735, 345, 754, -698, -911, -659, -84, -929, -629, -339, -832, -1122, -181, 34, -580, -812, -2952, -437, -2132, 46, -323, -318, -1608, -722, -380, -2552, -645, -1641, -541, -606, -382, 418, -725, -1360, -1354, -451, -86, 12, -189, -618, -61, -334, -135, 183, -460, -1359, -413, -304, -578, -853, -1848, 71, -1204, -134, -555, -338, -1462, -2160, -891, -904, 211, -32, -195, -1341, -74, -397, -1248, -3220, -1243, -908, -479, 276, 292, -742, -26, -580, -996, -352, -1376, -563, -977, -827, 875, -297, 173, -577, 835, -2242, -2, -733, -374, -299, -437, -42, -864, -503, -248, 99, -679, -1875, -373, -659, -1144, -903, -384, 839, -1874, -660, -664, -220, -731, -1553, -1793, -280, -310, -360, -1322, -131, -594, -559, -723, -340, -1015, 578, -1169, -1053, -805, -160, 389, -909, -67, -13, 115, -359, -367, -1332, -185, -424, 525, -69, -343, -1222, -909, -384, -3, -1173, 16, -113, 571, -1418, -652, -150, -1272, -752, -985, -946, -849, -696, -729, -347, -6, -189, -537, -1448, -310, -918, -390, -661, -843, -731, -1627, -611, 267, -255, -1247, -367, -315, -732, -598, -242, -360, -625, -1524, -848, -825, -617, -612, -301, -993, 704, -64, -106, -721, -947, -496, 233, 11, 587, 669, -393, -112, 136, 480, -1461, -1384, -658, -215, -585, -1574, -559, 307, -1160, -118, -746, -693, 95, -328, -697, -364, -1389, -564, -653, -791, -1021, -1562, -734, -504, 461, -789, -165, 64, -15, -1062, 125, -230, -774, -707, -1016, -1070, -1787, -731, -958, -178, -1027, -709, -420, 255, 119, 149, -1577, -99, -754, -541, -984, -646, -187, 399, 738, -262, -2025, -87, 208, -1334, -1469, 264, -3, -666, 117, -403, -716, -1119, -871, -383, -873, 643, -743, -610, -745, -301, 661, -84, -485, -1391, -497, -625, -809, 656, -487, -81, 30, -52, -1539, -1242, -494, -546, -1014, -267, -469, -386, 732, -514, -793, -1749, -217, -1852, -614, -1243, -514, -958, -1122, -593, 442, -430, 163, 66, -1731, -1092, -847, -640, -929, -908, -1244, -307, -1423, -581, -815, -133, 28, -664, -220, -475, 801, -931, -927, -207, -1233, -906, -456, -251, -793, -983, -475, -308, -259, -6, -1183, -510, -588, -1030, -92, 46, -508, -604, 306, -161, -398, -576, 36, 364, -322, 473, -555, -579, -653, -1293, 108, -837, -321, -629, 71, -1618, -1227, -693, -446, -1036, -471, -549, -438, -1259, -329, -652, -1148, -1775, 39, -746, 53, -1232, -282, -111, -1437, -183, -195, 341, -910, -1767, -1438, -227, 161, -146, 263, -874, 3083, -22, -782, -154, -421, -773, -484, -1789, -1315, -677, -680, -905, -543, -39, -1886, -1480, -607, -755, -1221, 206, -606, -153, -2164, -178, 154, -979, 184, -268, 155, -690, -300, -544, -25, 149, -509, -498, -1025, -1215, 156, -1213, 67, -626, -586, 410, 260, -1513, 63, -888, -1218, -1049, -64, -849, -400, -156, -702, -338, 882, -789, -747, -34, -88, -514, -548, -489, -1, -267, -709, -631, -297, -638, 61, -217, -340, -333, -420, -107, -874, -930, -455, 222, -1025, -81, 28, -987, -498, -470, 1033, -1657, -875, -367, -947, -1489, -1062, -367, 162, -246, -1501, -1254, -912, -714, -185, -279, -625, -671, -1378, 204, 321, -1216, -1209, -1171, -989, -293, -10, 199, -395, -10, 116, 1007, -1273, -404, -1856, -840, -666, -279, -154, -769, -973, -506, -200, -952, -724, -766, -1406, -1636, -950, -1411, -1097, -859, -358, 34, -272, 748, -1255, -315, -465, -59, -1410, 96, -1274, -203, -648, 29, -734, -1006, -750, -2428, -910, 523, -213, -1365, -1070, -430, -629, -1789, -162, -495, -781, -104, -706, -1406, 378, -340, -1288, 118, -365, -219, -450, -738, 64, -460, -1796, 106, -598, -1061, 3, -132, -416, -401, -1144, -104, -869, 207, -340, -836, -213, -1223, -90, -1977, -435, 334, 48, -751, -983, -1184, -121, -1021, -77, -702, -1165, -36, -2174, 1189, -346, 189, -1054, -881, -275, -193, 457, -874, -877, -507, -106, -872, -673, -740, -125, -719, 698, -836, -898, 335, -343, -215, -83, -381, -803, 337, -41, -1054, -1333, -379, -1500, -76, 452, -799, -712, -1415, -641, -321, -925, 1164, -184, -612, -1597, -781, -273, -1541, -662, -1665, -1016, -1113, 32, 32, 375, -911, -1233, -419, -248, -1137, -632, -801, -537, 620, -344, -792, -393, 243, -521, -1018, -107, -1052, -590, -385, 317, -1751, -1110, -936, -185, -638, -621, -1608, -1797, -1249, 17, -1071, -1673, -548, -304, -171, -1513, -321, -288, -682, -465, 104, -1078, -1047, 62, -392, 85, -1584, -363, -697, 420, -639, -1028, -115, -303, -1208, -1359, -3, -635, -393, -597, -1143, -597, -713, -790, -1482, -445, -128, -519, -110, -487, -677, -693, -218, -243, 214, -335, -464, -633, -130, -746, -1324, -1103, -150, 189, 54, -704, -86, -204, -37, -19, -127, -1107, -1834, -494, -1575, 256, -835, -886, -1314, -1440, 447, 344, -991, -57, -739, -191, 22, -677, -446, -537, -553, -690, -945, -596, -26, -108, -1756, -997, 348, -554, -1092, 72, -221, -143, -754, -1469, -192, 88, -210, -1339, -2328, -362, -512, -1069, -1078, 356, -1634, -740, -408, -146, -271, -104, -261, -416, -320, -626, -442, -100, -412, -285, -975, -241, -761, -219, -641, -848, -352, -863, -1656, -126, -1103, 576, -618, 889, -675, -351, 45, -403, -1618, -86, -109, -491, -1157, -424, -843, -667, -510, -1502, -393, 608, -454, -550, -77, -542, -346, 92, 315, -321, -1139, -568, 411, -324, -1137, -718, -658, -780, -70, -1343, -1472, -1026, -800, -1605, -1114, -687, -671, -503, -572, 223, -813, -979, 26, -345, 259, 9, -57, -1683, -31, -626, -646, -611, -650, -385, -915, 390, 206, -386, -45, -406, -288, -363, -1731, -13, -1020, -56, 185, -507, -312, -624, -253, -1176, 
    
    
    others => 0);
end gold_package;
