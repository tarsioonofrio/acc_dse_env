LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_signed.all;
	PACKAGE gold_package is
		type padroes is array(0 to 4000000) of integer;
		constant gold: padroes := ( 0, 0, 28, 
		111, 0, 0, 
		86, 61, 0, 
		
		0, 0, 0, 
		162, 37, 252, 
		147, 71, 0, 
		
		0, 0, 0, 
		0, 0, 8, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		182, 86, 0, 
		166, 88, 120, 
		58, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		153, 81, 45, 
		6, 186, 22, 
		129, 176, 213, 
		
		0, 0, 112, 
		76, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		14, 9, 0, 
		0, 0, 0, 
		0, 6, 0, 
		
		124, 18, 0, 
		0, 0, 0, 
		46, 229, 115, 
		
		0, 0, 195, 
		0, 0, 0, 
		12, 116, 154, 
		
		0, 0, 0, 
		52, 157, 82, 
		189, 0, 0, 
		
		0, 230, 255, 
		166, 140, 85, 
		0, 0, 98, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 21, 
		0, 0, 0, 
		0, 0, 0, 
		
		19, 189, 0, 
		15, 251, 66, 
		134, 103, 111, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 226, 69, 
		
		206, 135, 178, 
		86, 112, 10, 
		146, 191, 191, 
		
		0, 0, 0, 
		92, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		242, 129, 24, 
		157, 80, 0, 
		0, 0, 110, 
		
		0, 0, 96, 
		117, 46, 0, 
		233, 130, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		87, 0, 101, 
		0, 60, 12, 
		0, 43, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		196, 93, 0, 
		0, 0, 23, 
		105, 201, 106, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 242, 242, 
		
		0, 0, 66, 
		0, 0, 0, 
		0, 0, 0, 
		
		109, 69, 150, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 2, 
		
		120, 2, 6, 
		0, 0, 0, 
		0, 0, 0, 
		
		32, 134, 233, 
		114, 13, 115, 
		0, 0, 14, 
		
		0, 38, 34, 
		0, 0, 0, 
		195, 227, 223, 
		
		206, 81, 182, 
		29, 244, 191, 
		163, 172, 11, 
		
		0, 150, 0, 
		0, 35, 0, 
		0, 0, 0, 
		
		7, 113, 0, 
		88, 73, 45, 
		0, 0, 0, 
		
		0, 0, 1, 
		0, 104, 0, 
		0, 0, 0, 
		
		199, 71, 230, 
		164, 55, 38, 
		240, 133, 13, 
		
		0, 0, 135, 
		0, 0, 0, 
		0, 94, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		42, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		0, 33, 100, 
		109, 0, 0, 
		0, 0, 0, 
		
		90, 0, 0, 
		0, 0, 34, 
		0, 0, 0, 
		
		0, 0, 249, 
		0, 0, 0, 
		86, 3, 0, 
		
		53, 0, 14, 
		180, 68, 5, 
		235, 91, 0, 
		
		0, 0, 0, 
		20, 0, 0, 
		145, 126, 236, 
		
		87, 0, 0, 
		66, 104, 33, 
		206, 111, 131, 
		
		112, 117, 38, 
		54, 67, 60, 
		24, 237, 201, 
		
		0, 0, 0, 
		0, 0, 0, 
		0, 0, 0, 
		
		153, 141, 36, 
		32, 0, 57, 
		0, 0, 0, 
		
		0, 0, 79, 
		0, 0, 0, 
		0, 0, 217, 
		
		0, 0, 0, 
		0, 30, 0, 
		0, 0, 0, 
		
		253, 61, 0, 
		118, 224, 174, 
		134, 184, 170, 
		
		others=>0 );
END gold_package;
