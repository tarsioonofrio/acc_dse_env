library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package inmem_package is
  type mem is array(0 to 4000000) of integer;

  constant input_mem : mem := (
    -- bias
    -3217, 5289, -47477, 42653, 6831, -20502, -3370, 38122, -63349, 23279, -23287, 110672, -3692, 14946, -3151, 5559, 11161, 48525, 62764, 40712, -68182, -2256, 14330, -18239, -16858, -54280, -37951, 10828, 122620, 25588, -32934, 11479, -86074, -5725, -22567, -2736, 17616, 21823, -9002, 18815, 165760, -10303, 23535, 42713, -8069, 48783, 12392, -31424, -5489, 28243, 67204, 61608, 81473, 30341, -3996, 56384, 12784, -35831, 2234, 41161, -4031, 10214, 75192, -12807,

    -- weights
    -- filter=0 channel=0
    -11, 0, -3, -9, -25, 2, 9, 3, -18,
    -- filter=0 channel=1
    7, -6, -21, -5, 9, 3, -15, 2, -13,
    -- filter=0 channel=2
    -11, 6, -12, -4, 0, -14, 8, -6, 2,
    -- filter=0 channel=3
    -4, -9, -5, -2, -10, -4, -13, -25, -16,
    -- filter=0 channel=4
    -15, 6, 3, 2, -4, 6, -23, 5, -22,
    -- filter=0 channel=5
    5, 1, -19, 1, 6, -8, -27, 4, -2,
    -- filter=0 channel=6
    -27, -25, -24, 4, -3, 17, 1, 5, -11,
    -- filter=0 channel=7
    -11, -19, 5, -6, -1, -17, -17, -9, 10,
    -- filter=0 channel=8
    -17, 0, 7, -15, -8, -7, -17, -1, 0,
    -- filter=0 channel=9
    6, 5, -1, 9, 15, 14, -11, 0, 10,
    -- filter=0 channel=10
    -20, -21, -20, -19, -1, 5, 0, -1, -18,
    -- filter=0 channel=11
    -30, -30, -26, -27, -31, -16, 2, -9, 0,
    -- filter=0 channel=12
    -5, 9, -7, -27, -14, -21, 1, -11, 11,
    -- filter=0 channel=13
    -20, -9, 5, -13, 0, 5, 18, -19, -11,
    -- filter=0 channel=14
    -1, -15, -1, -15, -21, -6, -11, 0, 1,
    -- filter=0 channel=15
    -19, -4, -20, -19, -1, -19, -15, -9, -4,
    -- filter=0 channel=16
    -20, -19, 2, -31, -14, -2, 0, -1, -21,
    -- filter=0 channel=17
    -15, 19, -7, -1, 18, 5, -11, -19, 3,
    -- filter=0 channel=18
    -6, -23, 8, -5, -2, -4, -12, 3, -18,
    -- filter=0 channel=19
    -28, -18, -29, 3, 0, -11, -17, -23, -22,
    -- filter=0 channel=20
    -20, 0, 0, -17, 16, 15, 11, -25, 3,
    -- filter=0 channel=21
    9, -24, -32, -2, -24, -7, 15, -6, 8,
    -- filter=0 channel=22
    -11, 17, -26, 2, 19, 7, -4, 14, -6,
    -- filter=0 channel=23
    -24, -9, -11, -23, 5, 4, -1, -4, -27,
    -- filter=0 channel=24
    7, -14, 5, -2, 0, -9, 2, 0, -22,
    -- filter=0 channel=25
    2, -20, -10, 6, -7, -14, -13, -8, 7,
    -- filter=0 channel=26
    -33, 8, -17, 1, -10, -3, -11, -11, 4,
    -- filter=0 channel=27
    -23, -15, -22, -15, -26, -20, -4, -1, 0,
    -- filter=0 channel=28
    -15, 6, -30, -20, -11, 1, -8, -14, -26,
    -- filter=0 channel=29
    -3, -17, 2, 8, -29, 5, -10, -2, -14,
    -- filter=0 channel=30
    -7, 1, -21, 19, 7, -19, -17, -22, -2,
    -- filter=0 channel=31
    -22, -10, -22, -30, -19, -26, -14, 7, -5,
    -- filter=1 channel=0
    74, 23, -97, -48, 48, -83, -233, 133, 21,
    -- filter=1 channel=1
    -358, -168, -24, -34, 90, -195, 22, 160, -12,
    -- filter=1 channel=2
    40, 149, 33, -97, -13, 128, 99, 27, -77,
    -- filter=1 channel=3
    71, 71, 60, 66, 59, 66, -42, 71, 69,
    -- filter=1 channel=4
    -123, -119, 32, -48, 2, -66, 45, 322, 132,
    -- filter=1 channel=5
    11, 89, -44, -62, -92, 207, -159, -127, 0,
    -- filter=1 channel=6
    -186, 10, 17, 225, 85, 67, -54, -76, 30,
    -- filter=1 channel=7
    -80, 18, -136, -190, -382, 41, -27, -83, -143,
    -- filter=1 channel=8
    -172, 104, 65, -262, -150, 99, -32, -95, -242,
    -- filter=1 channel=9
    -44, -98, -112, -244, 36, -266, -47, 35, -78,
    -- filter=1 channel=10
    184, -97, -10, -92, -130, -135, -36, 121, -128,
    -- filter=1 channel=11
    -88, 111, -117, -109, -53, -26, 152, 143, 54,
    -- filter=1 channel=12
    80, 125, -86, -174, 194, -106, -9, -106, -107,
    -- filter=1 channel=13
    -1, -3, 2, -7, -17, -1, -12, -1, 15,
    -- filter=1 channel=14
    -117, 73, 20, 9, -161, 140, -23, 29, -258,
    -- filter=1 channel=15
    35, -28, 21, 103, -131, 110, 102, -69, 127,
    -- filter=1 channel=16
    -19, -11, 35, -88, -50, 58, 124, -203, 2,
    -- filter=1 channel=17
    -52, -59, -3, -4, -1, -246, 89, 77, 88,
    -- filter=1 channel=18
    30, -18, 152, -18, 39, 105, 99, -154, 1,
    -- filter=1 channel=19
    112, 30, -74, 231, -64, -153, 11, 44, 112,
    -- filter=1 channel=20
    -65, 28, -94, 32, 70, -20, 19, 103, 59,
    -- filter=1 channel=21
    162, 107, -172, -68, -167, -25, -181, 128, -82,
    -- filter=1 channel=22
    -400, -222, -265, 230, -47, 293, 57, 86, -150,
    -- filter=1 channel=23
    -9, 10, -352, -50, -201, 180, 27, -219, -98,
    -- filter=1 channel=24
    75, -4, 44, 94, 87, -24, 49, -15, 144,
    -- filter=1 channel=25
    13, 88, 57, 128, 81, -76, 43, -213, -36,
    -- filter=1 channel=26
    -175, 33, -48, -30, 105, -402, -39, -82, 122,
    -- filter=1 channel=27
    120, -188, 21, -5, 113, 91, 89, 2, -110,
    -- filter=1 channel=28
    43, -88, 112, 160, 141, 222, -187, -176, -152,
    -- filter=1 channel=29
    -26, -138, -229, -149, -393, -149, 16, -203, 22,
    -- filter=1 channel=30
    -17, 32, 142, -100, 194, -91, -213, 121, 31,
    -- filter=1 channel=31
    222, 31, 0, -59, -62, 119, -8, -169, -57,
    -- filter=2 channel=0
    -6, 47, -56, 55, 123, 98, -169, 88, 38,
    -- filter=2 channel=1
    91, -12, 171, 81, 264, 106, 46, -169, 132,
    -- filter=2 channel=2
    112, -196, -213, -46, -356, -206, 83, -42, 155,
    -- filter=2 channel=3
    114, -92, 314, 28, -207, -38, 164, -97, -153,
    -- filter=2 channel=4
    -173, 135, 184, 82, 51, -87, -41, 88, 78,
    -- filter=2 channel=5
    -544, 45, -60, 139, 30, -27, -159, 52, -63,
    -- filter=2 channel=6
    92, -6, 38, -98, -62, 65, -65, 15, -187,
    -- filter=2 channel=7
    99, 1, 103, -253, -207, -64, -64, 69, 85,
    -- filter=2 channel=8
    -101, 104, -50, 15, -92, -79, -190, 217, 33,
    -- filter=2 channel=9
    -14, -207, 216, 67, -160, 20, -40, 78, 42,
    -- filter=2 channel=10
    -20, 58, -92, -124, -131, -130, 11, 115, -5,
    -- filter=2 channel=11
    209, -251, 73, -53, -327, -250, 20, -4, -103,
    -- filter=2 channel=12
    -76, -21, 25, 225, 103, 38, -207, 19, 33,
    -- filter=2 channel=13
    25, -1, -10, -13, -19, 12, -12, 8, 7,
    -- filter=2 channel=14
    128, 142, 37, -80, 71, 9, -66, -38, -34,
    -- filter=2 channel=15
    -8, -393, -36, -269, 42, -57, -139, -128, -103,
    -- filter=2 channel=16
    169, 145, 133, 123, -32, -362, 28, -13, 171,
    -- filter=2 channel=17
    39, -859, 130, 38, -173, 228, -213, 306, 146,
    -- filter=2 channel=18
    -133, -124, -192, -160, 257, 204, -48, 204, -31,
    -- filter=2 channel=19
    -58, 168, 27, -31, -55, 86, 163, -31, -247,
    -- filter=2 channel=20
    16, 91, 37, -68, 199, -244, -377, -175, -198,
    -- filter=2 channel=21
    160, -665, -183, -173, -447, -138, -37, 149, 131,
    -- filter=2 channel=22
    -115, -254, -36, -277, -209, 8, -146, 3, 261,
    -- filter=2 channel=23
    99, -230, 16, 61, 94, 158, -223, 140, -103,
    -- filter=2 channel=24
    127, 143, -78, -133, 15, 339, 102, -120, -55,
    -- filter=2 channel=25
    109, -38, -268, -172, 37, -201, -73, -10, -55,
    -- filter=2 channel=26
    63, 116, -372, 105, 67, 46, -312, 244, -26,
    -- filter=2 channel=27
    -312, 70, 59, -40, -240, 17, -67, 229, 137,
    -- filter=2 channel=28
    -187, -267, -9, 102, -288, 101, 142, 188, -179,
    -- filter=2 channel=29
    146, 148, 108, -21, 97, 2, -122, 90, -263,
    -- filter=2 channel=30
    24, 31, -156, 82, -96, 200, -181, 12, -25,
    -- filter=2 channel=31
    95, -295, -116, 20, -36, 23, 187, -100, 58,
    -- filter=3 channel=0
    112, 61, -120, -1, -409, -291, -209, -324, -89,
    -- filter=3 channel=1
    7, 21, 137, 16, 191, 86, 160, 108, 39,
    -- filter=3 channel=2
    -61, 85, 67, 122, -86, -148, 88, 94, -33,
    -- filter=3 channel=3
    79, -78, -30, -37, 102, 24, 46, -118, -49,
    -- filter=3 channel=4
    61, 83, -8, 166, 133, -180, 103, -98, -84,
    -- filter=3 channel=5
    -112, -26, -38, -198, -74, -174, -295, -240, -44,
    -- filter=3 channel=6
    -21, -120, 224, -33, -182, 82, -176, -358, -216,
    -- filter=3 channel=7
    0, -122, -59, -204, -113, -184, -207, -362, -179,
    -- filter=3 channel=8
    4, -43, -41, -32, 75, -92, -62, -164, 103,
    -- filter=3 channel=9
    5, 53, -73, -34, -239, -193, -114, -206, -593,
    -- filter=3 channel=10
    45, -21, -1, -47, -273, -329, -178, -147, 33,
    -- filter=3 channel=11
    4, -17, 33, -1, 60, 170, -16, -90, 135,
    -- filter=3 channel=12
    -60, 28, 140, -6, 183, -16, 210, 163, 69,
    -- filter=3 channel=13
    0, 16, 15, -10, -17, -27, 0, -15, -1,
    -- filter=3 channel=14
    31, -3, -143, 71, -38, -186, 17, -44, 25,
    -- filter=3 channel=15
    -132, -81, 73, 92, -32, 82, 184, 18, -158,
    -- filter=3 channel=16
    86, -3, 97, -234, -164, -45, 23, -15, -217,
    -- filter=3 channel=17
    -92, -156, 48, -36, 209, 248, -113, 283, 52,
    -- filter=3 channel=18
    115, -121, -21, 0, -4, -22, -223, 99, -47,
    -- filter=3 channel=19
    -146, 106, -10, -99, 166, -7, 87, -69, 63,
    -- filter=3 channel=20
    21, 9, -21, 17, 4, -79, 26, 61, -79,
    -- filter=3 channel=21
    57, -18, 152, -44, 13, -16, 50, -118, -61,
    -- filter=3 channel=22
    23, 19, -95, 106, -246, -170, 7, -89, 42,
    -- filter=3 channel=23
    198, -168, -209, 34, 9, 95, -38, 231, 175,
    -- filter=3 channel=24
    123, -13, -101, 29, 120, 33, 45, 68, 59,
    -- filter=3 channel=25
    49, 41, 131, 1, -69, 56, 10, -35, -182,
    -- filter=3 channel=26
    -40, -39, -31, 116, -33, -75, 147, -34, 46,
    -- filter=3 channel=27
    77, 117, -2, 38, 285, 203, 124, 232, 70,
    -- filter=3 channel=28
    52, 17, 106, -58, 21, -72, -87, -65, 124,
    -- filter=3 channel=29
    10, 112, 59, 96, 165, 189, 307, 264, 26,
    -- filter=3 channel=30
    102, -9, 48, 5, -49, -54, -115, -11, -85,
    -- filter=3 channel=31
    -114, -4, 82, -103, 207, -63, 185, -71, -176,
    -- filter=4 channel=0
    -59, 116, 40, -151, 132, -219, 163, 174, 103,
    -- filter=4 channel=1
    67, -174, -53, 3, -146, -122, -127, 74, -67,
    -- filter=4 channel=2
    218, -241, 64, -157, -214, 134, -37, -162, -85,
    -- filter=4 channel=3
    -290, 42, -313, 19, 50, -163, -43, -202, 43,
    -- filter=4 channel=4
    -54, -6, -272, -42, 53, 79, 53, -274, 36,
    -- filter=4 channel=5
    269, -11, -255, -200, 4, 117, -1, -143, -204,
    -- filter=4 channel=6
    -260, -402, -559, -419, -79, -150, -22, 94, -185,
    -- filter=4 channel=7
    -55, 70, 182, -263, -160, -83, 16, -35, 13,
    -- filter=4 channel=8
    -140, 138, -95, -147, 124, 226, 111, -130, -97,
    -- filter=4 channel=9
    32, -92, -336, 23, -22, 92, 143, -3, 85,
    -- filter=4 channel=10
    -90, 13, -61, 169, 100, 61, 27, -7, 19,
    -- filter=4 channel=11
    -124, 40, 0, -179, -201, -17, 181, -129, 128,
    -- filter=4 channel=12
    145, 72, 83, -253, -21, 93, 249, 148, 114,
    -- filter=4 channel=13
    5, -6, 0, -18, 4, 5, -21, 2, -7,
    -- filter=4 channel=14
    39, 223, -59, -2, 14, 55, -100, 54, 94,
    -- filter=4 channel=15
    -161, 87, -40, -148, 23, -69, 83, -15, -181,
    -- filter=4 channel=16
    -78, -204, -262, -22, -43, 148, 50, -87, 26,
    -- filter=4 channel=17
    246, -39, 44, 54, 107, 90, 235, 82, -92,
    -- filter=4 channel=18
    -33, 145, -17, -198, 303, 265, 90, -33, 346,
    -- filter=4 channel=19
    207, -31, -900, -209, 29, -356, 129, 201, -115,
    -- filter=4 channel=20
    108, -39, -95, -199, 218, 123, -90, -177, -58,
    -- filter=4 channel=21
    141, -7, 3, 75, 59, 97, -104, -282, -329,
    -- filter=4 channel=22
    -87, 94, -101, 20, 190, 367, 231, -122, -356,
    -- filter=4 channel=23
    -129, -79, 170, 66, -226, 33, 92, 0, 72,
    -- filter=4 channel=24
    100, 14, -2, -136, -184, 42, 40, -161, 25,
    -- filter=4 channel=25
    -82, -27, -866, 96, 66, -345, 23, 47, -477,
    -- filter=4 channel=26
    157, -262, -263, -196, 45, 17, 440, -505, -28,
    -- filter=4 channel=27
    230, -92, -327, -188, -271, -268, -112, 63, 85,
    -- filter=4 channel=28
    123, 61, 197, -154, 185, -2, 89, -61, 82,
    -- filter=4 channel=29
    -208, -96, 88, 118, 150, 108, 56, -169, -78,
    -- filter=4 channel=30
    93, -51, -221, 84, 67, -215, -195, 18, -175,
    -- filter=4 channel=31
    -35, -124, -335, -103, 145, -258, -67, 8, -161,
    -- filter=5 channel=0
    43, 18, 11, 71, 237, 122, 50, 118, 26,
    -- filter=5 channel=1
    24, 65, -10, 138, 87, -31, 126, 13, 31,
    -- filter=5 channel=2
    38, 54, 139, -50, 93, -263, 134, 16, -26,
    -- filter=5 channel=3
    0, -175, 111, 24, -401, -236, 131, -188, -39,
    -- filter=5 channel=4
    9, -130, -11, 49, 20, 66, -29, 44, 95,
    -- filter=5 channel=5
    31, 25, -43, -23, 140, -63, 133, 12, -4,
    -- filter=5 channel=6
    63, 50, 36, -175, -19, 89, -180, -3, 136,
    -- filter=5 channel=7
    68, 112, -27, -66, -225, -82, 52, -5, 70,
    -- filter=5 channel=8
    -29, 128, -51, 6, 71, -279, -7, -127, 20,
    -- filter=5 channel=9
    52, -122, -46, 106, -161, 6, -26, 14, -26,
    -- filter=5 channel=10
    216, -140, -315, 115, 129, -184, 47, 53, 40,
    -- filter=5 channel=11
    -96, -108, 190, -120, -155, 52, 96, -126, 53,
    -- filter=5 channel=12
    -69, -51, 223, -187, -221, -48, 2, 56, -91,
    -- filter=5 channel=13
    2, -6, 12, 23, 27, -29, -14, 7, -5,
    -- filter=5 channel=14
    -22, -223, -14, -55, 170, 157, 40, 107, 74,
    -- filter=5 channel=15
    -136, -279, 205, -34, -403, -285, 7, -181, -177,
    -- filter=5 channel=16
    220, 44, 58, 154, -81, -21, -112, -345, 18,
    -- filter=5 channel=17
    -75, 10, 130, 86, -103, -251, -83, 10, -232,
    -- filter=5 channel=18
    -38, -25, -105, 68, 3, 80, -1, 107, 200,
    -- filter=5 channel=19
    103, -94, -84, -20, 23, -242, 100, 231, 45,
    -- filter=5 channel=20
    31, 129, -197, 43, -83, -124, 147, -31, -29,
    -- filter=5 channel=21
    81, 79, 23, -112, 66, -9, 204, -4, -182,
    -- filter=5 channel=22
    -226, -99, -27, -42, 61, 49, -192, -302, 120,
    -- filter=5 channel=23
    -112, -151, -17, 107, -38, -3, 35, 170, 206,
    -- filter=5 channel=24
    -140, -104, 21, -144, -213, 19, 227, 77, -110,
    -- filter=5 channel=25
    -49, 3, -10, -7, 68, -41, -120, -66, -51,
    -- filter=5 channel=26
    -35, -32, -43, -83, -21, 217, 38, 75, -49,
    -- filter=5 channel=27
    8, 18, -45, 90, -85, 63, 20, 9, 191,
    -- filter=5 channel=28
    73, 24, 24, -114, 0, 204, 21, -110, 121,
    -- filter=5 channel=29
    -35, -135, 100, 0, 57, 16, -58, -5, 65,
    -- filter=5 channel=30
    158, 33, -136, 46, -72, -254, -54, 10, -15,
    -- filter=5 channel=31
    -114, -91, 86, -47, -17, 16, 15, 43, 212,
    -- filter=6 channel=0
    4, -21, -13, -1, -10, 10, -6, -9, -33,
    -- filter=6 channel=1
    14, -17, -21, -17, -23, 6, 3, -25, -13,
    -- filter=6 channel=2
    7, -21, -12, -25, -30, -9, -11, -14, -13,
    -- filter=6 channel=3
    8, -19, -10, -6, -25, -18, -10, -3, -24,
    -- filter=6 channel=4
    -19, 5, -7, 3, 8, 8, 11, 5, -22,
    -- filter=6 channel=5
    11, -13, 5, 6, 5, -13, -2, 5, 5,
    -- filter=6 channel=6
    -21, 4, 3, -16, -11, 0, -13, 4, -17,
    -- filter=6 channel=7
    -16, 11, 10, -4, -2, -11, 10, -5, 3,
    -- filter=6 channel=8
    -14, -14, -2, 2, -1, -17, 12, -15, -26,
    -- filter=6 channel=9
    -22, -14, 13, 8, -8, -13, -7, -15, 0,
    -- filter=6 channel=10
    -28, -30, -8, -6, 3, 17, -14, -9, 3,
    -- filter=6 channel=11
    -25, -14, -7, -7, -8, -16, -32, -1, -34,
    -- filter=6 channel=12
    -2, -24, -3, -15, -13, -24, -8, 10, 10,
    -- filter=6 channel=13
    -16, -11, 2, -20, -5, 15, -2, 15, -19,
    -- filter=6 channel=14
    -23, 0, 10, 13, -28, -10, -6, -18, -21,
    -- filter=6 channel=15
    5, -24, -16, 1, 4, -7, -6, -24, -2,
    -- filter=6 channel=16
    -26, -18, -22, -21, 1, -6, -4, -20, 7,
    -- filter=6 channel=17
    0, -21, -3, -9, -1, 8, 15, 3, 13,
    -- filter=6 channel=18
    2, -10, -20, 0, -27, -9, 10, -17, 0,
    -- filter=6 channel=19
    -5, -2, 4, -13, -14, -12, 7, 11, 7,
    -- filter=6 channel=20
    1, -1, -23, -25, 13, -6, -9, 9, -25,
    -- filter=6 channel=21
    -17, -16, 8, -22, 7, 0, -5, -8, -14,
    -- filter=6 channel=22
    -11, 5, -22, -13, -9, -21, 8, 10, -6,
    -- filter=6 channel=23
    -16, -7, 9, -21, -22, -16, -11, 10, -20,
    -- filter=6 channel=24
    -4, -29, 3, 7, -7, 5, -16, 0, -4,
    -- filter=6 channel=25
    -10, -15, -2, 7, -9, -18, -2, -3, 8,
    -- filter=6 channel=26
    -6, 2, 4, 12, 2, 2, -22, 10, -31,
    -- filter=6 channel=27
    -24, 7, -23, -26, -26, -10, -27, 0, 5,
    -- filter=6 channel=28
    3, -23, -12, 6, -9, -11, 7, -12, -30,
    -- filter=6 channel=29
    4, -7, -11, -4, 8, -16, 1, 7, -25,
    -- filter=6 channel=30
    -11, -15, -10, -21, 13, -20, -22, 6, -18,
    -- filter=6 channel=31
    -5, -1, -11, -12, -20, -7, -19, -3, -6,
    -- filter=7 channel=0
    -53, -136, -125, -154, -315, -117, -265, -336, -133,
    -- filter=7 channel=1
    -64, -10, -79, 2, 32, -9, 48, 126, 23,
    -- filter=7 channel=2
    -143, 66, -89, -176, 215, 84, 196, -27, 100,
    -- filter=7 channel=3
    -169, -228, 125, -178, 16, 63, 161, -145, 40,
    -- filter=7 channel=4
    -65, -152, -15, 136, 43, 12, 147, 22, 92,
    -- filter=7 channel=5
    18, -67, -132, -13, -130, -113, -36, 4, -64,
    -- filter=7 channel=6
    98, -124, 1, 127, 150, -225, -67, 83, 116,
    -- filter=7 channel=7
    163, -53, 134, 96, 53, 81, 81, -8, -4,
    -- filter=7 channel=8
    95, -52, 8, -58, -60, 102, 92, -97, -154,
    -- filter=7 channel=9
    -121, -271, -110, -179, -388, -292, -131, 108, -137,
    -- filter=7 channel=10
    -109, -32, 49, 18, -104, -143, 34, -142, 57,
    -- filter=7 channel=11
    104, 74, 164, 21, 76, -8, -112, -51, 54,
    -- filter=7 channel=12
    -7, 91, 56, -80, -29, -42, -65, 112, 72,
    -- filter=7 channel=13
    -16, 5, 19, 12, 2, 15, -13, -32, -15,
    -- filter=7 channel=14
    -54, -108, -89, -31, 15, 38, -215, -40, 47,
    -- filter=7 channel=15
    -127, -318, 60, 69, -225, -222, 134, 8, 108,
    -- filter=7 channel=16
    165, 51, -78, 155, 46, 9, 160, 7, -470,
    -- filter=7 channel=17
    -162, -184, 253, 63, 188, -136, -78, 236, 56,
    -- filter=7 channel=18
    -68, -71, -46, -39, 13, 18, -53, -50, 150,
    -- filter=7 channel=19
    32, -242, 24, 120, -23, -16, 56, 25, 139,
    -- filter=7 channel=20
    -33, 61, 172, -77, -32, 5, 89, -120, -211,
    -- filter=7 channel=21
    105, -282, -174, -116, 140, -54, 272, -58, -65,
    -- filter=7 channel=22
    -151, 34, -218, -57, -42, -6, 141, -87, -61,
    -- filter=7 channel=23
    -36, -10, -100, 51, 43, -44, 78, 71, 128,
    -- filter=7 channel=24
    120, -30, -88, 111, -11, -64, 91, -15, 133,
    -- filter=7 channel=25
    -59, 41, -1, -161, 93, -139, -260, 254, -67,
    -- filter=7 channel=26
    -100, -43, 44, -138, 86, 145, 76, -125, 26,
    -- filter=7 channel=27
    136, 62, -11, -25, 77, 138, -134, 142, 266,
    -- filter=7 channel=28
    80, -9, -45, -22, -64, -87, 16, -66, -115,
    -- filter=7 channel=29
    25, 75, -22, 3, 292, 71, 132, 77, 48,
    -- filter=7 channel=30
    -90, -69, -150, 90, -101, -50, 110, 67, -105,
    -- filter=7 channel=31
    203, 30, -38, 49, 20, -9, 24, -127, 18,
    -- filter=8 channel=0
    15, 163, 45, -36, 107, 103, 19, 129, 112,
    -- filter=8 channel=1
    -180, 30, -157, 77, -78, 98, -26, -133, 18,
    -- filter=8 channel=2
    144, 11, -135, 51, 129, 30, -8, -11, -15,
    -- filter=8 channel=3
    15, 182, -107, 24, 285, 37, 12, 109, -58,
    -- filter=8 channel=4
    -10, 80, 21, 6, 80, 111, -111, -30, 116,
    -- filter=8 channel=5
    -4, 175, -45, 109, -46, -152, 39, 56, -105,
    -- filter=8 channel=6
    11, -105, 101, 97, -151, 143, -90, 74, -114,
    -- filter=8 channel=7
    -178, -23, 24, 118, -24, -26, 128, 163, -21,
    -- filter=8 channel=8
    -199, -42, 87, -247, -150, 75, 70, -58, 50,
    -- filter=8 channel=9
    44, 112, 10, -24, 8, 85, 61, 105, 63,
    -- filter=8 channel=10
    6, -118, 16, 123, -60, -139, 9, 209, 73,
    -- filter=8 channel=11
    -199, -23, -201, 5, 72, 136, -122, 5, 143,
    -- filter=8 channel=12
    100, -24, -154, -17, 92, -36, -105, 49, -5,
    -- filter=8 channel=13
    0, 6, -13, 7, -13, -12, -14, -9, 19,
    -- filter=8 channel=14
    21, -28, -11, 101, 35, 13, -73, 102, -35,
    -- filter=8 channel=15
    68, -111, 101, -96, -42, 90, -181, -200, -22,
    -- filter=8 channel=16
    134, 57, 0, -136, 9, -33, -17, 141, 157,
    -- filter=8 channel=17
    -859, -223, 31, 110, -1, 113, -92, 298, -89,
    -- filter=8 channel=18
    -69, 0, 11, -116, -117, 100, 151, -77, -21,
    -- filter=8 channel=19
    -99, 46, 204, -26, -176, 125, -155, 40, -77,
    -- filter=8 channel=20
    101, -32, -23, -44, 47, 15, -66, -29, 142,
    -- filter=8 channel=21
    236, -168, -187, -192, 49, -85, -284, 43, -137,
    -- filter=8 channel=22
    -200, 205, -2, 100, 43, -45, 117, -33, -92,
    -- filter=8 channel=23
    -87, -140, -176, 124, 12, 65, -44, 115, 128,
    -- filter=8 channel=24
    196, -80, 15, 170, 20, -57, 33, 29, 109,
    -- filter=8 channel=25
    -85, 129, -18, 38, 57, -179, -220, -30, -16,
    -- filter=8 channel=26
    75, 22, 69, 95, -18, -110, 134, 11, -214,
    -- filter=8 channel=27
    -44, -12, -89, 34, 37, 31, 163, 206, 215,
    -- filter=8 channel=28
    260, -213, 65, -267, 44, 15, -109, -77, 37,
    -- filter=8 channel=29
    -147, -292, -106, 48, 8, -151, -170, -30, 12,
    -- filter=8 channel=30
    13, 6, 22, -486, -16, -19, -76, -251, 38,
    -- filter=8 channel=31
    -66, -184, -44, -195, -92, 237, -199, 34, 227,
    -- filter=9 channel=0
    165, -17, -30, 112, -12, 17, 136, 59, 41,
    -- filter=9 channel=1
    -142, -86, -23, 99, -55, 96, -160, 100, 129,
    -- filter=9 channel=2
    -126, 102, 184, 90, 60, -96, -228, 123, -82,
    -- filter=9 channel=3
    -87, -136, 17, -403, -48, 27, -62, -68, 176,
    -- filter=9 channel=4
    -120, 89, -26, 78, -57, -10, 41, -86, -220,
    -- filter=9 channel=5
    168, -53, -62, -18, -17, 84, 23, -77, 192,
    -- filter=9 channel=6
    -27, -68, -39, 68, -146, 170, 11, -14, -102,
    -- filter=9 channel=7
    -140, -60, -68, -306, -117, -126, -181, 62, 226,
    -- filter=9 channel=8
    178, 0, -108, 138, 70, 31, -80, 21, -97,
    -- filter=9 channel=9
    126, 106, -280, -113, -3, -55, 42, 26, 76,
    -- filter=9 channel=10
    8, 64, 76, -155, -148, -138, -119, -114, -5,
    -- filter=9 channel=11
    -109, -106, 29, -244, -224, 128, -192, 101, 4,
    -- filter=9 channel=12
    61, 187, -14, 120, -67, -111, -202, -82, -41,
    -- filter=9 channel=13
    4, -7, -17, 1, -7, -15, -15, 9, 0,
    -- filter=9 channel=14
    52, 50, -11, 83, -131, 7, 97, 39, -96,
    -- filter=9 channel=15
    -115, -183, -224, -10, -32, -81, -180, 26, 41,
    -- filter=9 channel=16
    -65, 183, 86, 53, -170, 75, 1, -34, 39,
    -- filter=9 channel=17
    -557, -6, -151, -148, 170, 50, -307, 79, 210,
    -- filter=9 channel=18
    82, 161, 184, 29, 62, -39, -69, -186, 61,
    -- filter=9 channel=19
    -69, -41, -50, -151, 141, 13, -245, -86, -171,
    -- filter=9 channel=20
    -144, -35, 88, 200, 99, -29, -102, 58, -85,
    -- filter=9 channel=21
    -99, -113, 255, 164, -158, 65, -67, 109, 38,
    -- filter=9 channel=22
    58, 149, 153, -152, 14, 16, -270, 76, -193,
    -- filter=9 channel=23
    191, 71, -44, -96, -41, 50, 72, 125, 168,
    -- filter=9 channel=24
    29, -251, -209, -59, -136, 1, 98, -101, 163,
    -- filter=9 channel=25
    22, 115, 17, 112, 160, 5, -181, 91, 149,
    -- filter=9 channel=26
    221, 129, 30, -33, 109, 29, -16, -57, -18,
    -- filter=9 channel=27
    123, -7, -78, 12, -92, 25, 48, 26, 90,
    -- filter=9 channel=28
    -23, -219, -173, -161, 99, 50, 116, -7, -30,
    -- filter=9 channel=29
    110, -23, 73, -114, 103, 153, 62, -192, -60,
    -- filter=9 channel=30
    -160, -57, 129, 169, -185, 5, -80, 327, 8,
    -- filter=9 channel=31
    76, -79, 43, 7, -71, -73, 48, 32, 34,
    -- filter=10 channel=0
    69, -218, -33, 76, -100, -30, 68, 181, -151,
    -- filter=10 channel=1
    -124, -115, 93, -29, -22, 40, -61, -122, -27,
    -- filter=10 channel=2
    56, -73, 97, -253, 137, 320, 200, 121, -673,
    -- filter=10 channel=3
    48, 148, -22, -96, 145, 86, -89, -133, -139,
    -- filter=10 channel=4
    -185, 84, -32, 22, -221, 26, -13, 90, -122,
    -- filter=10 channel=5
    94, 153, 192, -183, 54, 88, -278, -268, -369,
    -- filter=10 channel=6
    85, 46, 92, -19, -56, -230, 145, -120, -147,
    -- filter=10 channel=7
    -107, 176, -315, -180, -31, 132, -118, -28, 57,
    -- filter=10 channel=8
    -127, 131, -58, -64, 43, -69, -151, -228, 41,
    -- filter=10 channel=9
    -300, -7, 25, -17, 101, 9, -59, 190, 107,
    -- filter=10 channel=10
    -41, -106, -211, 159, -1, -167, 4, 27, -34,
    -- filter=10 channel=11
    44, 79, -46, -130, -29, -83, -121, -93, 100,
    -- filter=10 channel=12
    -121, 7, -13, 177, 130, -102, 65, 68, -213,
    -- filter=10 channel=13
    -5, -10, 0, 4, 1, -15, -19, 19, -11,
    -- filter=10 channel=14
    -13, -267, -7, 126, -91, -51, -226, 165, -104,
    -- filter=10 channel=15
    43, -168, 100, -87, -209, 131, 62, 71, -13,
    -- filter=10 channel=16
    45, 64, 34, -53, -93, -242, -234, -181, 189,
    -- filter=10 channel=17
    -121, 112, 260, 338, -89, 66, 61, -5, -278,
    -- filter=10 channel=18
    -42, -8, -260, 386, 57, 219, 181, -481, -326,
    -- filter=10 channel=19
    -117, 17, -16, -83, -90, -74, 207, -334, -174,
    -- filter=10 channel=20
    52, 119, 2, -45, 27, -19, 79, -169, 103,
    -- filter=10 channel=21
    -299, -49, -14, -6, 113, 81, -483, -37, 2,
    -- filter=10 channel=22
    289, 155, 128, 182, 113, 76, 190, -116, 65,
    -- filter=10 channel=23
    45, -108, 293, 77, -309, -60, -97, 192, -335,
    -- filter=10 channel=24
    -166, -32, -110, -90, -226, -286, 194, -396, -75,
    -- filter=10 channel=25
    32, 94, -141, 123, -102, 79, 41, -887, -226,
    -- filter=10 channel=26
    -16, -231, 0, -46, 13, 104, 87, 3, -53,
    -- filter=10 channel=27
    53, 57, 159, -114, 2, -28, 172, -31, 41,
    -- filter=10 channel=28
    -375, -44, 152, 192, 121, 279, 99, -160, 63,
    -- filter=10 channel=29
    209, -94, 36, -29, -8, -73, -144, 74, 43,
    -- filter=10 channel=30
    208, -74, -45, 18, -66, -153, -26, -24, 59,
    -- filter=10 channel=31
    -56, 31, -59, 0, 222, -132, -42, -102, 90,
    -- filter=11 channel=0
    94, -33, 17, 143, 109, 40, 26, -133, 1,
    -- filter=11 channel=1
    1, -4, -67, -64, -13, 30, 254, -201, 113,
    -- filter=11 channel=2
    36, 182, 38, -204, -225, 79, -126, -254, 52,
    -- filter=11 channel=3
    -172, -63, -11, 107, -53, -109, -63, -19, 57,
    -- filter=11 channel=4
    -20, -80, -1, 2, 18, 36, -5, 66, -100,
    -- filter=11 channel=5
    14, 125, -39, -53, 53, 30, -53, -102, 86,
    -- filter=11 channel=6
    -157, -76, -91, -53, -100, -25, 11, -109, -61,
    -- filter=11 channel=7
    -29, -16, -97, 29, 150, 14, -172, 61, -39,
    -- filter=11 channel=8
    111, 32, -3, -15, 49, 57, 19, -2, 25,
    -- filter=11 channel=9
    45, 72, 60, 49, 93, -149, -69, -46, -51,
    -- filter=11 channel=10
    67, 226, 91, 70, 174, -29, -166, -116, 39,
    -- filter=11 channel=11
    212, -166, -13, 68, -7, -91, -14, -31, -117,
    -- filter=11 channel=12
    -58, 75, 22, -55, -88, 21, 8, -8, 82,
    -- filter=11 channel=13
    -6, 11, 0, 9, 18, -14, -13, 12, -9,
    -- filter=11 channel=14
    75, 154, 17, 9, 10, 3, -101, 23, -129,
    -- filter=11 channel=15
    -119, -50, 173, 73, -41, -77, 35, 96, -139,
    -- filter=11 channel=16
    -76, 85, 46, -83, -82, -273, -245, -293, -99,
    -- filter=11 channel=17
    50, -13, 24, -39, 7, 317, 24, -49, 83,
    -- filter=11 channel=18
    -57, 54, -38, -44, 28, -31, 36, 69, 68,
    -- filter=11 channel=19
    -164, 61, -139, -212, -80, -225, -133, -191, 1,
    -- filter=11 channel=20
    -106, -61, -98, -38, -80, 120, 69, 7, -183,
    -- filter=11 channel=21
    52, -135, 99, 37, -124, 55, 78, -83, -57,
    -- filter=11 channel=22
    12, 46, 3, 93, -77, -12, 160, 199, 44,
    -- filter=11 channel=23
    138, -96, 17, 14, 50, 27, 96, 47, -68,
    -- filter=11 channel=24
    -54, -18, -114, 89, 196, -36, -52, 24, 95,
    -- filter=11 channel=25
    34, 33, -31, -124, -94, -21, 163, -183, -11,
    -- filter=11 channel=26
    -83, 142, 23, -25, -205, -83, -82, -76, -41,
    -- filter=11 channel=27
    28, 110, 118, 37, 102, 186, -14, 0, -61,
    -- filter=11 channel=28
    -134, -58, -32, -10, 80, 70, 18, -127, 49,
    -- filter=11 channel=29
    -42, 43, 26, -259, -93, -23, -57, 94, -26,
    -- filter=11 channel=30
    130, -89, -10, 60, 91, 66, 69, -34, -40,
    -- filter=11 channel=31
    -39, -78, -89, -27, -66, 136, 107, 84, -15,
    -- filter=12 channel=0
    131, 38, -86, 64, 70, -40, 11, 112, 148,
    -- filter=12 channel=1
    -200, 65, 166, -136, -2, -11, 18, 60, -73,
    -- filter=12 channel=2
    -150, -103, 77, 104, -112, -106, -41, -105, -96,
    -- filter=12 channel=3
    44, 84, -29, 33, -25, -83, -203, -14, 95,
    -- filter=12 channel=4
    2, 101, 28, 37, -47, 31, 112, 47, 112,
    -- filter=12 channel=5
    25, -58, -24, -62, -2, 170, -14, -121, 122,
    -- filter=12 channel=6
    -266, -26, 30, -100, -257, -135, -69, -102, -224,
    -- filter=12 channel=7
    -53, 101, 45, -87, 194, -14, 98, -21, -8,
    -- filter=12 channel=8
    -27, -65, -95, 78, -55, -201, 10, -40, 121,
    -- filter=12 channel=9
    222, 47, -45, 164, 107, 3, 31, -22, -78,
    -- filter=12 channel=10
    104, 23, -35, -90, -6, -113, 23, -27, -20,
    -- filter=12 channel=11
    -88, -243, 86, 85, -140, -163, -16, 66, 1,
    -- filter=12 channel=12
    -53, -283, -33, -49, 164, 69, 36, 64, 127,
    -- filter=12 channel=13
    3, -8, 3, 26, -3, 16, 6, -21, -6,
    -- filter=12 channel=14
    9, 111, -62, 130, -10, 12, -72, 55, 123,
    -- filter=12 channel=15
    84, -1, -110, 71, -52, 118, 133, -75, 104,
    -- filter=12 channel=16
    -40, 14, -56, 74, -1, 52, 10, 76, -35,
    -- filter=12 channel=17
    -134, -86, 182, -218, -32, 21, 182, -153, 233,
    -- filter=12 channel=18
    39, -126, 69, -47, -30, -48, 70, -20, 166,
    -- filter=12 channel=19
    -55, -3, 60, 28, -43, 103, 28, -21, -175,
    -- filter=12 channel=20
    233, 23, 54, -58, -53, -107, -96, -239, 128,
    -- filter=12 channel=21
    51, -99, 54, -4, 0, 60, 145, -60, 12,
    -- filter=12 channel=22
    -52, 29, -22, 70, -36, 98, 85, 79, -176,
    -- filter=12 channel=23
    159, -87, 4, -100, -19, -17, 66, 63, 265,
    -- filter=12 channel=24
    -4, -157, 143, -193, -41, 51, -155, -124, -60,
    -- filter=12 channel=25
    146, 46, 89, 24, 119, 5, 100, 38, -51,
    -- filter=12 channel=26
    -122, 31, 249, -202, -16, 73, 92, -13, -78,
    -- filter=12 channel=27
    -44, -62, -123, -137, 64, 78, -192, -77, 92,
    -- filter=12 channel=28
    -148, -174, 170, -65, 59, 67, 46, 41, -193,
    -- filter=12 channel=29
    -151, 76, 130, -55, -4, 20, 207, 135, 38,
    -- filter=12 channel=30
    54, -115, -57, -28, 9, 113, -191, 19, -130,
    -- filter=12 channel=31
    52, -181, 104, -30, -14, -101, 135, 135, 24,
    -- filter=13 channel=0
    -50, 19, -31, 200, -9, -83, 0, -13, 42,
    -- filter=13 channel=1
    -75, -425, 4, -70, 62, -7, -147, 306, 132,
    -- filter=13 channel=2
    82, -300, -153, -2, -24, -630, -161, -260, -242,
    -- filter=13 channel=3
    39, -4, 51, -59, -99, 63, 108, 42, 219,
    -- filter=13 channel=4
    -192, -81, 20, 154, 120, -79, 156, -34, -85,
    -- filter=13 channel=5
    80, -49, -48, 182, 237, -22, -72, -36, -64,
    -- filter=13 channel=6
    44, 71, 124, 21, -140, 75, 45, -131, 56,
    -- filter=13 channel=7
    -178, 22, -149, 78, -128, -152, 17, 142, -28,
    -- filter=13 channel=8
    87, 184, 46, -89, -22, 101, 3, -77, 103,
    -- filter=13 channel=9
    116, 39, 39, 112, 35, 29, 50, 48, 8,
    -- filter=13 channel=10
    -94, -24, -147, 47, -8, 43, -76, 78, -196,
    -- filter=13 channel=11
    21, 213, 68, -52, -212, -1, 46, -246, 100,
    -- filter=13 channel=12
    4, -113, -51, -16, 136, 28, -1, -41, -54,
    -- filter=13 channel=13
    -12, -1, 10, 13, -11, 0, -10, -17, 12,
    -- filter=13 channel=14
    -124, -60, -8, 84, 23, -99, 18, 50, -122,
    -- filter=13 channel=15
    238, -53, -66, -260, 76, -73, 99, -78, -225,
    -- filter=13 channel=16
    -48, -291, -214, 16, 95, 52, 122, -144, -198,
    -- filter=13 channel=17
    319, 415, -150, 11, 99, 24, -98, -20, -117,
    -- filter=13 channel=18
    29, 33, 9, -73, -335, -326, 186, 77, 156,
    -- filter=13 channel=19
    165, 174, 142, -17, -275, -81, -143, 323, 4,
    -- filter=13 channel=20
    110, 125, 139, -8, -39, 104, -467, -205, 191,
    -- filter=13 channel=21
    48, 34, -7, -150, 80, -21, -163, 52, -152,
    -- filter=13 channel=22
    -4, 101, -164, -102, -138, 49, 53, 234, 5,
    -- filter=13 channel=23
    34, -197, -34, -86, -39, -282, 38, -228, 21,
    -- filter=13 channel=24
    30, 38, 34, 100, 157, -151, -11, 102, -12,
    -- filter=13 channel=25
    -140, -438, -1, -126, -78, -187, 31, -43, 42,
    -- filter=13 channel=26
    -291, 82, -36, -139, -99, 81, 214, -71, 250,
    -- filter=13 channel=27
    91, 91, 75, 50, 183, 62, 28, -112, 101,
    -- filter=13 channel=28
    17, 175, 27, -193, 48, 20, -169, -111, -4,
    -- filter=13 channel=29
    -88, -14, -99, -241, -195, -182, 38, -185, 54,
    -- filter=13 channel=30
    195, 2, -30, -46, 235, -56, -572, 161, -117,
    -- filter=13 channel=31
    153, -30, 3, 43, 162, -238, -132, -102, 30,
    -- filter=14 channel=0
    -13, -26, 2, -4, -14, 12, -35, 13, -7,
    -- filter=14 channel=1
    -15, -1, -13, -15, -22, -29, -9, 3, 14,
    -- filter=14 channel=2
    -32, -24, -37, -27, -3, -15, -14, -4, -10,
    -- filter=14 channel=3
    -4, -28, -24, -30, -20, -10, 13, -24, -6,
    -- filter=14 channel=4
    -27, -25, -8, -29, -21, -13, 4, -8, 7,
    -- filter=14 channel=5
    2, -11, -2, -34, -22, -13, 5, -17, -24,
    -- filter=14 channel=6
    -3, -19, 18, -33, -2, -2, 5, 0, -11,
    -- filter=14 channel=7
    -13, -15, -7, 4, -1, -10, 17, 4, 3,
    -- filter=14 channel=8
    -3, 1, -3, -10, -4, -1, -26, -33, -1,
    -- filter=14 channel=9
    -11, -16, -24, -21, 3, -28, -18, -10, 22,
    -- filter=14 channel=10
    -20, 8, 10, -14, -15, -8, -20, -30, -24,
    -- filter=14 channel=11
    -4, -11, -17, 3, -12, -15, -13, -33, 6,
    -- filter=14 channel=12
    -39, -6, -13, -12, 3, -21, -20, -38, -4,
    -- filter=14 channel=13
    7, 14, -6, 6, -17, -11, 5, 3, 0,
    -- filter=14 channel=14
    0, -16, 15, 10, -6, 4, 22, -11, -7,
    -- filter=14 channel=15
    -19, -26, -25, -7, 5, -27, 4, -12, 2,
    -- filter=14 channel=16
    -5, -16, 10, -9, -12, 10, -14, -2, -10,
    -- filter=14 channel=17
    17, -13, -11, -8, 17, -15, -21, 4, -13,
    -- filter=14 channel=18
    -22, 8, -18, 1, 10, -5, -2, -9, -21,
    -- filter=14 channel=19
    -22, -3, -27, 12, -1, -6, 20, -11, 1,
    -- filter=14 channel=20
    -30, -17, 0, -15, -6, 3, -1, -28, 0,
    -- filter=14 channel=21
    -2, -3, 0, 0, -16, -21, -22, -14, 0,
    -- filter=14 channel=22
    -18, -5, 10, -11, -24, -13, 0, 19, 11,
    -- filter=14 channel=23
    -9, -22, -16, 6, 2, -14, -7, -5, -27,
    -- filter=14 channel=24
    -11, -16, 11, -2, -24, -9, -2, 11, -6,
    -- filter=14 channel=25
    9, -19, -13, -6, 12, 6, -13, -2, -13,
    -- filter=14 channel=26
    -9, 0, -6, 0, 13, 4, 4, -13, 13,
    -- filter=14 channel=27
    -33, -10, -15, -19, -1, -5, -31, 4, 1,
    -- filter=14 channel=28
    -2, -13, 4, -24, -26, -11, -4, 4, -1,
    -- filter=14 channel=29
    8, -21, 3, -10, -15, 4, -16, 11, -17,
    -- filter=14 channel=30
    -8, 4, 10, 1, -7, -12, -12, 2, 12,
    -- filter=14 channel=31
    -21, -19, 7, -7, -28, -31, -25, 4, -19,
    -- filter=15 channel=0
    96, -73, 31, -82, 33, 66, -39, -127, -13,
    -- filter=15 channel=1
    -82, -80, 214, -127, 51, 13, -102, -100, -165,
    -- filter=15 channel=2
    -144, 163, -37, 37, 188, -107, -14, 19, -59,
    -- filter=15 channel=3
    -4, -111, 50, 130, 25, 21, 72, 5, 133,
    -- filter=15 channel=4
    -51, -185, -2, 39, -52, -139, 113, -30, 49,
    -- filter=15 channel=5
    60, 37, 26, -66, 220, 238, -38, -93, 128,
    -- filter=15 channel=6
    -115, 68, -190, -25, 53, 81, 63, -91, 188,
    -- filter=15 channel=7
    -89, -127, -8, 93, -19, 37, -103, 98, 246,
    -- filter=15 channel=8
    -8, 199, -41, -109, 167, -59, 10, -140, -195,
    -- filter=15 channel=9
    -47, 31, -10, -34, 94, 129, 132, -83, -29,
    -- filter=15 channel=10
    169, -4, 157, 70, 70, 82, 4, 145, 65,
    -- filter=15 channel=11
    69, 62, -101, 25, -84, -18, 3, 42, -224,
    -- filter=15 channel=12
    -33, -64, 87, 20, -35, 56, 101, -1, 48,
    -- filter=15 channel=13
    26, -5, 0, 10, 11, 15, 6, -13, -3,
    -- filter=15 channel=14
    -54, 61, 100, 45, -54, -26, -90, -47, 34,
    -- filter=15 channel=15
    -118, -67, 43, 40, -12, -23, -74, -60, 95,
    -- filter=15 channel=16
    -221, 35, -44, -147, -141, -138, 193, -92, -112,
    -- filter=15 channel=17
    166, 245, -444, 133, -92, -67, 112, -334, 29,
    -- filter=15 channel=18
    10, 135, 51, -51, 32, 134, -226, 103, 21,
    -- filter=15 channel=19
    13, -165, 279, -511, 70, -279, -28, -17, 122,
    -- filter=15 channel=20
    137, -156, -293, -51, -63, -83, 136, -94, -497,
    -- filter=15 channel=21
    33, 118, 3, -90, -25, -252, -49, -19, -62,
    -- filter=15 channel=22
    158, 5, 39, -32, -22, 182, 119, 114, 155,
    -- filter=15 channel=23
    67, -105, 32, -107, 70, 109, 73, -141, -98,
    -- filter=15 channel=24
    -43, -95, -50, 144, 146, 51, 57, 56, 306,
    -- filter=15 channel=25
    -175, -51, -62, -215, 91, -23, -37, 56, -77,
    -- filter=15 channel=26
    -138, 87, 100, -104, -1, -76, -26, -137, -25,
    -- filter=15 channel=27
    60, 32, 35, -15, -72, 38, -12, 73, 124,
    -- filter=15 channel=28
    54, 216, -185, 49, -76, -122, -24, -180, 34,
    -- filter=15 channel=29
    166, -55, 21, -135, -81, 210, -47, -49, -47,
    -- filter=15 channel=30
    167, 43, -82, 50, -38, 40, -99, 63, -74,
    -- filter=15 channel=31
    35, 161, -1, -145, -125, -75, -112, 99, -219,
    -- filter=16 channel=0
    -133, -99, 47, -275, 1, -13, -275, -18, -8,
    -- filter=16 channel=1
    59, 112, -46, -157, 160, 130, -90, -97, 99,
    -- filter=16 channel=2
    239, 50, -124, -6, -42, -19, -9, 48, 115,
    -- filter=16 channel=3
    -99, -142, -101, -44, 72, -51, 45, -11, 75,
    -- filter=16 channel=4
    47, -65, -219, -224, -323, -76, -759, -60, -2,
    -- filter=16 channel=5
    78, 147, 47, 175, 13, 95, -152, 149, -331,
    -- filter=16 channel=6
    42, -77, 54, -62, -4, -42, -74, 36, 101,
    -- filter=16 channel=7
    83, 36, 121, -96, 3, 33, -238, 156, -133,
    -- filter=16 channel=8
    -111, -24, -29, 26, -158, 16, -101, 248, -166,
    -- filter=16 channel=9
    72, -36, -225, -255, -130, -185, -234, -549, 99,
    -- filter=16 channel=10
    100, -20, -103, 10, 148, -150, -75, 106, 47,
    -- filter=16 channel=11
    55, 57, -41, -5, 71, 207, 67, 12, -98,
    -- filter=16 channel=12
    -35, 136, 82, -86, -60, -52, -61, -222, -195,
    -- filter=16 channel=13
    -8, -7, -9, -10, 19, 20, -13, -16, -12,
    -- filter=16 channel=14
    -179, -63, -61, -292, -35, -177, -289, -191, 104,
    -- filter=16 channel=15
    4, 71, -156, -4, -48, -109, 131, 186, -202,
    -- filter=16 channel=16
    -86, -68, 132, -98, -136, 47, 56, -201, -215,
    -- filter=16 channel=17
    48, 274, 143, 169, -111, -282, 316, -90, -14,
    -- filter=16 channel=18
    -69, -54, -31, 78, 81, 107, 254, 32, -7,
    -- filter=16 channel=19
    0, -31, -131, 222, -40, 146, -63, 143, 54,
    -- filter=16 channel=20
    -212, 38, -167, -11, 78, 122, -170, 42, 69,
    -- filter=16 channel=21
    -70, 87, 74, -142, -67, -157, -221, 28, -65,
    -- filter=16 channel=22
    -170, 133, -100, -160, 42, -73, -4, 49, 106,
    -- filter=16 channel=23
    -76, 83, 100, 121, -124, 336, 58, -253, -24,
    -- filter=16 channel=24
    -25, -29, 149, 26, -55, 14, 63, -8, 102,
    -- filter=16 channel=25
    -49, -166, 168, 205, -178, 49, 0, -45, 35,
    -- filter=16 channel=26
    -14, -70, 58, -114, 81, 73, 76, -137, 55,
    -- filter=16 channel=27
    59, 45, -12, 101, -155, -33, 205, -35, 35,
    -- filter=16 channel=28
    -9, 65, -3, -51, -43, -122, 58, -8, 33,
    -- filter=16 channel=29
    -62, 89, 86, 71, -8, 197, 23, -121, 100,
    -- filter=16 channel=30
    -91, 89, -9, 47, -33, -34, 185, 21, -181,
    -- filter=16 channel=31
    126, 29, 68, 116, -143, -28, 114, -12, 48,
    -- filter=17 channel=0
    -255, -107, -47, -179, -47, -242, -119, -11, -20,
    -- filter=17 channel=1
    -51, -68, -125, 239, 20, -114, 75, -69, 108,
    -- filter=17 channel=2
    -11, -5, -211, 104, -166, -52, 12, -118, -139,
    -- filter=17 channel=3
    128, 81, 66, 106, -121, -184, -109, -109, 131,
    -- filter=17 channel=4
    12, 183, 125, 206, 35, -40, 66, -39, -116,
    -- filter=17 channel=5
    -217, -126, 144, -21, -46, 16, 108, 47, -47,
    -- filter=17 channel=6
    75, -6, 46, -25, -357, -181, -18, -27, -56,
    -- filter=17 channel=7
    -83, -176, -217, 28, -99, -159, 85, 17, -139,
    -- filter=17 channel=8
    98, -2, -190, -125, 44, 69, 19, -102, 223,
    -- filter=17 channel=9
    -78, -122, -30, 47, 108, 28, 179, 92, -97,
    -- filter=17 channel=10
    -177, -114, -35, -180, 24, -16, -49, -46, 71,
    -- filter=17 channel=11
    78, -105, -76, 176, -57, -204, 44, -82, 35,
    -- filter=17 channel=12
    29, 82, 3, -123, 52, -39, 130, 39, 22,
    -- filter=17 channel=13
    -12, 15, -5, -15, -11, 13, -7, 6, -7,
    -- filter=17 channel=14
    39, 90, 11, -8, 0, -5, -52, 102, 59,
    -- filter=17 channel=15
    84, 18, -55, -13, 30, 62, 94, -48, -63,
    -- filter=17 channel=16
    31, -108, -14, 20, 28, 69, 48, -62, 64,
    -- filter=17 channel=17
    270, -64, 45, -71, 55, -175, 185, -11, 109,
    -- filter=17 channel=18
    84, -112, -119, 126, -86, 25, 42, -217, 3,
    -- filter=17 channel=19
    46, 115, -6, 35, -191, -128, 163, 128, -128,
    -- filter=17 channel=20
    31, 71, 107, 71, -197, 22, 128, -22, 129,
    -- filter=17 channel=21
    -80, 120, 63, 3, -113, 44, -125, -145, 100,
    -- filter=17 channel=22
    247, 229, -111, 19, -59, 89, 151, 97, -212,
    -- filter=17 channel=23
    -46, -67, 127, 39, -129, -10, -144, -7, 0,
    -- filter=17 channel=24
    121, -206, 77, 131, -75, 166, 8, -234, -43,
    -- filter=17 channel=25
    17, 18, 35, 52, 54, 84, 75, -52, -16,
    -- filter=17 channel=26
    -118, 59, 5, -17, -206, 112, 240, -3, 15,
    -- filter=17 channel=27
    66, -11, -24, 62, -26, 0, 41, 184, -28,
    -- filter=17 channel=28
    -19, -102, 50, -33, -25, 102, 42, 35, -84,
    -- filter=17 channel=29
    159, 94, -76, 40, 138, 3, 253, 174, -97,
    -- filter=17 channel=30
    -191, -132, 141, 35, -178, 7, -23, -7, 7,
    -- filter=17 channel=31
    10, -50, -14, -15, 143, -23, -172, -18, 247,
    -- filter=18 channel=0
    -179, -5, -101, 111, 82, 0, 93, 51, -71,
    -- filter=18 channel=1
    37, 15, 20, 80, 149, 0, 110, 112, -117,
    -- filter=18 channel=2
    37, -32, 186, -94, 57, 93, -82, -296, -323,
    -- filter=18 channel=3
    31, 124, -47, 152, -203, -105, -160, 38, -68,
    -- filter=18 channel=4
    -138, -329, -335, -132, -150, -131, -140, -180, -18,
    -- filter=18 channel=5
    -178, -88, 68, 75, 146, 92, -61, 130, 63,
    -- filter=18 channel=6
    144, -77, -37, 192, 96, -138, 47, 15, -23,
    -- filter=18 channel=7
    55, -181, 63, -26, 23, 16, 85, 70, -69,
    -- filter=18 channel=8
    -38, -10, -135, -93, -6, -169, -68, -226, 81,
    -- filter=18 channel=9
    -118, -95, 16, -87, -136, -188, -116, -52, 122,
    -- filter=18 channel=10
    -163, 193, 102, 237, 85, -62, -141, 12, 65,
    -- filter=18 channel=11
    -24, 54, 86, 63, -81, 117, -64, -57, 168,
    -- filter=18 channel=12
    -106, 49, 51, -210, -136, -243, -95, -174, 245,
    -- filter=18 channel=13
    11, -23, 1, -13, -3, -13, -6, 13, 31,
    -- filter=18 channel=14
    -130, -44, -296, 111, -64, 36, -17, 98, -162,
    -- filter=18 channel=15
    -39, 22, -238, -154, 137, -253, 3, -6, 33,
    -- filter=18 channel=16
    -62, 125, 371, 177, 28, 7, -31, -2, 34,
    -- filter=18 channel=17
    -147, 2, -187, 0, -152, 115, -111, -155, -137,
    -- filter=18 channel=18
    -193, 47, 8, 44, 96, -146, 307, -178, -111,
    -- filter=18 channel=19
    -42, 326, -74, -61, -124, -299, -141, -194, 218,
    -- filter=18 channel=20
    -115, -134, -108, -101, 185, 132, -4, -31, 20,
    -- filter=18 channel=21
    -33, 67, -74, -120, -78, 246, -38, -38, -266,
    -- filter=18 channel=22
    0, -36, 133, 82, -76, -101, -26, 84, -23,
    -- filter=18 channel=23
    -36, 152, -99, -54, 6, -77, 41, -174, 86,
    -- filter=18 channel=24
    175, -320, -183, -2, 109, -249, 150, 26, 66,
    -- filter=18 channel=25
    -59, -230, 173, -24, 12, -210, 0, 27, 45,
    -- filter=18 channel=26
    -99, 40, -20, -77, 62, -145, -10, -174, 31,
    -- filter=18 channel=27
    15, 10, 75, 34, 111, 35, 124, -171, -96,
    -- filter=18 channel=28
    62, -174, 80, 125, 104, -18, 86, -123, -108,
    -- filter=18 channel=29
    68, 28, -18, 155, -44, -107, 78, -160, 35,
    -- filter=18 channel=30
    -190, 15, -14, -62, 142, 42, 104, -48, -26,
    -- filter=18 channel=31
    128, -92, 60, 37, 36, -6, -1, -205, -46,
    -- filter=19 channel=0
    -116, -127, 39, 1, 86, 198, 5, 118, 91,
    -- filter=19 channel=1
    4, -123, 46, 51, -151, -44, -15, -154, -35,
    -- filter=19 channel=2
    136, -99, 62, 9, 266, -118, -100, -28, 0,
    -- filter=19 channel=3
    -114, 138, 91, -127, -76, 32, 6, -111, -29,
    -- filter=19 channel=4
    -45, -102, -132, 85, -12, -173, -66, -296, 111,
    -- filter=19 channel=5
    30, 36, 90, -284, 74, -77, -43, 136, -87,
    -- filter=19 channel=6
    -143, -358, -207, 57, -123, -11, 131, -180, -137,
    -- filter=19 channel=7
    -17, -144, 37, -175, 56, -3, -65, -145, 97,
    -- filter=19 channel=8
    -115, -165, 129, -349, 74, 118, -116, 63, -30,
    -- filter=19 channel=9
    -105, 30, 60, 34, 118, 8, -24, -92, -35,
    -- filter=19 channel=10
    28, -85, 139, -110, 24, 192, -6, 151, 47,
    -- filter=19 channel=11
    73, -94, -71, 204, -122, -11, -122, -26, 102,
    -- filter=19 channel=12
    -169, -58, 63, 1, 187, 215, -218, 55, 61,
    -- filter=19 channel=13
    -1, 0, -3, 19, -5, -1, -14, -5, -19,
    -- filter=19 channel=14
    5, -151, 87, -58, -39, -75, 86, -5, 7,
    -- filter=19 channel=15
    -36, -205, -22, 128, -55, 80, -67, -50, -22,
    -- filter=19 channel=16
    86, 157, 31, -248, 169, 194, -85, 73, 203,
    -- filter=19 channel=17
    124, -18, 47, 236, 65, -195, 65, 123, -84,
    -- filter=19 channel=18
    -187, -105, -55, 154, 19, 169, -83, -44, -68,
    -- filter=19 channel=19
    -94, 31, 28, -16, 58, -3, 53, 22, 9,
    -- filter=19 channel=20
    -120, 52, -205, 52, -81, -89, -66, 79, -39,
    -- filter=19 channel=21
    8, 132, 103, 133, 98, -88, 40, -109, -143,
    -- filter=19 channel=22
    154, -20, 130, 126, 51, 137, 13, 21, -8,
    -- filter=19 channel=23
    -29, 79, -120, 90, -5, 15, -141, -111, 32,
    -- filter=19 channel=24
    48, 185, -8, 46, -81, -48, 49, 24, -165,
    -- filter=19 channel=25
    -70, -195, 31, 100, 38, 6, -63, 71, -22,
    -- filter=19 channel=26
    -39, -32, -161, 66, -82, 126, 117, 26, 28,
    -- filter=19 channel=27
    -310, -164, 26, 83, -219, -205, -96, -28, -156,
    -- filter=19 channel=28
    36, 207, 51, -82, -60, -33, 8, 43, 60,
    -- filter=19 channel=29
    -32, -96, 95, -121, -84, -94, -83, -80, 135,
    -- filter=19 channel=30
    74, 16, 54, 53, 22, 86, 17, 155, -29,
    -- filter=19 channel=31
    -33, -44, 35, -88, 129, 111, 2, 127, -35,
    -- filter=20 channel=0
    62, 116, 45, 85, 102, 138, -91, 86, -50,
    -- filter=20 channel=1
    131, 28, -14, 138, 146, 135, 168, 162, 40,
    -- filter=20 channel=2
    47, 31, -186, -103, 8, -102, 122, 210, -295,
    -- filter=20 channel=3
    -85, -108, -196, 24, 218, 139, 121, -21, 134,
    -- filter=20 channel=4
    -84, 123, 115, -50, 152, 47, 60, -194, 149,
    -- filter=20 channel=5
    135, 2, -7, 67, -80, -66, -181, -18, -394,
    -- filter=20 channel=6
    -36, -9, -25, 18, -6, -142, 99, -303, 41,
    -- filter=20 channel=7
    -361, -251, 2, -186, 143, 92, 15, 25, 143,
    -- filter=20 channel=8
    77, 97, 26, -94, -76, -95, -272, 77, -78,
    -- filter=20 channel=9
    178, 46, 28, -50, 80, 5, -112, -202, -84,
    -- filter=20 channel=10
    24, -87, -23, 87, -92, 126, -105, 48, 169,
    -- filter=20 channel=11
    -11, -99, -19, 87, 0, -19, -90, 9, 11,
    -- filter=20 channel=12
    -30, 116, 73, 0, 4, -212, -180, -119, 96,
    -- filter=20 channel=13
    17, 12, 0, 4, -15, 9, -8, -19, -6,
    -- filter=20 channel=14
    10, 212, 91, 140, -32, -85, -130, -225, -173,
    -- filter=20 channel=15
    -130, -335, -21, -2, 10, 121, 149, 86, 123,
    -- filter=20 channel=16
    88, -48, -54, -256, -110, -39, 50, 51, -55,
    -- filter=20 channel=17
    119, -106, -138, 44, -79, -96, -90, 128, 86,
    -- filter=20 channel=18
    -26, 66, -163, -108, -21, 113, 31, -97, 63,
    -- filter=20 channel=19
    10, -168, 58, -90, 65, 136, -178, 129, -20,
    -- filter=20 channel=20
    -134, 98, -5, -87, -251, 66, 66, -101, 112,
    -- filter=20 channel=21
    -15, -176, 67, 18, 9, 131, -171, -20, 116,
    -- filter=20 channel=22
    119, -96, -6, -40, -140, -158, 69, -35, -71,
    -- filter=20 channel=23
    -136, -89, -32, 68, 186, -39, -10, 20, -28,
    -- filter=20 channel=24
    -144, -100, -38, -19, 30, 104, 199, 255, 272,
    -- filter=20 channel=25
    4, 78, -194, -206, -146, 7, 218, 43, 17,
    -- filter=20 channel=26
    95, 112, 69, -75, -17, -46, -28, -76, 142,
    -- filter=20 channel=27
    128, 149, 98, -63, 165, -27, -28, -141, 4,
    -- filter=20 channel=28
    130, 7, -6, 66, -154, -65, -89, 97, 5,
    -- filter=20 channel=29
    176, 89, 12, 58, 11, -149, 28, 46, 25,
    -- filter=20 channel=30
    -101, -275, -124, 16, 13, 18, -31, -122, 195,
    -- filter=20 channel=31
    -17, -25, -12, -16, -89, 37, 111, 36, 34,
    -- filter=21 channel=0
    -7, 17, -2, -11, -17, 3, -2, -26, -2,
    -- filter=21 channel=1
    -26, 7, -22, 11, -11, -21, 2, -32, -1,
    -- filter=21 channel=2
    -2, 1, -2, -5, 13, 3, -8, -9, 2,
    -- filter=21 channel=3
    -28, 0, -6, 7, -10, -7, 2, 4, -12,
    -- filter=21 channel=4
    14, -1, -24, -14, -1, -17, -8, 11, 14,
    -- filter=21 channel=5
    -25, -20, -17, -2, -3, 0, -20, -28, 2,
    -- filter=21 channel=6
    -3, -10, 2, -31, -11, -22, 0, 18, -25,
    -- filter=21 channel=7
    6, -22, 10, -8, 3, 17, 3, -18, 2,
    -- filter=21 channel=8
    3, 5, 13, -4, -8, -7, -23, -3, -21,
    -- filter=21 channel=9
    -21, -12, -13, -6, 0, -18, -11, -24, 0,
    -- filter=21 channel=10
    -6, -4, -14, -15, -21, 7, -12, 11, -23,
    -- filter=21 channel=11
    3, 0, -10, -17, -22, -10, -12, 11, -13,
    -- filter=21 channel=12
    4, -7, -9, -15, -16, 9, -35, 12, -14,
    -- filter=21 channel=13
    -3, 14, 4, 14, -7, 8, -17, 15, -19,
    -- filter=21 channel=14
    0, -11, -5, -7, 5, -4, 14, -17, -5,
    -- filter=21 channel=15
    -27, -10, -3, -25, 0, 7, -26, -13, -21,
    -- filter=21 channel=16
    -22, -1, -14, -7, -4, -3, 0, -4, 0,
    -- filter=21 channel=17
    5, -21, -3, 0, 15, -1, 19, 6, 11,
    -- filter=21 channel=18
    -3, 0, -10, -14, -24, -19, 1, -7, -3,
    -- filter=21 channel=19
    0, 7, 0, -12, -11, -9, -17, 1, -5,
    -- filter=21 channel=20
    -8, 0, -5, 0, 7, -14, -24, -19, 10,
    -- filter=21 channel=21
    3, -6, -11, -10, -8, -18, 10, -17, -25,
    -- filter=21 channel=22
    -24, 10, -6, -6, -2, -2, -1, -11, -18,
    -- filter=21 channel=23
    -22, -20, -15, -24, -13, -2, -9, 1, -4,
    -- filter=21 channel=24
    3, -20, -9, -11, 19, -1, 2, -7, -22,
    -- filter=21 channel=25
    -14, 1, 8, 12, 8, 5, -26, 10, -7,
    -- filter=21 channel=26
    0, 0, -23, -28, -3, -28, 0, -12, 1,
    -- filter=21 channel=27
    3, -15, 7, -6, -4, 0, -20, -10, -2,
    -- filter=21 channel=28
    -1, -11, 6, 0, -12, 8, 2, -18, 0,
    -- filter=21 channel=29
    6, 3, 7, 1, 1, 10, -19, -27, 0,
    -- filter=21 channel=30
    17, 20, -22, -14, -3, 5, -17, -15, 0,
    -- filter=21 channel=31
    7, -13, -29, 9, -32, 4, -33, -10, -8,
    -- filter=22 channel=0
    33, -124, -99, -1, -70, 1, -30, -110, -36,
    -- filter=22 channel=1
    -14, 171, -14, -139, 58, 46, -17, -90, -198,
    -- filter=22 channel=2
    76, 78, -42, 15, 44, 75, 0, -123, 97,
    -- filter=22 channel=3
    -130, 134, -75, 47, 100, 38, 13, -31, -187,
    -- filter=22 channel=4
    16, 1, -17, -45, 32, -113, -92, 142, 117,
    -- filter=22 channel=5
    0, 7, -127, 138, 7, -26, -14, 8, 81,
    -- filter=22 channel=6
    -47, -71, 83, -291, 17, 27, -192, 201, 84,
    -- filter=22 channel=7
    46, 90, -17, 102, 221, 7, -48, -72, -55,
    -- filter=22 channel=8
    -101, 16, -220, -143, 9, 72, -45, -139, 130,
    -- filter=22 channel=9
    -35, -302, -82, 41, -86, -174, -16, 117, 165,
    -- filter=22 channel=10
    -62, -31, 200, 10, -3, -54, 19, 56, 11,
    -- filter=22 channel=11
    -81, 126, -54, 152, 131, 22, -208, -169, 17,
    -- filter=22 channel=12
    41, -310, -180, 20, 8, -89, 160, 256, 18,
    -- filter=22 channel=13
    12, -6, -7, 13, -21, 9, 20, 6, -1,
    -- filter=22 channel=14
    -94, -150, -104, -64, 38, 86, -2, -105, -71,
    -- filter=22 channel=15
    -81, 252, -163, -112, 0, -24, 32, -296, -186,
    -- filter=22 channel=16
    63, 93, -7, 41, 59, 133, 5, 57, -25,
    -- filter=22 channel=17
    -50, -197, -184, -129, 366, -109, 56, -131, 179,
    -- filter=22 channel=18
    -143, 58, -24, -191, 13, -166, -24, 63, -209,
    -- filter=22 channel=19
    -78, 67, -11, -59, 52, 84, -163, 66, -24,
    -- filter=22 channel=20
    52, 175, 59, 115, 61, 3, -61, -164, -123,
    -- filter=22 channel=21
    -219, -161, -218, -55, 220, -92, 5, 11, -30,
    -- filter=22 channel=22
    87, -54, 210, 54, 41, -86, -77, 67, 90,
    -- filter=22 channel=23
    -35, -85, -252, 118, 101, -41, 84, 8, 18,
    -- filter=22 channel=24
    -175, 46, 92, -124, 78, 122, 69, 54, 42,
    -- filter=22 channel=25
    -13, 92, -20, -11, -135, 65, -59, -49, 132,
    -- filter=22 channel=26
    17, 249, 32, -59, 72, 109, -87, -406, -174,
    -- filter=22 channel=27
    94, -239, -119, 111, -31, -140, 119, -31, 105,
    -- filter=22 channel=28
    -224, -199, -314, 6, -216, -44, 236, 127, 92,
    -- filter=22 channel=29
    76, -229, -63, 83, 121, 63, 8, -131, 69,
    -- filter=22 channel=30
    -13, -122, -359, 190, 150, -97, -102, 134, 7,
    -- filter=22 channel=31
    95, -333, -81, -156, 223, 10, -129, 253, 90,
    -- filter=23 channel=0
    62, -74, 43, 67, 32, 195, -67, -59, 153,
    -- filter=23 channel=1
    59, -44, 68, 41, 49, -61, -74, -20, 130,
    -- filter=23 channel=2
    46, -24, -39, 54, 55, -231, -169, -128, 58,
    -- filter=23 channel=3
    295, -141, -68, -280, 74, -69, 118, 105, -123,
    -- filter=23 channel=4
    116, -169, -2, -64, -170, 9, 16, 4, -8,
    -- filter=23 channel=5
    -104, -361, -152, 125, -117, -36, 114, -60, -95,
    -- filter=23 channel=6
    -128, -107, 72, -245, 42, -111, 84, -62, -145,
    -- filter=23 channel=7
    277, -33, -80, 160, 39, 122, 153, -30, 55,
    -- filter=23 channel=8
    63, -90, -61, -48, -119, -66, -144, -49, -73,
    -- filter=23 channel=9
    89, 40, 67, 6, 67, 99, -118, 68, -115,
    -- filter=23 channel=10
    176, 25, 180, 3, 109, -7, 25, 25, 69,
    -- filter=23 channel=11
    -49, -25, 0, -15, -165, 197, 60, 23, -4,
    -- filter=23 channel=12
    43, 36, 59, -20, 245, 150, 165, 185, -33,
    -- filter=23 channel=13
    3, -20, 4, -30, 0, 23, -9, -6, -24,
    -- filter=23 channel=14
    155, -55, 125, -130, -118, -59, -115, -172, 75,
    -- filter=23 channel=15
    -15, 124, -190, -31, 94, 42, -131, 130, -35,
    -- filter=23 channel=16
    -331, -126, -86, -161, -144, -82, -225, 52, 21,
    -- filter=23 channel=17
    -135, 122, -9, -66, 127, -148, 89, 7, 183,
    -- filter=23 channel=18
    -124, 44, -224, 2, 103, 195, 108, -24, 49,
    -- filter=23 channel=19
    -25, 168, -22, -55, 207, 120, 217, -264, 65,
    -- filter=23 channel=20
    -112, -254, 30, -210, 272, -24, -4, 54, -54,
    -- filter=23 channel=21
    270, -142, -62, -275, 16, 149, 115, -200, 193,
    -- filter=23 channel=22
    185, -111, 4, -39, -131, -72, -145, 117, -671,
    -- filter=23 channel=23
    97, -5, -107, -31, 96, -63, 130, -103, 85,
    -- filter=23 channel=24
    -81, -223, -23, -23, 26, 149, 200, -82, -79,
    -- filter=23 channel=25
    -297, -9, -520, -152, -69, 134, 35, -160, 110,
    -- filter=23 channel=26
    2, -80, -142, -161, 77, -48, 61, 194, 163,
    -- filter=23 channel=27
    16, 6, -245, -26, -193, -305, 44, -37, -2,
    -- filter=23 channel=28
    -251, -10, -161, -117, -285, -30, -74, 177, -374,
    -- filter=23 channel=29
    100, 198, 86, 58, 31, 80, 45, 22, 66,
    -- filter=23 channel=30
    -336, -109, 75, -242, -271, 55, -60, -7, 90,
    -- filter=23 channel=31
    -161, 94, 162, -28, -5, 89, -53, -148, 1,
    -- filter=24 channel=0
    112, -173, 48, 59, -103, -7, -170, 55, 17,
    -- filter=24 channel=1
    -154, 63, -50, -55, 51, -181, 302, 43, 118,
    -- filter=24 channel=2
    34, 27, -219, -101, -12, 39, 128, 96, 30,
    -- filter=24 channel=3
    1, -51, 155, -136, -90, 4, -62, 24, -123,
    -- filter=24 channel=4
    120, 0, -84, 48, -108, -182, 21, -157, 38,
    -- filter=24 channel=5
    129, -58, -64, 13, 35, -123, 134, -82, -131,
    -- filter=24 channel=6
    52, 127, -187, -40, -36, -55, 1, -55, -72,
    -- filter=24 channel=7
    16, -192, -115, -75, -79, 2, -11, -75, 21,
    -- filter=24 channel=8
    18, -110, -86, -134, -118, 20, 182, 183, -49,
    -- filter=24 channel=9
    146, -136, 19, -86, -28, -129, 184, 37, 68,
    -- filter=24 channel=10
    -8, -11, 72, 17, 88, 214, 64, -104, 1,
    -- filter=24 channel=11
    -227, -8, -11, -32, -8, 43, 114, 144, 40,
    -- filter=24 channel=12
    -9, 129, 51, 129, 69, 45, -27, 65, -49,
    -- filter=24 channel=13
    -10, -4, -7, 0, -6, 17, -14, 0, 0,
    -- filter=24 channel=14
    -137, -118, -47, 71, -27, -98, 78, 14, 61,
    -- filter=24 channel=15
    -80, -101, 111, -107, -156, -34, 100, 51, 80,
    -- filter=24 channel=16
    68, -102, 41, -11, -73, 31, 111, 57, -15,
    -- filter=24 channel=17
    -135, 210, -190, 104, 72, 50, 206, 190, 80,
    -- filter=24 channel=18
    169, 91, -41, 98, -255, 65, -45, -23, 10,
    -- filter=24 channel=19
    105, 19, 100, -42, 33, -38, 67, -233, 22,
    -- filter=24 channel=20
    -130, -200, -51, -166, 91, 24, 53, 250, 99,
    -- filter=24 channel=21
    54, -121, -229, 11, 173, 22, -122, -63, 148,
    -- filter=24 channel=22
    83, -183, -3, -63, 7, 75, 110, -142, -201,
    -- filter=24 channel=23
    -239, 11, 126, -8, 7, 116, 51, -99, -74,
    -- filter=24 channel=24
    -108, 358, 31, 37, 108, -24, -290, 106, 163,
    -- filter=24 channel=25
    -45, -160, 9, 141, 77, 48, 99, -174, 90,
    -- filter=24 channel=26
    -176, 56, 166, 146, 152, -31, -6, -1, -221,
    -- filter=24 channel=27
    22, 56, 47, 12, 97, -136, -56, -105, 13,
    -- filter=24 channel=28
    197, 88, -118, -171, 135, 141, -130, -181, 3,
    -- filter=24 channel=29
    -49, 55, 36, -172, -32, 142, -244, -111, 28,
    -- filter=24 channel=30
    -362, 71, -97, -342, 111, -16, -19, 61, 31,
    -- filter=24 channel=31
    137, 92, 259, 59, 105, -88, -241, -550, -64,
    -- filter=25 channel=0
    152, 179, -48, 28, 113, 91, -93, 0, -58,
    -- filter=25 channel=1
    58, 82, 125, -164, 16, -47, -384, 24, -243,
    -- filter=25 channel=2
    -103, -43, 161, 286, 156, 66, 13, -31, 39,
    -- filter=25 channel=3
    20, 188, 37, -49, 70, 98, -10, -88, -35,
    -- filter=25 channel=4
    -12, 147, 35, 70, 162, -1, 209, -25, 103,
    -- filter=25 channel=5
    -1, -166, -21, -234, -43, 98, -255, -54, -19,
    -- filter=25 channel=6
    -78, -134, 95, -78, -12, 35, 157, -7, 74,
    -- filter=25 channel=7
    -12, -100, -128, 78, 112, -23, 108, 70, -142,
    -- filter=25 channel=8
    69, -157, -234, 10, 69, 8, -46, -80, 69,
    -- filter=25 channel=9
    98, 122, 166, 252, 224, 11, 4, 16, -94,
    -- filter=25 channel=10
    -16, 95, -17, 89, 49, -5, -67, 14, -62,
    -- filter=25 channel=11
    -14, -161, -99, 82, 83, -134, 165, 88, -25,
    -- filter=25 channel=12
    12, 67, 167, 16, 61, -74, -133, -131, -6,
    -- filter=25 channel=13
    21, 20, 16, 13, -15, -8, -7, -1, -8,
    -- filter=25 channel=14
    27, 152, 53, 67, 112, 206, -224, -174, -48,
    -- filter=25 channel=15
    -41, 72, -189, 94, 49, -35, 153, 14, -49,
    -- filter=25 channel=16
    23, -97, 151, 38, -28, -49, 116, -16, 11,
    -- filter=25 channel=17
    -236, 131, 110, 97, -96, 223, -57, 100, 356,
    -- filter=25 channel=18
    -45, -332, -85, -116, 59, 0, 18, -25, 80,
    -- filter=25 channel=19
    123, 84, -182, 113, 78, 91, 55, 74, 85,
    -- filter=25 channel=20
    -112, 21, -54, 68, 69, 25, -50, -73, 89,
    -- filter=25 channel=21
    16, 80, 43, 59, 152, 52, 96, -66, -228,
    -- filter=25 channel=22
    28, -207, -74, -110, 29, 25, -48, -237, 29,
    -- filter=25 channel=23
    -134, 8, -88, 165, 128, -8, 38, 38, 0,
    -- filter=25 channel=24
    -65, 60, -165, 168, 89, -32, -25, 142, -3,
    -- filter=25 channel=25
    -15, 41, -14, -129, -187, -238, 117, 130, -57,
    -- filter=25 channel=26
    3, 20, -39, -1, -3, 27, -123, 82, -150,
    -- filter=25 channel=27
    -199, 74, -17, -46, -168, -235, -159, -405, 13,
    -- filter=25 channel=28
    73, -85, -91, 39, 36, 98, -2, 6, 60,
    -- filter=25 channel=29
    53, 66, -15, -60, -72, 51, -29, -250, -23,
    -- filter=25 channel=30
    -1, 104, -31, 133, 104, 82, 53, -3, -83,
    -- filter=25 channel=31
    22, 7, 109, -116, -152, -152, 153, -40, -169,
    -- filter=26 channel=0
    -22, -24, -14, 142, -16, -163, 4, 61, -33,
    -- filter=26 channel=1
    178, -130, -41, 58, 91, -3, -164, 16, 177,
    -- filter=26 channel=2
    -89, 44, 136, -113, -17, 17, -115, 5, 134,
    -- filter=26 channel=3
    -159, 87, -39, -33, 184, -191, 115, 80, -5,
    -- filter=26 channel=4
    -219, 109, -114, -3, -61, -68, -10, -29, 158,
    -- filter=26 channel=5
    68, -17, -157, 172, -66, 83, 30, 103, 23,
    -- filter=26 channel=6
    101, 19, -116, 107, 38, -53, 156, 92, -19,
    -- filter=26 channel=7
    7, 81, -88, 63, -58, 37, -52, 28, -124,
    -- filter=26 channel=8
    -96, -191, -125, 116, -106, -67, 101, -175, -27,
    -- filter=26 channel=9
    10, 87, 14, -2, 157, 15, -97, -80, -34,
    -- filter=26 channel=10
    -33, 83, 97, 12, 60, 13, -31, 49, -190,
    -- filter=26 channel=11
    117, -18, -217, -64, -201, -70, 32, 4, 88,
    -- filter=26 channel=12
    -25, 85, 135, -64, 1, 72, 22, 159, 71,
    -- filter=26 channel=13
    -3, -4, 8, -1, -14, 7, 0, 1, 2,
    -- filter=26 channel=14
    -74, 9, -131, -87, -51, -111, 74, 98, 52,
    -- filter=26 channel=15
    -37, -71, 156, -18, 15, -15, 125, 83, -242,
    -- filter=26 channel=16
    91, -93, -29, -100, 161, -144, 14, -226, -43,
    -- filter=26 channel=17
    121, 55, -108, 57, 182, -53, -197, 5, 109,
    -- filter=26 channel=18
    -76, 67, -17, 31, 62, 35, -155, -5, 13,
    -- filter=26 channel=19
    -3, -130, 103, -39, 140, 38, 69, 24, 90,
    -- filter=26 channel=20
    -30, 186, 114, -334, -123, 215, 143, 61, -62,
    -- filter=26 channel=21
    246, -126, -142, 21, -38, -205, 4, -177, -191,
    -- filter=26 channel=22
    -167, 8, 213, 68, -12, -34, -45, -21, 25,
    -- filter=26 channel=23
    172, 100, -44, 138, 34, -92, 137, -43, 55,
    -- filter=26 channel=24
    -59, 142, -75, 173, 56, -322, 59, -149, -8,
    -- filter=26 channel=25
    161, -16, 99, -185, 72, -58, -266, 63, -78,
    -- filter=26 channel=26
    -89, -49, 92, -220, 30, 216, -184, -233, 240,
    -- filter=26 channel=27
    -7, 102, -38, -23, -17, -81, -270, -146, 118,
    -- filter=26 channel=28
    -21, 12, 65, 79, 118, -470, 139, -3, 125,
    -- filter=26 channel=29
    211, 77, -18, -22, -7, -65, 62, -83, -71,
    -- filter=26 channel=30
    175, -256, 48, 8, -103, -83, -36, 164, 137,
    -- filter=26 channel=31
    113, 54, -179, 157, 205, -233, 70, 5, -176,
    -- filter=27 channel=0
    -152, -126, 17, 153, -99, 5, 43, 108, 134,
    -- filter=27 channel=1
    -138, -6, -212, -85, 75, -115, 107, 147, 87,
    -- filter=27 channel=2
    34, 164, -245, 143, 259, 25, -438, -15, 70,
    -- filter=27 channel=3
    13, -88, -206, -71, 6, -220, -109, -59, -42,
    -- filter=27 channel=4
    4, 2, -47, -246, 55, -106, 31, 104, 114,
    -- filter=27 channel=5
    -63, -157, 27, 135, -62, -103, 27, 141, 183,
    -- filter=27 channel=6
    52, -49, 97, -45, 165, 30, 5, 170, 83,
    -- filter=27 channel=7
    0, -168, -61, -103, -219, -128, -205, -148, 187,
    -- filter=27 channel=8
    79, 80, -139, 114, 43, 14, 208, 9, 129,
    -- filter=27 channel=9
    -30, 49, 108, 122, 55, -106, 11, 44, -60,
    -- filter=27 channel=10
    -52, 38, -44, 73, -4, -79, 22, -76, -198,
    -- filter=27 channel=11
    -110, 97, 37, -3, 17, 99, 60, -150, -46,
    -- filter=27 channel=12
    -73, 139, -13, 140, -145, 67, 1, 0, -185,
    -- filter=27 channel=13
    12, 5, 15, 3, -11, -21, -11, -16, -19,
    -- filter=27 channel=14
    4, 56, 82, -7, 187, -25, -13, 204, 246,
    -- filter=27 channel=15
    -60, 109, 132, -110, 81, 98, -127, -226, -90,
    -- filter=27 channel=16
    40, 329, -70, -25, 176, 150, -232, -283, -63,
    -- filter=27 channel=17
    -34, 79, 193, 150, -183, -94, 3, -135, -82,
    -- filter=27 channel=18
    -141, -49, -154, -121, -29, 109, -71, -124, -195,
    -- filter=27 channel=19
    -37, 189, 22, -75, 110, 146, -117, -115, 140,
    -- filter=27 channel=20
    130, 62, 51, -101, 38, 141, -353, -34, -103,
    -- filter=27 channel=21
    -4, 129, 138, -127, 89, 37, -205, -188, -96,
    -- filter=27 channel=22
    26, 196, -46, 54, 206, -4, -238, 144, -10,
    -- filter=27 channel=23
    102, -99, 70, 124, -192, -207, 10, 55, 81,
    -- filter=27 channel=24
    -36, -50, -89, -155, -272, 117, 126, 47, -373,
    -- filter=27 channel=25
    97, -193, 157, -119, -206, 45, 166, -46, -141,
    -- filter=27 channel=26
    -109, -83, -9, 78, 91, -6, -215, 0, 25,
    -- filter=27 channel=27
    -53, -127, -3, -43, 70, 32, -141, 48, 133,
    -- filter=27 channel=28
    -149, -4, 2, -12, 93, -27, -181, 43, 246,
    -- filter=27 channel=29
    137, 79, 43, 22, 53, -146, 23, 85, 28,
    -- filter=27 channel=30
    -81, -20, -130, -59, -150, 21, -365, -162, -329,
    -- filter=27 channel=31
    143, 83, -7, -63, -90, -36, 85, -104, 65,
    -- filter=28 channel=0
    65, -44, 119, -135, 64, 102, -7, -20, 23,
    -- filter=28 channel=1
    -3, 265, -11, 34, -84, -123, -11, -43, 6,
    -- filter=28 channel=2
    -8, 49, 18, -5, 45, 176, -8, -24, -73,
    -- filter=28 channel=3
    2, -227, -67, 24, -130, -133, 55, -76, -32,
    -- filter=28 channel=4
    109, -67, -115, 87, 78, -9, 67, 48, -102,
    -- filter=28 channel=5
    97, 74, -66, -247, 94, -13, 85, 74, 102,
    -- filter=28 channel=6
    79, -235, -141, -243, 20, -21, 32, -24, -30,
    -- filter=28 channel=7
    89, 40, 25, -133, -81, -122, -116, -218, -142,
    -- filter=28 channel=8
    -116, 91, 32, 20, -244, 35, -72, 109, -76,
    -- filter=28 channel=9
    121, -87, 26, -95, -17, 58, 9, -70, 58,
    -- filter=28 channel=10
    -69, 123, 217, -63, -86, 206, 77, 47, 88,
    -- filter=28 channel=11
    -21, -13, -189, 86, 82, -129, 213, 3, 26,
    -- filter=28 channel=12
    -23, -23, 58, 58, -55, 70, 52, 144, 56,
    -- filter=28 channel=13
    1, 10, -8, -8, 21, 16, 21, -7, 9,
    -- filter=28 channel=14
    45, -153, -102, -38, 34, 15, 18, -3, 111,
    -- filter=28 channel=15
    -23, 23, 64, -54, 14, 65, -115, 65, 45,
    -- filter=28 channel=16
    5, -110, -496, -78, -132, -170, -33, -95, -267,
    -- filter=28 channel=17
    -40, -34, -225, -1, -285, -185, -52, -34, -231,
    -- filter=28 channel=18
    -104, -59, -65, 193, -84, 25, 55, -60, 2,
    -- filter=28 channel=19
    261, -68, -115, -188, -239, 54, 194, -95, 6,
    -- filter=28 channel=20
    -65, -26, 56, -30, -201, 112, 89, 19, 43,
    -- filter=28 channel=21
    -320, 26, -20, 70, 12, -290, -46, -44, -196,
    -- filter=28 channel=22
    57, -167, 97, 229, -15, -61, -91, 17, -54,
    -- filter=28 channel=23
    66, -39, 18, -20, 51, -154, -17, -145, 14,
    -- filter=28 channel=24
    105, 19, 102, -158, -125, -13, -184, -56, -158,
    -- filter=28 channel=25
    -283, -262, -76, -261, -223, -90, -1, -173, -277,
    -- filter=28 channel=26
    42, -326, -29, -158, -152, -42, -52, 7, -295,
    -- filter=28 channel=27
    70, -49, 241, 4, 75, 150, -54, -111, 68,
    -- filter=28 channel=28
    121, -20, -104, 106, -84, -40, 67, -72, 71,
    -- filter=28 channel=29
    70, 51, 12, -108, -33, -16, -83, -45, -108,
    -- filter=28 channel=30
    -136, 226, 28, 174, -43, -137, -19, -27, 39,
    -- filter=28 channel=31
    -80, 97, 28, 3, 5, 139, 32, 18, -20,
    -- filter=29 channel=0
    15, -18, 6, 63, -90, 135, -205, 124, 209,
    -- filter=29 channel=1
    -30, 81, -76, -313, 225, -154, 91, 176, -159,
    -- filter=29 channel=2
    76, -117, -155, 35, -2, 7, -100, 163, -70,
    -- filter=29 channel=3
    171, 29, -148, 0, 102, -23, -14, 189, -18,
    -- filter=29 channel=4
    25, -3, 10, -29, 55, 1, 47, 30, 131,
    -- filter=29 channel=5
    -60, -18, 108, -212, -210, 97, -213, -107, -68,
    -- filter=29 channel=6
    -192, 50, 108, -131, -243, -108, -69, -50, -77,
    -- filter=29 channel=7
    6, -243, 44, -216, -144, -306, -335, -96, -148,
    -- filter=29 channel=8
    112, -257, 112, 74, -56, -256, 10, -23, -39,
    -- filter=29 channel=9
    227, 248, -11, 13, 240, 41, -58, -34, -11,
    -- filter=29 channel=10
    -74, 148, 102, -111, 41, 219, -129, 66, 4,
    -- filter=29 channel=11
    -226, -41, 150, 17, 43, 54, 15, -26, -43,
    -- filter=29 channel=12
    -48, 0, -160, 63, -28, -26, -17, 15, -207,
    -- filter=29 channel=13
    12, -5, 4, 8, 4, -16, -9, 6, 6,
    -- filter=29 channel=14
    -33, -67, 92, 65, 181, 71, -82, -57, 173,
    -- filter=29 channel=15
    89, -84, -111, 33, 50, 57, 26, 82, -125,
    -- filter=29 channel=16
    1, 19, 0, -135, -82, 24, -49, -84, -52,
    -- filter=29 channel=17
    0, -57, -243, -41, -354, -164, 323, 194, 10,
    -- filter=29 channel=18
    37, -104, 116, 53, -27, -152, -177, 127, 77,
    -- filter=29 channel=19
    198, 35, -185, -10, 68, -107, 54, 88, -52,
    -- filter=29 channel=20
    34, 51, -7, 184, 50, -111, -28, 55, 0,
    -- filter=29 channel=21
    101, -113, -99, 0, 112, -71, -9, -106, -90,
    -- filter=29 channel=22
    40, -89, -20, 107, 80, -157, -187, -298, 5,
    -- filter=29 channel=23
    -161, -51, 123, 99, 13, -25, -20, 65, 90,
    -- filter=29 channel=24
    -70, 99, -100, 57, -56, -155, 11, 31, 74,
    -- filter=29 channel=25
    -4, 8, -34, -73, -88, -185, 0, 14, -6,
    -- filter=29 channel=26
    -51, 0, 124, 219, -21, -104, -108, 184, 246,
    -- filter=29 channel=27
    -46, -42, 116, -162, -134, 48, 11, 94, 16,
    -- filter=29 channel=28
    100, 106, 33, -207, 69, -6, 30, 24, 174,
    -- filter=29 channel=29
    -31, -155, 18, 36, 98, -41, 137, -39, 61,
    -- filter=29 channel=30
    -140, -117, -55, -226, 276, 142, -158, -7, -122,
    -- filter=29 channel=31
    -64, -117, 8, -56, 4, 106, -145, -177, 193,
    -- filter=30 channel=0
    -75, 140, 173, -1, 109, 82, -463, -149, -49,
    -- filter=30 channel=1
    -105, -18, 47, 89, -84, 63, -145, 0, -97,
    -- filter=30 channel=2
    -147, 48, 81, 60, 159, -112, -11, 79, -256,
    -- filter=30 channel=3
    88, -127, -50, 99, -48, -109, -20, -214, 127,
    -- filter=30 channel=4
    14, 34, 98, -12, -6, -319, -150, 43, 160,
    -- filter=30 channel=5
    -120, -79, -65, -170, -58, -23, 38, -99, -166,
    -- filter=30 channel=6
    -53, -91, 14, 73, -86, 114, 24, -95, 195,
    -- filter=30 channel=7
    -17, 27, 2, -14, -320, -14, -131, -21, 108,
    -- filter=30 channel=8
    -8, -16, 253, 1, -313, -92, -395, 110, 135,
    -- filter=30 channel=9
    161, 80, -184, -54, 126, 23, -342, -124, 61,
    -- filter=30 channel=10
    -255, 207, 69, -389, -212, -13, -168, -321, 31,
    -- filter=30 channel=11
    -83, -234, -38, 24, 66, 216, -55, 18, 101,
    -- filter=30 channel=12
    97, -123, -314, -114, 31, 2, -22, 14, -43,
    -- filter=30 channel=13
    12, 11, 13, 7, 10, 6, -7, -9, -3,
    -- filter=30 channel=14
    -1, 83, 111, -24, 160, 85, -218, -6, 34,
    -- filter=30 channel=15
    -160, -342, -87, -60, -192, -129, 67, 84, 140,
    -- filter=30 channel=16
    -230, 23, -102, 149, 61, 7, 98, -105, -233,
    -- filter=30 channel=17
    -306, 116, -209, -613, -474, 42, 135, 306, 104,
    -- filter=30 channel=18
    -83, -144, 99, 65, -4, 106, -327, -202, 77,
    -- filter=30 channel=19
    65, 9, -116, -15, 134, 106, 127, 25, 130,
    -- filter=30 channel=20
    20, -103, 188, 397, -178, -15, -71, 52, -141,
    -- filter=30 channel=21
    56, 51, 68, 37, -8, -87, 40, -56, 55,
    -- filter=30 channel=22
    158, -231, 123, -259, 17, -55, -60, 176, -478,
    -- filter=30 channel=23
    -53, 174, -73, -18, 122, -9, 158, -42, -119,
    -- filter=30 channel=24
    -129, -81, -94, 232, -37, -290, 239, 109, -18,
    -- filter=30 channel=25
    48, -180, -64, -33, -72, -212, -80, 211, 130,
    -- filter=30 channel=26
    93, -320, -50, -107, -119, 282, 68, -70, 78,
    -- filter=30 channel=27
    54, 104, -100, 75, 121, -79, 257, 126, 136,
    -- filter=30 channel=28
    0, 28, 55, -99, -99, -24, -63, 79, -260,
    -- filter=30 channel=29
    -40, -30, -62, 84, 105, 152, 138, 130, 1,
    -- filter=30 channel=30
    121, -69, 18, -180, -78, -38, -100, 13, -175,
    -- filter=30 channel=31
    -179, 127, -14, -97, 142, -203, 28, 101, 251,
    -- filter=31 channel=0
    81, 97, 51, 168, -20, -92, 43, -82, -30,
    -- filter=31 channel=1
    -59, -106, 159, 70, -242, 128, 200, -273, 38,
    -- filter=31 channel=2
    80, 105, 105, 91, -74, -125, -27, -31, -9,
    -- filter=31 channel=3
    -33, 200, -185, 235, 37, -135, -110, -444, -166,
    -- filter=31 channel=4
    -21, 104, 48, -88, 18, 72, -112, -79, 9,
    -- filter=31 channel=5
    -142, 9, -24, -15, 85, 48, 32, -147, 53,
    -- filter=31 channel=6
    -202, -29, -19, 25, -194, 26, 149, -116, 143,
    -- filter=31 channel=7
    -295, -95, -9, -293, -225, -8, -174, -5, 139,
    -- filter=31 channel=8
    -136, -321, -69, 13, 100, -21, 32, 139, -70,
    -- filter=31 channel=9
    138, -24, -273, -14, 63, 258, 202, -52, 14,
    -- filter=31 channel=10
    -8, 171, -20, -115, -73, -71, -55, 78, 124,
    -- filter=31 channel=11
    -127, 21, -132, -86, -150, 9, 103, 128, 58,
    -- filter=31 channel=12
    260, 105, -3, 52, -44, -39, -15, -12, -44,
    -- filter=31 channel=13
    -7, 9, -5, -19, -6, 13, -2, 20, -12,
    -- filter=31 channel=14
    90, 65, 70, 105, -32, -61, -21, -77, 46,
    -- filter=31 channel=15
    106, 18, 155, 1, 63, -73, 43, -116, -205,
    -- filter=31 channel=16
    69, 75, 14, -47, -73, 73, -88, -72, 18,
    -- filter=31 channel=17
    134, 18, 209, -178, 302, 39, -204, -178, -280,
    -- filter=31 channel=18
    -141, 164, -225, 5, 184, -75, -8, 140, -143,
    -- filter=31 channel=19
    -338, -158, -118, -283, 110, -191, -132, -197, 219,
    -- filter=31 channel=20
    -2, 120, 50, 108, -1, 50, 192, 58, 23,
    -- filter=31 channel=21
    -10, 63, -55, -259, 19, -61, -459, 65, 373,
    -- filter=31 channel=22
    -3, 25, 8, -57, 36, 134, -92, 321, -31,
    -- filter=31 channel=23
    253, 74, -74, -253, -27, -50, -116, 30, -221,
    -- filter=31 channel=24
    -77, 18, 80, 55, 32, 8, -1, -35, 125,
    -- filter=31 channel=25
    -34, 174, 87, -130, 61, 87, 194, -25, 38,
    -- filter=31 channel=26
    1, -1, 65, -7, 140, 154, -148, -114, -255,
    -- filter=31 channel=27
    63, 92, 62, -44, -21, 102, -19, -4, 116,
    -- filter=31 channel=28
    52, -118, -60, 74, 3, -52, 173, -286, 106,
    -- filter=31 channel=29
    -238, -205, -23, 64, -205, -79, 12, 73, -275,
    -- filter=31 channel=30
    -81, 157, -115, -144, -296, 40, -96, -4, -89,
    -- filter=31 channel=31
    -122, 21, -114, 2, 78, -150, -333, -67, 48,
    -- filter=32 channel=0
    -358, -374, -161, -156, -258, -256, 23, -27, -162,
    -- filter=32 channel=1
    68, -810, 359, 183, 174, -132, 18, 189, 199,
    -- filter=32 channel=2
    192, 123, -338, -12, 1, -30, -9, 87, 33,
    -- filter=32 channel=3
    -48, 36, 148, -56, 28, 162, -25, 39, 81,
    -- filter=32 channel=4
    232, -415, 56, 2, 241, -57, 4, 19, -151,
    -- filter=32 channel=5
    -410, -223, -349, -146, -127, 20, 104, 36, 164,
    -- filter=32 channel=6
    -9, -236, 29, -18, -70, -16, 90, -73, -16,
    -- filter=32 channel=7
    -108, -405, -46, -140, 96, 49, 42, -76, 151,
    -- filter=32 channel=8
    -63, 250, 11, 128, -43, -177, 70, -127, 224,
    -- filter=32 channel=9
    13, -561, -36, -104, 66, 284, -77, -154, 172,
    -- filter=32 channel=10
    -76, -58, 112, -199, -89, 138, 40, -205, 242,
    -- filter=32 channel=11
    56, -176, -52, 0, 20, 112, 70, 53, 33,
    -- filter=32 channel=12
    -48, -156, -435, 268, 270, -415, -78, -66, 145,
    -- filter=32 channel=13
    -19, 11, 17, -14, 4, 13, -10, 0, -15,
    -- filter=32 channel=14
    -195, -261, -55, 58, -265, -78, 125, -81, -12,
    -- filter=32 channel=15
    -74, 97, 188, 16, 87, 18, 17, -22, 7,
    -- filter=32 channel=16
    121, -171, -9, -61, -11, 115, -206, -94, 121,
    -- filter=32 channel=17
    298, -269, 28, -72, 28, 55, -191, 96, 140,
    -- filter=32 channel=18
    -8, -35, -53, -57, 18, 83, -20, 14, 0,
    -- filter=32 channel=19
    22, -393, 171, -74, 152, -37, 15, 60, 99,
    -- filter=32 channel=20
    32, 54, -107, -175, 68, -122, -71, -14, 158,
    -- filter=32 channel=21
    -155, 205, 108, 107, 40, -48, -68, 10, -83,
    -- filter=32 channel=22
    65, -197, 31, -66, -310, 465, -76, -31, 106,
    -- filter=32 channel=23
    119, -178, -594, 6, 137, 97, 102, 8, -181,
    -- filter=32 channel=24
    -110, 224, 178, -74, -29, 121, 100, -94, -183,
    -- filter=32 channel=25
    110, -278, -5, 174, 74, -66, -8, 40, 13,
    -- filter=32 channel=26
    -26, 31, -83, 163, -50, -131, 11, 44, 27,
    -- filter=32 channel=27
    103, 73, -137, 75, 55, -22, 52, -33, 138,
    -- filter=32 channel=28
    220, 4, -89, -73, 136, 23, 64, -11, -6,
    -- filter=32 channel=29
    -245, -281, -281, 215, -112, 102, 5, 101, -54,
    -- filter=32 channel=30
    -284, 149, 63, 20, -62, -34, -132, -8, -55,
    -- filter=32 channel=31
    -55, -23, 140, 10, 1, -160, 11, -134, 74,
    -- filter=33 channel=0
    115, 111, 130, 92, 151, 96, 20, 108, 130,
    -- filter=33 channel=1
    -16, -91, 68, -91, -126, 122, -90, 38, -7,
    -- filter=33 channel=2
    42, 5, -131, -212, 105, 167, -41, 134, 73,
    -- filter=33 channel=3
    -34, -52, -62, 3, 4, -19, 82, -67, 89,
    -- filter=33 channel=4
    -86, -153, -73, -119, -213, -275, -76, -164, -255,
    -- filter=33 channel=5
    117, -67, 137, 136, 114, -3, 225, 153, -29,
    -- filter=33 channel=6
    13, 1, 55, 67, -105, -105, -24, -106, -30,
    -- filter=33 channel=7
    40, 137, 48, 120, 136, 46, 107, -3, 97,
    -- filter=33 channel=8
    121, 66, 89, -11, 20, 71, 5, -150, 79,
    -- filter=33 channel=9
    47, -19, 46, -108, -1, -126, 68, 25, -158,
    -- filter=33 channel=10
    49, 132, 11, 242, 275, 170, 154, 132, 142,
    -- filter=33 channel=11
    -101, -116, 29, -136, -64, -150, -61, -8, -34,
    -- filter=33 channel=12
    45, -15, 52, -64, -1, -100, 52, -283, -97,
    -- filter=33 channel=13
    1, 4, -18, 9, -8, -3, 8, 26, 5,
    -- filter=33 channel=14
    -9, -9, -26, -55, -12, -113, -18, -8, -39,
    -- filter=33 channel=15
    78, -51, 85, -117, -99, 79, 28, -34, 92,
    -- filter=33 channel=16
    0, 133, 103, 20, 191, 34, -42, -82, 28,
    -- filter=33 channel=17
    -19, -348, -6, 136, 140, -269, 145, 225, -87,
    -- filter=33 channel=18
    7, 168, -101, 69, -2, -49, -82, 163, 144,
    -- filter=33 channel=19
    197, 72, -6, 57, 98, -31, -58, 133, 42,
    -- filter=33 channel=20
    -102, 155, -42, -102, 12, -103, -84, 57, -23,
    -- filter=33 channel=21
    4, 5, -4, -167, 6, 35, -152, -125, -9,
    -- filter=33 channel=22
    -120, 108, -38, -106, -2, 21, 213, -299, -8,
    -- filter=33 channel=23
    -27, -93, 38, -59, -48, -240, 82, 54, -194,
    -- filter=33 channel=24
    6, -53, -9, 31, 47, 37, -69, 20, -5,
    -- filter=33 channel=25
    4, -158, -115, -52, -10, -34, -87, -164, -50,
    -- filter=33 channel=26
    133, 18, 70, -32, -129, 92, -201, 45, -103,
    -- filter=33 channel=27
    -80, -67, -147, 0, -438, -31, -69, -42, -205,
    -- filter=33 channel=28
    -74, -2, -92, -72, -16, 41, 46, 60, 120,
    -- filter=33 channel=29
    -201, 84, -74, -159, -55, -82, 3, -271, -218,
    -- filter=33 channel=30
    -37, -135, -125, 160, 1, -1, -34, 258, 151,
    -- filter=33 channel=31
    -70, 159, 72, -12, 8, -15, -178, -93, 97,
    -- filter=34 channel=0
    -162, -79, -49, -48, 127, 75, -112, -135, 96,
    -- filter=34 channel=1
    -201, 161, -43, -110, -40, -172, 73, -24, -28,
    -- filter=34 channel=2
    103, 15, -36, -19, -3, -85, 10, -102, -13,
    -- filter=34 channel=3
    159, -184, -54, 264, 104, -56, -32, 27, -122,
    -- filter=34 channel=4
    -86, -28, -1, 95, 279, 122, 29, 45, -14,
    -- filter=34 channel=5
    -75, -78, 163, -94, 31, 10, 0, 26, 46,
    -- filter=34 channel=6
    40, -44, 10, 41, 86, 36, 167, -17, -113,
    -- filter=34 channel=7
    37, -120, 70, -53, -19, -157, 128, 10, -85,
    -- filter=34 channel=8
    -20, 117, 37, -330, -164, 13, 24, 204, -61,
    -- filter=34 channel=9
    -253, -5, -33, 19, 279, 256, -223, 134, 98,
    -- filter=34 channel=10
    -2, -15, -44, 24, -201, -67, 0, 145, 163,
    -- filter=34 channel=11
    41, 183, 37, 6, -218, -159, 149, 40, -13,
    -- filter=34 channel=12
    91, -79, -89, 65, 0, 15, -33, -41, -10,
    -- filter=34 channel=13
    8, 15, -20, 9, 18, -20, -19, 10, 7,
    -- filter=34 channel=14
    -53, -23, 59, -33, 15, 79, -193, -11, 239,
    -- filter=34 channel=15
    48, 86, -99, 111, 144, -20, -228, -129, 174,
    -- filter=34 channel=16
    89, 168, 110, 15, -114, -86, -86, 56, 145,
    -- filter=34 channel=17
    -18, -443, 7, 284, -246, 171, -95, 299, -74,
    -- filter=34 channel=18
    32, 29, -103, 18, -43, 26, -71, -123, -151,
    -- filter=34 channel=19
    206, -48, -127, -159, 35, -43, 22, 7, 127,
    -- filter=34 channel=20
    64, 138, -230, 66, -190, -204, -71, 12, -44,
    -- filter=34 channel=21
    91, -74, 108, 19, -36, -117, 123, -342, 79,
    -- filter=34 channel=22
    114, -69, -22, 89, 108, -19, -165, 121, 178,
    -- filter=34 channel=23
    31, 97, -126, -126, -82, -13, 73, 30, 150,
    -- filter=34 channel=24
    -140, 9, -154, -194, 214, -494, -23, 184, -150,
    -- filter=34 channel=25
    165, -15, -34, 28, 12, -90, 105, -61, -86,
    -- filter=34 channel=26
    29, 55, 57, 103, 95, -41, 44, -11, -143,
    -- filter=34 channel=27
    49, -73, -6, 115, -177, -111, -32, 112, 208,
    -- filter=34 channel=28
    -136, -198, 85, -58, 26, -60, 56, -66, 10,
    -- filter=34 channel=29
    60, -206, 166, -48, 3, 7, -32, 139, 24,
    -- filter=34 channel=30
    46, 95, -115, -62, -117, -221, 182, 131, 138,
    -- filter=34 channel=31
    -16, 33, -41, 166, 100, -5, -157, -74, -253,
    -- filter=35 channel=0
    2, -5, 12, -25, 5, -14, -21, -3, -21,
    -- filter=35 channel=1
    1, 6, -20, 2, -24, -2, -27, -1, -2,
    -- filter=35 channel=2
    -14, -16, 6, -34, -11, -13, -10, -18, 0,
    -- filter=35 channel=3
    -10, 14, -5, -7, 7, -9, -19, -10, 2,
    -- filter=35 channel=4
    8, 0, 5, -27, -21, -22, -25, 4, -25,
    -- filter=35 channel=5
    -12, -14, -2, -5, 9, 5, -13, -16, 12,
    -- filter=35 channel=6
    -16, -16, -4, -24, 12, -16, -5, -9, 9,
    -- filter=35 channel=7
    -13, -12, 16, -17, -1, 9, -24, -21, -14,
    -- filter=35 channel=8
    -29, 7, -5, -27, -6, -11, -8, -16, 0,
    -- filter=35 channel=9
    -17, -27, 1, -17, -26, 1, 5, -20, 9,
    -- filter=35 channel=10
    7, -8, -21, -11, 0, 4, -18, -21, -1,
    -- filter=35 channel=11
    1, -17, 1, -15, -24, -4, -31, -30, -19,
    -- filter=35 channel=12
    0, -23, -1, 0, -17, -28, -5, -17, -11,
    -- filter=35 channel=13
    -17, -3, 1, -12, 7, 6, -16, 9, 22,
    -- filter=35 channel=14
    -5, -12, -2, -22, -23, 14, -5, -13, 1,
    -- filter=35 channel=15
    -7, -16, -7, -19, -28, -9, 10, 0, -24,
    -- filter=35 channel=16
    -20, 7, -20, 4, -21, 0, -23, -12, -13,
    -- filter=35 channel=17
    1, -27, -4, 11, -10, 8, -3, -3, -17,
    -- filter=35 channel=18
    2, 9, 1, -23, 13, -9, -2, 13, 8,
    -- filter=35 channel=19
    2, -11, -11, 2, -17, -6, 9, -14, -24,
    -- filter=35 channel=20
    -23, -18, 9, 2, -14, -18, -8, -6, -26,
    -- filter=35 channel=21
    -8, -1, 6, 3, 8, -6, -4, -10, -12,
    -- filter=35 channel=22
    12, 14, -1, -20, 12, 3, -25, -10, -6,
    -- filter=35 channel=23
    -26, -19, -25, -10, -11, -8, -28, -17, -12,
    -- filter=35 channel=24
    -7, -13, -2, -12, -8, 9, -13, -17, -5,
    -- filter=35 channel=25
    2, 0, -16, 0, 11, 7, 9, -4, -19,
    -- filter=35 channel=26
    16, 4, -29, 18, -11, -13, -5, -9, 12,
    -- filter=35 channel=27
    -9, 7, -15, -6, 2, -12, 5, -24, -8,
    -- filter=35 channel=28
    5, 8, -23, 4, -19, 0, -14, -2, 10,
    -- filter=35 channel=29
    -7, 7, -31, 16, -4, -10, -9, -5, 7,
    -- filter=35 channel=30
    9, -20, -20, 4, 1, 5, -15, -22, 11,
    -- filter=35 channel=31
    -3, -1, -18, -13, -25, -29, -18, -20, -32,
    -- filter=36 channel=0
    62, -11, -86, -18, -45, 116, 87, 137, 102,
    -- filter=36 channel=1
    130, -65, 50, -18, 151, -426, -29, 40, -33,
    -- filter=36 channel=2
    -129, 153, 56, 113, -88, -136, 307, -174, -375,
    -- filter=36 channel=3
    -29, -32, 154, -205, -90, -86, -10, -82, 24,
    -- filter=36 channel=4
    -174, 89, 120, -240, 153, 112, -32, 10, 20,
    -- filter=36 channel=5
    23, -173, -193, 84, 20, -22, 100, 38, 150,
    -- filter=36 channel=6
    -48, 1, -130, -10, 124, -32, -23, 23, -21,
    -- filter=36 channel=7
    54, -209, -1, 43, -88, -37, 240, -51, -38,
    -- filter=36 channel=8
    -139, 6, 96, 67, -70, 255, -50, 141, -62,
    -- filter=36 channel=9
    -56, -44, -121, 26, 111, 86, -3, -40, -9,
    -- filter=36 channel=10
    14, -295, -241, 18, -58, -74, -10, 131, 133,
    -- filter=36 channel=11
    163, 53, -90, 11, 22, 145, 11, 4, -176,
    -- filter=36 channel=12
    29, 147, 13, 34, 14, 16, -153, -105, -51,
    -- filter=36 channel=13
    -23, 4, 4, -6, -8, -14, -4, 8, -9,
    -- filter=36 channel=14
    -100, 140, -17, -16, 161, 40, 64, 48, 20,
    -- filter=36 channel=15
    -104, 84, 220, -23, 3, 213, -13, 0, 94,
    -- filter=36 channel=16
    -104, -250, -299, -151, -83, -33, -42, 6, 24,
    -- filter=36 channel=17
    191, -38, 18, 156, 130, 0, 6, 4, -194,
    -- filter=36 channel=18
    37, -203, 42, 132, 92, 107, 26, 154, -38,
    -- filter=36 channel=19
    -23, -15, -55, -156, 98, 40, 79, -116, 11,
    -- filter=36 channel=20
    149, -141, -180, -24, -89, -11, 212, 79, -194,
    -- filter=36 channel=21
    -88, 86, 137, 12, 67, -40, -168, -81, 125,
    -- filter=36 channel=22
    126, -173, -13, -278, 32, 88, -216, 147, 97,
    -- filter=36 channel=23
    -8, -35, -31, 105, -72, 20, -41, 72, 27,
    -- filter=36 channel=24
    -113, 73, -142, -70, -33, -298, 39, -63, -97,
    -- filter=36 channel=25
    -57, 77, 17, 39, -51, -29, 77, 63, -266,
    -- filter=36 channel=26
    60, -70, 43, 114, -101, -14, -86, -174, -80,
    -- filter=36 channel=27
    -55, 47, 18, -76, -23, 13, -210, -10, -12,
    -- filter=36 channel=28
    113, 31, -117, -80, 79, 2, 51, -29, 66,
    -- filter=36 channel=29
    155, -38, 127, -51, 1, -4, -104, 145, 55,
    -- filter=36 channel=30
    108, -16, -110, -20, 20, -126, -92, -72, 137,
    -- filter=36 channel=31
    17, 101, -70, -89, -62, -74, 111, -4, 143,
    -- filter=37 channel=0
    182, 83, -19, -227, -371, -113, -162, -236, -113,
    -- filter=37 channel=1
    -47, 101, 5, 32, -177, 157, 39, 81, -90,
    -- filter=37 channel=2
    -71, -13, 5, -72, -58, 122, 194, 67, -29,
    -- filter=37 channel=3
    84, -67, 298, 43, -34, 44, 33, -97, -158,
    -- filter=37 channel=4
    -193, -49, -23, 15, -270, -92, 118, -178, -114,
    -- filter=37 channel=5
    164, 94, 155, -60, 82, 25, -4, 57, 12,
    -- filter=37 channel=6
    104, 83, 87, 210, 165, -73, -64, 95, 18,
    -- filter=37 channel=7
    143, -85, -16, -10, -31, 125, -56, -79, -42,
    -- filter=37 channel=8
    81, -64, -66, -112, -40, -6, -232, 46, -38,
    -- filter=37 channel=9
    19, 6, -69, -407, -107, -134, 2, -153, 173,
    -- filter=37 channel=10
    65, -36, -76, 61, 120, 69, -10, 106, 0,
    -- filter=37 channel=11
    98, 98, -5, 86, -189, -68, 11, -11, -66,
    -- filter=37 channel=12
    -12, -51, -140, 46, -181, 76, 24, 173, 16,
    -- filter=37 channel=13
    7, -8, -11, -13, -18, -17, 5, 16, 27,
    -- filter=37 channel=14
    81, 32, 144, -13, -303, -275, -118, -98, -86,
    -- filter=37 channel=15
    -65, -127, -233, 23, -30, -3, -46, -52, 72,
    -- filter=37 channel=16
    -71, -122, 70, 4, -21, -214, 198, -36, -75,
    -- filter=37 channel=17
    -107, 177, 63, -197, 85, 9, -97, 62, -51,
    -- filter=37 channel=18
    4, 57, -79, 55, -139, 109, -260, -110, 172,
    -- filter=37 channel=19
    66, 88, -82, -185, -117, 53, -346, 246, -185,
    -- filter=37 channel=20
    -94, -4, 86, 106, 200, 11, -124, -152, 38,
    -- filter=37 channel=21
    -234, 17, -112, 100, -55, 55, 157, 197, -111,
    -- filter=37 channel=22
    274, -67, 9, 128, 65, 68, -139, -6, 42,
    -- filter=37 channel=23
    50, 85, 69, 56, 52, -44, -39, -154, -58,
    -- filter=37 channel=24
    134, -103, -56, -148, 200, -29, 91, 69, 79,
    -- filter=37 channel=25
    116, -128, 95, 95, -133, -47, -134, -176, -188,
    -- filter=37 channel=26
    92, -12, 67, 119, 27, 68, 57, 20, -83,
    -- filter=37 channel=27
    136, -63, 32, 59, 105, -82, -2, -56, 7,
    -- filter=37 channel=28
    70, 189, -132, -19, -146, -249, -64, 7, 87,
    -- filter=37 channel=29
    122, -64, 77, -128, -269, 42, 33, -157, 64,
    -- filter=37 channel=30
    -154, 225, 16, 40, -75, 12, 28, -5, -7,
    -- filter=37 channel=31
    -28, -72, -49, 226, -34, 145, -65, -70, 86,
    -- filter=38 channel=0
    -27, -200, -99, -14, 90, 174, 72, -31, 97,
    -- filter=38 channel=1
    -246, -391, 258, 83, -7, -458, -138, 139, 267,
    -- filter=38 channel=2
    -61, 146, 55, 8, 52, -61, -154, 254, 92,
    -- filter=38 channel=3
    -220, -199, 93, -65, 133, -48, 100, 46, 112,
    -- filter=38 channel=4
    75, -159, 2, -172, 146, -412, -269, -153, 70,
    -- filter=38 channel=5
    -112, 186, -36, -28, -61, -125, -19, -15, -19,
    -- filter=38 channel=6
    -9, -103, -420, -57, -83, -458, -24, -72, 84,
    -- filter=38 channel=7
    -111, -18, 51, -119, 81, -118, -4, 64, 139,
    -- filter=38 channel=8
    -44, -94, -30, -77, -161, -264, 82, 132, 1,
    -- filter=38 channel=9
    99, 42, -60, 83, 87, 24, -57, -90, 75,
    -- filter=38 channel=10
    17, 108, -251, -64, -78, -332, -74, -225, 8,
    -- filter=38 channel=11
    11, 80, 15, 130, 23, -7, 10, 13, -201,
    -- filter=38 channel=12
    107, 38, -105, 140, -106, -58, -146, 96, -122,
    -- filter=38 channel=13
    -4, 0, -1, -8, -14, 1, 11, -10, -9,
    -- filter=38 channel=14
    -114, 76, -148, -65, 85, 70, 61, 79, -13,
    -- filter=38 channel=15
    130, -133, 137, -105, -141, 70, -163, 20, 150,
    -- filter=38 channel=16
    -22, 48, -33, -69, -361, -22, -83, 269, -9,
    -- filter=38 channel=17
    83, 88, 111, 36, -49, -9, 37, 76, 186,
    -- filter=38 channel=18
    -163, -372, 117, -3, 24, 105, 182, -65, 26,
    -- filter=38 channel=19
    114, -65, -101, 199, 71, 7, 40, -183, 50,
    -- filter=38 channel=20
    -58, 241, -33, 30, -289, 87, -100, 66, -149,
    -- filter=38 channel=21
    51, 47, -37, -138, 41, 26, 3, -135, 133,
    -- filter=38 channel=22
    151, -168, -33, 158, -97, 223, 147, -407, 53,
    -- filter=38 channel=23
    -171, 6, -206, -172, 8, 23, -212, -62, -3,
    -- filter=38 channel=24
    25, -45, 133, 45, -63, -72, 143, 76, -260,
    -- filter=38 channel=25
    27, 20, 209, -66, 6, 20, 69, -52, -360,
    -- filter=38 channel=26
    195, -61, 38, -213, 84, 193, -149, -68, 31,
    -- filter=38 channel=27
    -73, 15, 17, -12, -307, 33, 67, -99, 59,
    -- filter=38 channel=28
    -23, -89, -200, 78, -28, 119, 192, 99, -48,
    -- filter=38 channel=29
    -268, -33, -88, 60, 45, -76, 94, -36, 62,
    -- filter=38 channel=30
    179, 98, 35, -7, -282, -94, 4, 121, -228,
    -- filter=38 channel=31
    83, -282, 119, 45, 179, 30, -105, -35, -102,
    -- filter=39 channel=0
    9, -223, 19, -6, 40, 36, -34, 71, 6,
    -- filter=39 channel=1
    10, 86, -148, 63, -79, 190, -133, 160, 173,
    -- filter=39 channel=2
    -112, -49, -1, 10, -36, -97, 287, 3, -123,
    -- filter=39 channel=3
    -49, -46, 9, -77, -37, 66, -74, 114, -89,
    -- filter=39 channel=4
    -39, -70, -4, -61, -34, 14, 52, -69, -61,
    -- filter=39 channel=5
    -294, 34, 7, -143, -26, 116, 116, -216, -331,
    -- filter=39 channel=6
    86, -52, 100, -55, -248, 52, -181, -158, 65,
    -- filter=39 channel=7
    -87, -239, -17, 98, -51, -147, 136, 215, -51,
    -- filter=39 channel=8
    -103, -56, -89, -13, -131, 54, 67, 19, 156,
    -- filter=39 channel=9
    128, 191, -64, -14, -68, -70, 94, -88, -40,
    -- filter=39 channel=10
    61, -20, 62, 54, 93, 33, 92, 80, -136,
    -- filter=39 channel=11
    -76, -309, -270, -44, 117, 179, 221, 123, 67,
    -- filter=39 channel=12
    -40, -114, -42, 126, 45, 47, 148, 58, 35,
    -- filter=39 channel=13
    -17, -3, -21, 12, -20, -13, 32, -14, -19,
    -- filter=39 channel=14
    55, 54, -48, 94, -58, 46, -29, 85, 75,
    -- filter=39 channel=15
    12, -117, -250, -63, 104, -17, 165, 214, 154,
    -- filter=39 channel=16
    -110, -50, -150, 57, -45, -146, -89, -190, -63,
    -- filter=39 channel=17
    -38, 8, -94, -118, 43, -11, -86, 117, 281,
    -- filter=39 channel=18
    -63, 78, -53, -274, -85, -312, -108, 123, -218,
    -- filter=39 channel=19
    60, -88, 16, -34, 117, -20, 47, 174, 48,
    -- filter=39 channel=20
    57, 52, -178, -82, 26, -126, 34, -48, 5,
    -- filter=39 channel=21
    36, 19, 135, -72, 104, 54, -95, -302, -65,
    -- filter=39 channel=22
    10, 211, 187, -75, -36, 232, -134, 103, -258,
    -- filter=39 channel=23
    -51, -33, 17, -220, -4, -91, 116, 5, -1,
    -- filter=39 channel=24
    61, -210, -111, 41, 29, -92, -114, 16, 97,
    -- filter=39 channel=25
    271, 33, -162, -52, 56, -800, -296, 180, -86,
    -- filter=39 channel=26
    21, -347, -154, -90, 60, -195, 19, -149, -47,
    -- filter=39 channel=27
    26, -71, 14, 101, -210, -81, -8, -53, -40,
    -- filter=39 channel=28
    -21, 64, 225, -24, 19, 108, 14, -80, -116,
    -- filter=39 channel=29
    69, -160, -91, 49, -97, -56, 45, 68, 186,
    -- filter=39 channel=30
    -18, -207, 85, 17, 41, -70, 22, -71, -109,
    -- filter=39 channel=31
    -57, 144, 212, -49, -170, -181, -8, 140, -145,
    -- filter=40 channel=0
    54, -68, -96, 94, -142, -93, 139, -97, -9,
    -- filter=40 channel=1
    126, -35, -78, 110, -244, -48, 101, -175, 122,
    -- filter=40 channel=2
    73, -131, 259, 54, -7, -8, -171, -113, -55,
    -- filter=40 channel=3
    -70, 45, -287, -155, 18, -24, -105, 24, -33,
    -- filter=40 channel=4
    -120, -50, -103, -216, -269, 79, -124, -40, -136,
    -- filter=40 channel=5
    125, 3, -69, 49, -58, -97, 3, 25, -82,
    -- filter=40 channel=6
    65, -9, -123, 60, -39, 52, 72, -34, 26,
    -- filter=40 channel=7
    -45, -80, -57, -206, -30, -33, -125, 74, 84,
    -- filter=40 channel=8
    29, 43, -31, 26, -53, -16, 53, 29, 117,
    -- filter=40 channel=9
    27, -193, -9, -65, -295, -282, -51, -52, -207,
    -- filter=40 channel=10
    123, 0, -62, 30, 56, -92, -58, -82, 0,
    -- filter=40 channel=11
    -8, 114, 20, 6, 132, 202, 111, -66, 128,
    -- filter=40 channel=12
    -17, -39, -5, -364, -156, -198, -174, -88, 39,
    -- filter=40 channel=13
    8, -3, 0, -5, -20, 11, -8, 7, -19,
    -- filter=40 channel=14
    46, -120, 65, 77, -147, -24, 41, 53, -98,
    -- filter=40 channel=15
    -93, 61, -60, -54, -54, 144, 33, -199, -172,
    -- filter=40 channel=16
    -99, 52, 1, -165, -72, 55, -156, -121, -136,
    -- filter=40 channel=17
    -130, -194, 47, 33, -347, 68, -50, -357, 103,
    -- filter=40 channel=18
    -22, 118, -184, -180, -7, -238, -110, -16, 53,
    -- filter=40 channel=19
    98, -53, -170, 5, 12, 65, -117, -162, 20,
    -- filter=40 channel=20
    62, 105, -48, -106, -75, 93, -55, 19, 52,
    -- filter=40 channel=21
    56, 104, 55, -60, -68, 280, -94, -54, 38,
    -- filter=40 channel=22
    -68, -172, -113, 63, 17, 97, 12, 14, -101,
    -- filter=40 channel=23
    -8, -56, -14, -75, 96, -19, 83, 181, 75,
    -- filter=40 channel=24
    -83, -62, -60, -166, 148, 59, 28, 102, 131,
    -- filter=40 channel=25
    33, 34, -89, -246, 9, -75, 139, -84, 47,
    -- filter=40 channel=26
    30, 44, -44, -46, 5, -119, 107, 138, 72,
    -- filter=40 channel=27
    -39, -16, -11, -25, -242, -50, 24, -149, -186,
    -- filter=40 channel=28
    -138, -3, 24, -126, 13, 75, 34, -82, 57,
    -- filter=40 channel=29
    10, 6, -10, -110, -64, 1, 26, 66, -54,
    -- filter=40 channel=30
    -81, 11, -137, -71, 16, -8, 29, -73, 37,
    -- filter=40 channel=31
    -161, 9, -74, -140, 143, -61, 58, 123, 191,
    -- filter=41 channel=0
    73, -139, -54, 33, 154, -88, 73, -25, 31,
    -- filter=41 channel=1
    -157, -65, -73, -113, -224, -23, -41, -73, -25,
    -- filter=41 channel=2
    25, -31, -84, 174, 91, -216, 54, 142, -192,
    -- filter=41 channel=3
    119, -128, 45, -2, 142, -9, -145, -77, -158,
    -- filter=41 channel=4
    -134, 173, 83, 5, 126, 96, -137, -13, -101,
    -- filter=41 channel=5
    105, 35, 34, 102, 65, 216, -2, 42, 131,
    -- filter=41 channel=6
    -68, 85, 92, -44, -125, 171, -140, -19, 33,
    -- filter=41 channel=7
    -133, -101, -59, -189, -145, 17, -269, -55, 111,
    -- filter=41 channel=8
    63, -17, 27, 54, 25, -14, -100, 116, -88,
    -- filter=41 channel=9
    122, 189, 10, -21, -181, 197, -312, -46, -95,
    -- filter=41 channel=10
    -15, -186, 170, 182, 67, -94, 129, -85, 82,
    -- filter=41 channel=11
    -2, 191, -88, 174, -183, -92, -53, 71, -27,
    -- filter=41 channel=12
    149, -130, -80, 149, 179, 198, 25, 69, 256,
    -- filter=41 channel=13
    23, -8, 13, -28, -12, -4, -16, 16, -9,
    -- filter=41 channel=14
    -116, -68, -8, -2, -83, 31, -80, -35, -8,
    -- filter=41 channel=15
    0, -43, -128, 200, -7, -167, 97, -59, 39,
    -- filter=41 channel=16
    39, 116, -20, -69, -206, 149, 29, 56, 17,
    -- filter=41 channel=17
    185, 137, 65, 8, -135, 83, -511, -21, 256,
    -- filter=41 channel=18
    -51, -197, 95, 28, 18, -213, 113, 3, -78,
    -- filter=41 channel=19
    -87, 57, -79, 136, -96, 25, -46, 32, -57,
    -- filter=41 channel=20
    16, -178, 3, 142, -120, 10, 46, -77, -125,
    -- filter=41 channel=21
    27, -92, 149, -133, 57, -27, 27, -272, -70,
    -- filter=41 channel=22
    -81, -145, 119, -75, 63, 19, -108, -43, -97,
    -- filter=41 channel=23
    27, 26, 121, -72, -100, 49, -181, -223, 177,
    -- filter=41 channel=24
    48, 34, 3, -134, 256, -89, 62, 75, -24,
    -- filter=41 channel=25
    -151, 13, -75, 53, 182, 24, -39, 23, 122,
    -- filter=41 channel=26
    52, -1, -41, -8, 35, 0, -46, -62, 97,
    -- filter=41 channel=27
    -88, 53, 142, -210, 0, 169, -139, 141, 12,
    -- filter=41 channel=28
    133, -48, -43, 64, -11, -71, -102, 254, -50,
    -- filter=41 channel=29
    -98, 0, 106, -28, -143, 15, 151, 91, 11,
    -- filter=41 channel=30
    70, -124, -47, -252, 158, 132, -159, 179, -86,
    -- filter=41 channel=31
    -55, -70, -132, 157, -121, -26, 70, 24, -60,
    -- filter=42 channel=0
    -114, -26, -55, 86, -184, -245, 27, 45, 61,
    -- filter=42 channel=1
    -65, 126, -12, -43, -227, 41, 128, -173, -303,
    -- filter=42 channel=2
    -11, -7, -23, -60, 51, 71, -106, 203, -89,
    -- filter=42 channel=3
    -73, 250, 202, 2, -83, 46, -169, 31, -227,
    -- filter=42 channel=4
    -71, -30, 137, -37, 26, -61, 42, 129, 75,
    -- filter=42 channel=5
    34, -65, -73, 48, -118, -199, -46, -64, -139,
    -- filter=42 channel=6
    178, -15, -263, 205, -347, -9, -141, -18, -188,
    -- filter=42 channel=7
    56, 132, -6, 84, -19, -27, 154, 49, -154,
    -- filter=42 channel=8
    34, 13, -122, 51, -365, -56, -48, -178, -89,
    -- filter=42 channel=9
    39, -58, 36, -17, 70, -136, 95, 83, 211,
    -- filter=42 channel=10
    -83, 13, -44, 91, -218, -224, 99, -61, -69,
    -- filter=42 channel=11
    14, -32, 126, 70, -4, 200, 18, 97, 47,
    -- filter=42 channel=12
    -118, 89, -93, -33, 39, 182, 5, 189, 115,
    -- filter=42 channel=13
    -7, -7, 3, 1, -4, 19, 24, 2, -16,
    -- filter=42 channel=14
    63, -36, 125, 98, 30, -44, 50, 4, 27,
    -- filter=42 channel=15
    -219, -77, -7, -87, 26, 56, -145, 35, 148,
    -- filter=42 channel=16
    45, 203, 154, 7, 102, -31, 4, 25, 20,
    -- filter=42 channel=17
    58, 10, -7, 0, 280, -58, -68, 36, -59,
    -- filter=42 channel=18
    -7, 99, -69, -80, -5, -86, -116, -169, -21,
    -- filter=42 channel=19
    64, 12, -119, 123, -126, -213, -143, 15, -129,
    -- filter=42 channel=20
    -149, -68, 147, 249, -110, -211, 49, -63, -106,
    -- filter=42 channel=21
    121, -149, 52, 92, -72, 109, -54, 213, 106,
    -- filter=42 channel=22
    68, -8, 4, -11, -90, -14, 51, 112, -106,
    -- filter=42 channel=23
    112, -98, 91, 73, 51, -94, -162, 54, 113,
    -- filter=42 channel=24
    -170, -5, 61, 97, -153, 27, 106, -50, -86,
    -- filter=42 channel=25
    -113, -9, 22, -87, 168, 122, -171, -22, 261,
    -- filter=42 channel=26
    138, 97, 69, -64, -25, 26, -137, -127, 14,
    -- filter=42 channel=27
    138, 33, 56, 7, 8, 33, 171, -54, 177,
    -- filter=42 channel=28
    46, 0, -102, 24, 52, -46, 27, -66, -46,
    -- filter=42 channel=29
    89, -118, 14, -127, 29, 71, -188, -167, 203,
    -- filter=42 channel=30
    -46, 184, 126, -41, 10, -20, 6, -108, -139,
    -- filter=42 channel=31
    -52, 10, -39, -27, -124, 50, -117, 158, 35,
    -- filter=43 channel=0
    69, -332, 94, -111, -268, 52, -17, -60, 29,
    -- filter=43 channel=1
    -50, 81, -161, -9, -140, -75, -21, -30, 56,
    -- filter=43 channel=2
    30, -83, 3, -68, 80, 35, -111, 280, -207,
    -- filter=43 channel=3
    177, -43, 49, -91, 6, -145, -67, -54, -277,
    -- filter=43 channel=4
    -102, -66, 137, -45, -639, -47, -23, -61, -61,
    -- filter=43 channel=5
    82, -116, -114, -52, 76, -202, 117, 131, -31,
    -- filter=43 channel=6
    145, 164, -242, 42, 180, -118, 39, 30, 27,
    -- filter=43 channel=7
    59, 87, 41, 129, 130, 155, -34, -77, 52,
    -- filter=43 channel=8
    -150, 33, -137, 40, -50, 146, 59, -97, 133,
    -- filter=43 channel=9
    -73, -5, 141, -12, -190, -106, 114, -78, -201,
    -- filter=43 channel=10
    -12, 135, -81, 99, -32, -52, 88, -44, 108,
    -- filter=43 channel=11
    -58, -250, 11, 117, 77, 124, 68, 45, 12,
    -- filter=43 channel=12
    -27, 39, 97, 87, 94, 133, -92, 10, -138,
    -- filter=43 channel=13
    8, -12, 7, 1, -1, 10, 17, -6, -8,
    -- filter=43 channel=14
    -250, -269, -49, -248, -142, -94, 55, 14, 122,
    -- filter=43 channel=15
    93, 31, 90, -103, 16, 151, -281, -28, -185,
    -- filter=43 channel=16
    106, 73, 7, -13, 130, -23, 99, -48, -210,
    -- filter=43 channel=17
    210, -148, 81, -3, 17, 37, -15, 49, -17,
    -- filter=43 channel=18
    -161, 9, -5, 135, 72, -63, -246, 49, -19,
    -- filter=43 channel=19
    166, -133, 116, 35, -284, 224, -12, -120, 8,
    -- filter=43 channel=20
    -20, 146, 74, -48, -122, 13, -132, 65, -7,
    -- filter=43 channel=21
    68, -113, 54, 75, -262, -59, 146, -85, 125,
    -- filter=43 channel=22
    80, 126, -89, -25, -50, 22, 43, 0, 232,
    -- filter=43 channel=23
    89, -183, -182, -46, -76, -198, 34, 47, 39,
    -- filter=43 channel=24
    -62, 24, 150, 180, 29, -55, 80, -39, -200,
    -- filter=43 channel=25
    -42, 51, 191, -140, -58, 53, 38, 26, -13,
    -- filter=43 channel=26
    -37, 111, 134, -85, -11, 31, -119, 170, -71,
    -- filter=43 channel=27
    -321, -145, -134, -75, -131, -170, -47, -174, -124,
    -- filter=43 channel=28
    56, -79, -21, 62, 33, 5, -188, -103, -103,
    -- filter=43 channel=29
    -48, 107, -171, -111, 103, 36, -60, 66, 221,
    -- filter=43 channel=30
    113, -64, 109, 37, -99, 72, -47, -74, -37,
    -- filter=43 channel=31
    -191, 7, 121, -24, 70, 86, 17, 172, -6,
    -- filter=44 channel=0
    9, 96, -21, 2, 62, 47, -62, 48, 103,
    -- filter=44 channel=1
    117, 67, -35, 245, -87, 72, 13, 32, -15,
    -- filter=44 channel=2
    65, -29, 36, 224, -100, 3, 57, -246, -244,
    -- filter=44 channel=3
    52, -98, -8, 13, -90, -139, 11, -234, 44,
    -- filter=44 channel=4
    48, 109, 37, -58, 11, -9, 92, 66, -94,
    -- filter=44 channel=5
    -39, 15, 52, -39, 75, -37, -14, -61, -46,
    -- filter=44 channel=6
    -7, 47, 108, -189, -22, -18, -197, -205, -18,
    -- filter=44 channel=7
    112, 136, -11, -25, -70, 189, -84, -15, 58,
    -- filter=44 channel=8
    -109, -23, 0, -17, -155, 44, 64, 81, -3,
    -- filter=44 channel=9
    162, 116, 48, -351, 73, 53, -95, 27, 6,
    -- filter=44 channel=10
    22, 44, 25, 11, 75, -50, -43, -76, -69,
    -- filter=44 channel=11
    199, -210, 53, -68, -93, 52, -34, -11, -8,
    -- filter=44 channel=12
    12, 156, -150, 41, 134, -153, 126, -94, -10,
    -- filter=44 channel=13
    2, 25, 18, 8, 14, 1, -4, -15, 1,
    -- filter=44 channel=14
    -8, 13, -44, -58, -108, 18, -37, 38, -143,
    -- filter=44 channel=15
    148, -67, -194, 125, -85, 160, 28, -6, -16,
    -- filter=44 channel=16
    72, 70, -74, 61, 2, -13, 102, 139, -88,
    -- filter=44 channel=17
    -374, 201, -138, 56, -229, 209, 3, 179, -42,
    -- filter=44 channel=18
    -104, -114, -22, -72, -254, 114, 52, -132, -21,
    -- filter=44 channel=19
    235, -23, -279, 197, -80, 69, 51, -43, -4,
    -- filter=44 channel=20
    229, 124, -199, 205, -2, -223, 108, -137, 4,
    -- filter=44 channel=21
    -208, 25, -54, 166, -68, 117, 21, -166, 39,
    -- filter=44 channel=22
    -95, -29, 113, -12, 142, 38, -21, 105, 83,
    -- filter=44 channel=23
    122, -96, -133, -68, -170, -16, -8, -121, -115,
    -- filter=44 channel=24
    271, 34, 17, 8, 114, -153, -75, -7, -248,
    -- filter=44 channel=25
    66, -88, -101, -5, -157, 160, 40, -39, -137,
    -- filter=44 channel=26
    8, -140, -126, 37, 170, -301, 121, 7, 21,
    -- filter=44 channel=27
    -101, 156, 38, -15, -27, 3, -1, -25, -40,
    -- filter=44 channel=28
    -44, 222, 81, 52, -37, -85, -75, -124, -57,
    -- filter=44 channel=29
    -56, -188, 51, 212, -56, -69, 248, 126, 26,
    -- filter=44 channel=30
    -26, 82, 6, -178, 94, -43, 26, 137, -56,
    -- filter=44 channel=31
    -13, 69, 200, -96, 51, -2, -5, 160, 18,
    -- filter=45 channel=0
    54, 8, -139, -46, 61, -83, 75, 91, 30,
    -- filter=45 channel=1
    -85, -62, 138, 23, -22, -83, 61, 90, 11,
    -- filter=45 channel=2
    -18, -4, -161, 21, 62, -193, 238, 113, 11,
    -- filter=45 channel=3
    -66, 23, -91, -41, -61, -52, 34, -66, 188,
    -- filter=45 channel=4
    -128, -114, 53, -43, -29, 105, -126, 165, -46,
    -- filter=45 channel=5
    25, -22, -118, 96, 146, 75, 72, -66, -26,
    -- filter=45 channel=6
    -204, -159, 174, -177, -83, 83, -98, 61, 70,
    -- filter=45 channel=7
    92, -23, 5, 79, -28, -35, 215, -4, -18,
    -- filter=45 channel=8
    44, 3, -26, -55, -95, 66, -32, -52, 28,
    -- filter=45 channel=9
    -12, -174, 44, -31, -46, 108, -99, 3, 19,
    -- filter=45 channel=10
    122, 31, -5, -72, -154, -109, -8, -128, 15,
    -- filter=45 channel=11
    30, -37, -28, -143, 96, 80, 21, 87, -10,
    -- filter=45 channel=12
    -25, -64, 209, 231, 189, 28, 221, -46, -40,
    -- filter=45 channel=13
    19, 27, -3, -15, 14, -18, -4, 8, 5,
    -- filter=45 channel=14
    -7, -70, -83, 87, -35, -119, -92, 178, 141,
    -- filter=45 channel=15
    45, -24, 62, 59, -228, -128, -9, 16, -75,
    -- filter=45 channel=16
    120, 70, 129, 38, 100, 89, -62, -105, 49,
    -- filter=45 channel=17
    259, 58, -182, 111, 236, -256, -44, 118, 146,
    -- filter=45 channel=18
    -115, 130, -132, 142, 134, -11, 12, 61, -125,
    -- filter=45 channel=19
    43, -36, 97, -233, -167, -75, -109, -46, -270,
    -- filter=45 channel=20
    -50, -92, 219, -82, 77, -50, -120, -26, 52,
    -- filter=45 channel=21
    -225, 161, 211, -57, 24, -42, 30, -8, -109,
    -- filter=45 channel=22
    -113, 102, 75, 184, 89, 1, 101, -127, -23,
    -- filter=45 channel=23
    60, 81, -24, -1, -53, -72, -72, 57, -59,
    -- filter=45 channel=24
    146, -77, 152, -314, -25, -39, -18, -5, -161,
    -- filter=45 channel=25
    22, -115, 111, 27, -27, -98, -9, 71, 6,
    -- filter=45 channel=26
    -75, -94, -168, 9, -240, -27, 254, -32, -239,
    -- filter=45 channel=27
    -56, -105, -83, 13, 175, 114, -1, 40, -99,
    -- filter=45 channel=28
    -56, 33, 95, -160, 181, 120, -236, -66, 99,
    -- filter=45 channel=29
    -111, -6, -32, -375, -187, 4, -97, -159, -187,
    -- filter=45 channel=30
    -174, 46, 9, 133, 186, -170, -259, -55, 92,
    -- filter=45 channel=31
    -13, 184, 67, -105, 140, 126, -108, 52, -10,
    -- filter=46 channel=0
    -268, 30, -55, 66, 12, -16, -38, -17, 36,
    -- filter=46 channel=1
    -3, -286, -76, 102, -317, -124, 57, -187, 109,
    -- filter=46 channel=2
    33, -135, 16, -244, 21, 42, -249, 23, 169,
    -- filter=46 channel=3
    -3, -110, 45, 109, 128, 48, 39, -66, -4,
    -- filter=46 channel=4
    -1, 20, 84, 112, 37, 120, -67, 153, 120,
    -- filter=46 channel=5
    -198, -119, -128, 21, 30, -116, 44, -324, -96,
    -- filter=46 channel=6
    65, 47, 124, 35, -33, -132, -142, 66, -79,
    -- filter=46 channel=7
    -81, -72, -70, -355, -94, -119, -187, -152, -35,
    -- filter=46 channel=8
    -153, -196, 66, -96, -148, 70, 217, -95, -66,
    -- filter=46 channel=9
    -99, 84, -19, 187, 105, 10, 105, 215, 241,
    -- filter=46 channel=10
    -28, 104, -17, -162, 0, 21, -37, -104, -33,
    -- filter=46 channel=11
    -111, -37, -8, -51, 127, -13, -111, -208, 55,
    -- filter=46 channel=12
    97, 18, -16, 88, 89, -206, 173, -51, -43,
    -- filter=46 channel=13
    -10, 18, -21, 1, -1, 0, -8, 10, -17,
    -- filter=46 channel=14
    -159, 13, -66, -52, 62, 84, 159, 227, 140,
    -- filter=46 channel=15
    50, -111, 78, -6, 184, 37, 93, -41, 47,
    -- filter=46 channel=16
    -12, 28, 9, 54, -83, 0, -102, -14, -80,
    -- filter=46 channel=17
    -73, 136, -158, -210, 161, -784, 21, 241, 114,
    -- filter=46 channel=18
    18, 142, 9, 0, -87, 65, -21, -74, -99,
    -- filter=46 channel=19
    -11, -2, 35, 6, -152, 57, -157, 136, -23,
    -- filter=46 channel=20
    -74, -176, 195, 84, 65, -98, 17, -167, 165,
    -- filter=46 channel=21
    48, 30, -26, -12, -98, 26, 139, 52, -6,
    -- filter=46 channel=22
    149, 145, -132, 92, 97, -22, 23, 37, -58,
    -- filter=46 channel=23
    206, -88, -273, 84, -46, -72, 30, 271, 34,
    -- filter=46 channel=24
    198, 41, 36, 136, -14, -222, -82, -78, 4,
    -- filter=46 channel=25
    18, -18, -51, 36, -80, 60, 93, 18, -8,
    -- filter=46 channel=26
    137, -25, -57, 261, -148, -53, -125, -61, 51,
    -- filter=46 channel=27
    -113, -17, 43, -34, -304, -80, 95, 61, -63,
    -- filter=46 channel=28
    98, -50, 145, -259, 87, 0, 84, 243, 239,
    -- filter=46 channel=29
    -105, -90, -5, -360, -217, 30, -37, -186, -177,
    -- filter=46 channel=30
    -135, -93, 194, -17, 17, -151, 35, -94, 125,
    -- filter=46 channel=31
    1, -56, 13, 80, -82, 20, 31, -43, -82,
    -- filter=47 channel=0
    35, -164, -101, 87, -178, -180, 121, -66, -90,
    -- filter=47 channel=1
    14, 144, -58, 247, 59, 107, -173, 56, 62,
    -- filter=47 channel=2
    255, 206, -113, -217, -23, -79, 46, 205, -179,
    -- filter=47 channel=3
    42, 161, -181, 74, -508, -76, -145, -105, -345,
    -- filter=47 channel=4
    25, 25, 9, 258, 275, -2, 29, 35, 23,
    -- filter=47 channel=5
    108, -100, -7, 0, 46, 37, 29, -173, -216,
    -- filter=47 channel=6
    -7, -62, -168, -58, -98, 101, 86, -243, 15,
    -- filter=47 channel=7
    105, 161, -650, 111, -30, -53, 168, 78, 80,
    -- filter=47 channel=8
    42, 30, -132, -13, 17, -102, 15, -47, 150,
    -- filter=47 channel=9
    33, -183, 6, 55, 19, -9, 223, 396, -58,
    -- filter=47 channel=10
    -17, 97, 30, -396, -64, -80, 134, 69, 136,
    -- filter=47 channel=11
    -159, 235, -82, 32, 76, -67, -36, 54, 23,
    -- filter=47 channel=12
    -107, -6, 18, -121, 233, 15, -375, -117, 172,
    -- filter=47 channel=13
    7, -12, -11, -7, -5, -8, -9, -3, -8,
    -- filter=47 channel=14
    51, 8, -69, 25, 103, -167, 58, 67, -128,
    -- filter=47 channel=15
    -17, -248, -70, -310, 120, -56, -150, 9, 65,
    -- filter=47 channel=16
    -160, -17, -377, -110, -109, 120, 166, -175, 176,
    -- filter=47 channel=17
    -118, -188, -121, -173, 245, 9, 107, -246, 7,
    -- filter=47 channel=18
    61, 75, -337, -647, -190, 10, -471, -178, 225,
    -- filter=47 channel=19
    26, 74, 28, 20, -64, -137, 22, 54, -71,
    -- filter=47 channel=20
    -49, 53, 58, 123, 33, 215, -152, -264, 26,
    -- filter=47 channel=21
    -260, 271, 58, 129, 52, 60, -145, 148, 172,
    -- filter=47 channel=22
    -90, -54, -62, -300, -212, 85, 45, -596, -30,
    -- filter=47 channel=23
    -185, 98, -11, -50, 140, 59, 13, 112, -137,
    -- filter=47 channel=24
    -72, -112, -61, -104, -199, 159, 60, -262, -196,
    -- filter=47 channel=25
    -86, 61, 140, -198, -298, 190, -101, 212, 106,
    -- filter=47 channel=26
    61, 51, 168, -171, -115, -167, 152, -79, -298,
    -- filter=47 channel=27
    -197, -306, 54, -87, -293, 209, 23, -43, 110,
    -- filter=47 channel=28
    -49, 47, -51, -50, 73, 21, 38, -269, -77,
    -- filter=47 channel=29
    -121, -92, -132, -62, 241, -99, -78, 126, 106,
    -- filter=47 channel=30
    23, 75, -185, 115, -270, 94, 34, -5, 38,
    -- filter=47 channel=31
    -107, 137, -167, 281, -82, -367, -131, -5, -16,
    -- filter=48 channel=0
    80, -211, -75, 95, -178, -139, 2, 75, -125,
    -- filter=48 channel=1
    -44, -172, 87, -21, -211, -6, -54, -27, 9,
    -- filter=48 channel=2
    -241, 37, 252, -212, 185, 38, -38, -177, 149,
    -- filter=48 channel=3
    77, 209, 93, -23, -89, 19, -94, -1, -99,
    -- filter=48 channel=4
    -153, -21, -190, -26, 28, -237, 175, 155, -58,
    -- filter=48 channel=5
    -40, -74, 107, -309, 41, 121, -18, -77, -114,
    -- filter=48 channel=6
    -97, 25, 59, -9, -24, 125, -121, 0, 121,
    -- filter=48 channel=7
    53, -165, -101, -21, -107, 122, -24, -76, 79,
    -- filter=48 channel=8
    3, 23, 72, -91, 0, 109, -29, -100, 0,
    -- filter=48 channel=9
    -22, 193, 55, 26, -12, -19, 94, -132, -82,
    -- filter=48 channel=10
    79, -7, -126, -79, 4, -45, -4, 40, -33,
    -- filter=48 channel=11
    -501, -112, 308, -86, -74, 263, -21, -147, 311,
    -- filter=48 channel=12
    -14, 170, -120, -42, -42, 46, -57, -99, 149,
    -- filter=48 channel=13
    1, 19, 3, 5, -3, -14, -25, -6, 0,
    -- filter=48 channel=14
    -30, -39, 63, 161, 316, -78, 38, 23, -450,
    -- filter=48 channel=15
    -64, 182, -59, 18, 54, 125, -97, -150, -26,
    -- filter=48 channel=16
    -100, -95, 60, -145, 139, -53, -138, 79, -256,
    -- filter=48 channel=17
    -105, 125, 47, -56, -181, 127, -292, -117, -168,
    -- filter=48 channel=18
    142, 8, -167, 35, -220, -274, -50, -4, 66,
    -- filter=48 channel=19
    66, 205, -77, 28, 32, -47, 38, -100, 105,
    -- filter=48 channel=20
    -11, -142, 70, -82, -49, 150, 24, -42, -89,
    -- filter=48 channel=21
    42, -26, 203, -158, 107, -61, -96, 83, -123,
    -- filter=48 channel=22
    42, -33, -28, 191, 42, -67, -66, -48, 91,
    -- filter=48 channel=23
    -34, -216, 156, -111, 74, -109, 22, 159, 35,
    -- filter=48 channel=24
    -48, 61, -71, 79, 112, -294, 100, 34, 65,
    -- filter=48 channel=25
    175, 69, -89, 11, -110, 63, 148, 71, -36,
    -- filter=48 channel=26
    -74, 27, 139, 56, 42, 78, -70, 36, 42,
    -- filter=48 channel=27
    40, 210, -101, -80, 71, -112, -30, 35, -196,
    -- filter=48 channel=28
    13, 256, -144, -12, 135, -323, -51, 3, -182,
    -- filter=48 channel=29
    -80, 70, -27, 61, 136, -103, 53, 95, -46,
    -- filter=48 channel=30
    87, -239, 83, 39, 35, -20, -34, -5, 21,
    -- filter=48 channel=31
    -58, 7, -60, -53, -9, -181, 87, 54, 83,
    -- filter=49 channel=0
    30, 87, 168, 179, 134, 236, -93, 118, 96,
    -- filter=49 channel=1
    -24, -28, -101, 34, 218, -81, 33, 28, -193,
    -- filter=49 channel=2
    102, -41, -12, -187, 137, 170, 30, -180, 84,
    -- filter=49 channel=3
    -308, -62, 123, -161, -12, -122, 158, -103, -110,
    -- filter=49 channel=4
    102, 83, -71, 54, -74, -53, -157, -89, 69,
    -- filter=49 channel=5
    19, 74, -21, 103, -73, -2, 27, 114, -12,
    -- filter=49 channel=6
    -114, 5, 61, -103, -11, -156, 95, 57, 58,
    -- filter=49 channel=7
    24, 104, 53, -259, 98, -28, 36, 4, -61,
    -- filter=49 channel=8
    14, 119, -25, 123, -47, -37, 0, 11, -70,
    -- filter=49 channel=9
    -16, 3, -30, 90, -4, -171, -272, 34, 42,
    -- filter=49 channel=10
    -88, 41, -289, 16, 21, 107, -1, 70, 100,
    -- filter=49 channel=11
    -2, 2, -60, 198, 10, -167, 11, 6, 30,
    -- filter=49 channel=12
    -69, 32, -7, -14, 132, 51, -109, -69, -101,
    -- filter=49 channel=13
    -3, -6, -10, -23, 13, 2, -8, 23, -11,
    -- filter=49 channel=14
    -28, 69, 140, -159, -72, -54, -112, 35, 117,
    -- filter=49 channel=15
    43, -284, 72, 57, -111, -19, 86, -143, 25,
    -- filter=49 channel=16
    1, 101, 181, -63, 82, 124, 30, -6, 117,
    -- filter=49 channel=17
    -176, 103, 178, -269, 78, 84, 132, 105, -108,
    -- filter=49 channel=18
    -164, -27, -52, -74, 143, -56, -13, 11, 68,
    -- filter=49 channel=19
    -152, -62, -41, -279, -10, -10, -39, 100, 52,
    -- filter=49 channel=20
    59, 112, 110, -68, 229, -37, -68, -44, 107,
    -- filter=49 channel=21
    133, 23, -4, -13, 38, 181, 157, -311, -129,
    -- filter=49 channel=22
    -114, -156, 145, -312, 100, -307, -19, 134, -100,
    -- filter=49 channel=23
    57, -41, -37, 29, -74, -16, -56, 109, -299,
    -- filter=49 channel=24
    39, 77, -313, -2, -51, 103, 54, -4, -63,
    -- filter=49 channel=25
    -36, 37, -1, -64, -58, -177, 54, -78, 114,
    -- filter=49 channel=26
    -31, -149, 51, 87, 48, -100, 107, -14, -123,
    -- filter=49 channel=27
    61, 196, 113, -237, -47, -15, -140, -256, -230,
    -- filter=49 channel=28
    12, -125, 61, -57, 17, -38, -110, 32, 61,
    -- filter=49 channel=29
    -103, 67, 131, -98, 36, 36, 62, -184, 0,
    -- filter=49 channel=30
    -27, -197, -234, -79, 153, -59, 142, -129, -117,
    -- filter=49 channel=31
    -41, -120, 36, 30, 87, 142, 58, 73, 120,
    -- filter=50 channel=0
    83, 157, -33, 43, 92, 111, -22, -87, 88,
    -- filter=50 channel=1
    -84, 20, 152, 31, -52, 19, -70, -15, 209,
    -- filter=50 channel=2
    -289, 176, 21, 157, -80, 15, 51, 76, -117,
    -- filter=50 channel=3
    51, 17, -261, -103, -327, -111, -121, -25, -51,
    -- filter=50 channel=4
    51, 78, -37, 24, -2, -10, -68, -239, 4,
    -- filter=50 channel=5
    -207, -127, -83, 24, -2, 105, 113, -155, 144,
    -- filter=50 channel=6
    -88, -79, 60, 109, 5, -6, -46, 208, -105,
    -- filter=50 channel=7
    -94, 99, -297, 103, 48, -56, 73, 139, -22,
    -- filter=50 channel=8
    26, -9, 70, -23, 111, 37, -80, 4, 35,
    -- filter=50 channel=9
    80, 37, 45, -35, -40, -86, 39, -174, -88,
    -- filter=50 channel=10
    88, 23, -13, -179, -5, -102, 32, 21, 60,
    -- filter=50 channel=11
    134, 46, 84, -87, -137, -38, 84, 116, 61,
    -- filter=50 channel=12
    11, -249, -17, 13, -55, -143, 40, -11, -275,
    -- filter=50 channel=13
    2, 6, -9, -17, -8, 12, -2, 2, 5,
    -- filter=50 channel=14
    30, -49, 23, 88, 72, 68, -133, -67, 81,
    -- filter=50 channel=15
    158, 25, -163, -147, -147, 41, -42, -182, 85,
    -- filter=50 channel=16
    88, 7, 134, -112, -313, 91, -74, -207, -19,
    -- filter=50 channel=17
    120, 119, 7, 10, -21, -43, 113, -212, -164,
    -- filter=50 channel=18
    58, -106, -48, -78, 110, 154, -96, 268, -132,
    -- filter=50 channel=19
    17, 99, -128, -141, 234, -55, -49, -124, -35,
    -- filter=50 channel=20
    -6, -122, 97, -273, -42, -139, 254, -10, 42,
    -- filter=50 channel=21
    12, -120, 98, 0, 38, 94, 281, -276, -39,
    -- filter=50 channel=22
    46, 91, 23, 115, 4, 82, -54, -48, 34,
    -- filter=50 channel=23
    80, 61, -89, 59, 49, -106, 21, -59, 33,
    -- filter=50 channel=24
    -404, -99, -244, -436, -189, -277, 138, -320, -92,
    -- filter=50 channel=25
    -254, -77, -221, 124, -30, 86, 260, 194, 42,
    -- filter=50 channel=26
    -92, -6, 68, -169, -9, -3, 52, 4, 118,
    -- filter=50 channel=27
    97, -40, 64, 46, -23, -108, 57, -128, 4,
    -- filter=50 channel=28
    33, 61, 25, 120, 15, -177, 149, -18, -127,
    -- filter=50 channel=29
    -110, 35, -39, 12, -21, 37, 78, -147, -296,
    -- filter=50 channel=30
    -312, -3, -131, -4, -145, 8, 33, -35, 114,
    -- filter=50 channel=31
    32, -6, 208, -108, 16, -78, -298, 173, 31,
    -- filter=51 channel=0
    124, -29, -104, 111, -55, 118, -86, -76, 161,
    -- filter=51 channel=1
    -572, -349, 120, 53, 13, 12, 65, 97, 79,
    -- filter=51 channel=2
    24, 29, -48, -206, -138, 105, -26, 112, -22,
    -- filter=51 channel=3
    -98, 203, -91, -143, -63, 47, 125, -224, 37,
    -- filter=51 channel=4
    -213, -152, -324, 204, -17, -100, 197, -179, 19,
    -- filter=51 channel=5
    -47, -60, -15, 185, 145, -23, 125, 25, 65,
    -- filter=51 channel=6
    -265, 158, -4, 141, 11, -50, 90, 120, 25,
    -- filter=51 channel=7
    -209, 29, 133, -55, -35, -135, -154, 39, 94,
    -- filter=51 channel=8
    -190, 125, -67, -37, 90, 57, 78, -31, 83,
    -- filter=51 channel=9
    -147, -271, -119, -22, -50, -33, 113, 124, 18,
    -- filter=51 channel=10
    -103, -36, -85, -209, 67, 5, -123, -105, 179,
    -- filter=51 channel=11
    -60, -38, -43, 60, 38, -80, 117, -63, -18,
    -- filter=51 channel=12
    -81, -49, -118, -140, -152, -160, 29, 141, -25,
    -- filter=51 channel=13
    -3, -17, -13, 12, -11, -9, -14, 7, 0,
    -- filter=51 channel=14
    -35, 160, 119, 138, -102, 54, -160, -183, 51,
    -- filter=51 channel=15
    21, 98, -93, -171, 122, -72, 16, -91, 86,
    -- filter=51 channel=16
    63, 22, -15, -157, -103, 147, 35, -170, -58,
    -- filter=51 channel=17
    -87, -185, 15, -66, 231, 125, -25, -135, 123,
    -- filter=51 channel=18
    -168, 39, -79, -418, 110, 141, -148, 88, 202,
    -- filter=51 channel=19
    87, -45, -179, -36, 90, -113, -25, 8, -17,
    -- filter=51 channel=20
    -127, -226, 121, -204, 19, 157, 57, -49, 26,
    -- filter=51 channel=21
    -105, -673, -192, -226, -46, 151, -149, 108, 39,
    -- filter=51 channel=22
    -121, -133, 320, -111, 198, 126, -5, 98, 78,
    -- filter=51 channel=23
    136, -187, -101, 2, 16, -176, 65, 131, -49,
    -- filter=51 channel=24
    -58, 64, -44, -81, -23, 36, 239, 66, -64,
    -- filter=51 channel=25
    -164, -84, 115, -60, 72, -58, -18, 102, -16,
    -- filter=51 channel=26
    4, -18, -33, -46, 17, 130, -11, 170, -92,
    -- filter=51 channel=27
    38, -80, -109, -42, 10, -97, 57, 78, 72,
    -- filter=51 channel=28
    -99, -112, 85, -8, 205, -129, -96, -94, 62,
    -- filter=51 channel=29
    1, -56, -141, -122, 46, -8, 194, 30, 129,
    -- filter=51 channel=30
    19, -197, 148, 90, 9, -71, -169, -27, 31,
    -- filter=51 channel=31
    -38, -66, -13, -19, -91, 2, 15, 60, 137,
    -- filter=52 channel=0
    82, 70, 55, 24, 18, -42, -25, -8, 107,
    -- filter=52 channel=1
    83, 92, 149, 110, 23, 177, 112, -39, -239,
    -- filter=52 channel=2
    -94, 147, 60, -53, -6, 59, 61, -11, -36,
    -- filter=52 channel=3
    72, 27, -146, 18, 28, -153, 58, -32, 34,
    -- filter=52 channel=4
    -27, 122, 75, 135, 3, -168, -19, -148, -225,
    -- filter=52 channel=5
    122, 35, 25, 33, -69, -85, 58, -123, 109,
    -- filter=52 channel=6
    13, 74, 157, -48, 48, 13, 141, 94, 2,
    -- filter=52 channel=7
    -156, -7, -91, -84, -242, -264, -26, -143, -205,
    -- filter=52 channel=8
    -27, 65, -54, -64, 115, 109, -75, -114, -98,
    -- filter=52 channel=9
    -36, -36, 76, -168, -196, 1, -425, -161, -260,
    -- filter=52 channel=10
    60, -102, 7, 0, -97, -143, 224, -178, -6,
    -- filter=52 channel=11
    36, -82, 36, 58, -56, -86, 166, 132, 24,
    -- filter=52 channel=12
    -42, 18, -7, -211, -294, -138, -126, -298, -142,
    -- filter=52 channel=13
    15, 29, 12, 13, 8, 0, 18, -8, -13,
    -- filter=52 channel=14
    95, 2, 76, -4, -7, -32, 7, 146, 118,
    -- filter=52 channel=15
    248, 39, -6, -43, 153, -86, -111, -127, -1,
    -- filter=52 channel=16
    -84, -84, -202, -229, -116, 43, -226, -27, -4,
    -- filter=52 channel=17
    -37, -114, 62, -82, 14, -132, -199, 100, -40,
    -- filter=52 channel=18
    -131, -37, -36, -6, 81, -23, -187, 151, 24,
    -- filter=52 channel=19
    -89, 47, 190, -196, -215, 109, 33, -125, -257,
    -- filter=52 channel=20
    -33, -82, -95, -99, -132, -30, 188, 1, 17,
    -- filter=52 channel=21
    -92, 53, -185, 47, 47, -1, 87, 55, 146,
    -- filter=52 channel=22
    137, -227, 98, 32, 61, 138, 122, 74, -36,
    -- filter=52 channel=23
    6, 9, 23, -6, 135, -81, -133, 239, 4,
    -- filter=52 channel=24
    76, -62, -134, -19, -71, 24, 404, 10, 19,
    -- filter=52 channel=25
    -179, -48, -102, 40, 118, -26, 60, 47, -8,
    -- filter=52 channel=26
    -52, 248, -59, 47, -194, -48, -161, -296, -26,
    -- filter=52 channel=27
    -20, 121, 52, -31, 100, -65, 115, 0, -65,
    -- filter=52 channel=28
    -66, 102, 10, -158, -32, -17, -13, 176, -125,
    -- filter=52 channel=29
    86, 31, 119, -74, 10, 35, -45, -70, -73,
    -- filter=52 channel=30
    -62, 1, 154, -310, -10, 86, -7, -34, 143,
    -- filter=52 channel=31
    -75, -109, 137, -130, -7, -49, 140, 30, 143,
    -- filter=53 channel=0
    -36, 1, -274, 100, 101, -102, 50, 109, 143,
    -- filter=53 channel=1
    -189, -26, 141, -52, -105, 34, 38, 35, 9,
    -- filter=53 channel=2
    25, -46, 15, -45, 196, 66, 27, -110, -183,
    -- filter=53 channel=3
    -276, 74, 122, 102, 144, -75, -105, -162, -196,
    -- filter=53 channel=4
    -367, 76, 165, -7, 127, -7, 196, 33, 120,
    -- filter=53 channel=5
    -25, 42, -170, -71, -30, -182, -58, -17, -72,
    -- filter=53 channel=6
    -37, -66, -201, 207, 106, 8, -149, 28, 5,
    -- filter=53 channel=7
    28, 188, 52, -60, -207, 165, 117, -37, 104,
    -- filter=53 channel=8
    72, -147, -33, -34, 119, -87, -5, 57, 32,
    -- filter=53 channel=9
    -114, -366, -45, 2, 38, 43, 0, 151, 57,
    -- filter=53 channel=10
    3, -32, -86, -94, -60, 19, 107, 22, -35,
    -- filter=53 channel=11
    119, 121, 189, -159, -208, -184, -99, -3, 130,
    -- filter=53 channel=12
    -21, -141, -42, 55, 78, 146, -11, -83, -136,
    -- filter=53 channel=13
    -5, 11, -19, 23, 27, -3, -10, 14, -4,
    -- filter=53 channel=14
    0, 68, -24, -102, 76, -4, 55, 63, -89,
    -- filter=53 channel=15
    -90, 127, -118, 117, -156, -5, -6, 51, 154,
    -- filter=53 channel=16
    62, 138, -195, -142, -163, 53, 37, 85, -59,
    -- filter=53 channel=17
    59, 64, 12, -307, 12, -459, 94, -228, 58,
    -- filter=53 channel=18
    -15, -26, -365, 97, 17, 99, -149, -202, 168,
    -- filter=53 channel=19
    33, 24, 6, 83, -101, -78, -240, -135, 142,
    -- filter=53 channel=20
    26, -222, 40, 104, -51, -117, 73, 22, 101,
    -- filter=53 channel=21
    -158, -177, -210, 136, 89, 1, -53, 3, -5,
    -- filter=53 channel=22
    -141, -21, 0, -114, -84, 190, -33, 210, -68,
    -- filter=53 channel=23
    150, 158, 128, -197, -183, 153, -145, -86, -29,
    -- filter=53 channel=24
    281, -87, 36, -55, 67, 8, 47, -124, 78,
    -- filter=53 channel=25
    111, -98, -71, 93, 110, -32, -37, -111, -130,
    -- filter=53 channel=26
    216, 39, -5, 80, 183, -94, -40, -439, -227,
    -- filter=53 channel=27
    -208, -109, -50, -227, 105, -1, 150, 28, -121,
    -- filter=53 channel=28
    60, -223, -52, 14, 99, -156, 124, 12, 134,
    -- filter=53 channel=29
    -6, 183, 149, -248, 84, 124, -71, -67, -87,
    -- filter=53 channel=30
    -61, -11, -8, -71, 240, 216, -277, -156, -108,
    -- filter=53 channel=31
    -262, -96, 27, -47, 272, 49, 5, -100, -59,
    -- filter=54 channel=0
    7, 0, -26, -7, -4, 0, -10, -7, 3,
    -- filter=54 channel=1
    -24, -2, -25, -24, -27, -23, 11, -20, -25,
    -- filter=54 channel=2
    9, 0, -16, 10, 11, -4, 4, -20, 4,
    -- filter=54 channel=3
    11, 14, 3, -22, -19, 10, 3, -17, 10,
    -- filter=54 channel=4
    -25, -6, -9, -31, 0, -4, 2, 5, -23,
    -- filter=54 channel=5
    -4, -24, -35, 22, -19, 5, -4, 10, 3,
    -- filter=54 channel=6
    -29, -16, -18, -19, -5, -27, -32, 2, -11,
    -- filter=54 channel=7
    -5, 7, -21, -33, -28, -5, 0, -9, -15,
    -- filter=54 channel=8
    -34, -1, -39, -15, -34, -30, -32, -4, -20,
    -- filter=54 channel=9
    15, -17, 5, -18, 0, 0, -13, -21, -8,
    -- filter=54 channel=10
    13, -11, -24, -19, -12, 3, -32, 0, -14,
    -- filter=54 channel=11
    -3, -18, 3, 9, 2, -15, -1, -2, 5,
    -- filter=54 channel=12
    -17, -13, 9, -1, -8, 5, -9, -26, 7,
    -- filter=54 channel=13
    8, -12, -21, -5, 0, -18, 3, -20, 0,
    -- filter=54 channel=14
    -33, -19, 1, -23, -2, -7, -9, 8, -34,
    -- filter=54 channel=15
    -29, -24, -4, -16, -6, -21, 0, -12, 8,
    -- filter=54 channel=16
    0, -9, -17, -23, 6, -7, -23, -5, -4,
    -- filter=54 channel=17
    17, -17, 8, 19, 6, 6, 7, -1, 5,
    -- filter=54 channel=18
    8, 3, -15, 6, -25, -11, -17, -13, -5,
    -- filter=54 channel=19
    -6, -11, -33, -5, -14, -4, -24, -4, 4,
    -- filter=54 channel=20
    -29, -13, -9, -1, -17, 3, 15, 19, -17,
    -- filter=54 channel=21
    -2, -12, -18, -31, -9, -20, -37, -1, -7,
    -- filter=54 channel=22
    -16, -26, -25, -22, -21, -21, 11, 13, -8,
    -- filter=54 channel=23
    -37, -32, -32, 20, -19, -5, -14, -15, -23,
    -- filter=54 channel=24
    -15, -6, -4, -30, -31, -28, -23, -11, -27,
    -- filter=54 channel=25
    -5, -3, 6, 3, 7, 16, -3, -15, 16,
    -- filter=54 channel=26
    -1, -22, -3, 12, -2, 10, -11, -21, -3,
    -- filter=54 channel=27
    -17, -28, -1, -5, 2, -25, -17, -1, -2,
    -- filter=54 channel=28
    -17, 0, -5, 12, -29, -6, 8, 3, 5,
    -- filter=54 channel=29
    -18, -5, -8, 2, -14, -1, 5, -11, 3,
    -- filter=54 channel=30
    6, -16, -4, 4, -13, 4, -2, -18, 9,
    -- filter=54 channel=31
    0, 0, 9, 3, -9, -22, -3, -43, 3,
    -- filter=55 channel=0
    -48, -118, -60, -13, -397, -34, -64, -158, -59,
    -- filter=55 channel=1
    -308, -54, 47, 141, -101, 133, -111, 133, 41,
    -- filter=55 channel=2
    -178, 80, -61, 23, -19, -32, -134, 101, 86,
    -- filter=55 channel=3
    -126, -7, -205, 34, -70, -98, 180, 1, -57,
    -- filter=55 channel=4
    -157, -218, 84, 7, 158, -58, 147, -397, -7,
    -- filter=55 channel=5
    -242, -31, -94, -460, -10, -20, -173, 102, -121,
    -- filter=55 channel=6
    -237, 248, -19, -110, -41, -37, 194, -89, 24,
    -- filter=55 channel=7
    -215, 28, -18, -40, -509, -270, -284, -154, 124,
    -- filter=55 channel=8
    -293, -22, -30, 16, -261, -53, -51, -25, 103,
    -- filter=55 channel=9
    -135, -31, 24, 174, -62, -75, 174, 194, 0,
    -- filter=55 channel=10
    -114, -123, 69, 156, -126, -83, 88, -113, -149,
    -- filter=55 channel=11
    -75, 122, 47, -94, 16, 20, -101, -4, -69,
    -- filter=55 channel=12
    -111, -4, -171, 223, 196, -14, 67, -367, 18,
    -- filter=55 channel=13
    8, 12, -2, -17, 15, -3, -11, -6, 8,
    -- filter=55 channel=14
    -84, -83, 197, 0, 73, 82, -113, -83, -41,
    -- filter=55 channel=15
    101, 130, -77, 143, -62, -93, 94, 53, 150,
    -- filter=55 channel=16
    99, 40, 0, 31, -364, -63, 37, -15, -219,
    -- filter=55 channel=17
    20, 96, -196, 95, 185, -27, 59, 46, 242,
    -- filter=55 channel=18
    35, 61, -38, -175, -20, 6, 40, 47, 222,
    -- filter=55 channel=19
    -91, -102, -6, -121, 116, 51, 15, -114, 68,
    -- filter=55 channel=20
    -378, -4, 104, -2, -93, -28, -14, 26, -10,
    -- filter=55 channel=21
    165, -3, 97, -80, 129, -62, 27, -22, -164,
    -- filter=55 channel=22
    -123, -115, -31, 155, -17, 86, 235, 40, 197,
    -- filter=55 channel=23
    50, -175, 164, 51, -31, -18, 76, -38, 39,
    -- filter=55 channel=24
    -81, 67, 58, 188, 71, 128, -316, 46, 137,
    -- filter=55 channel=25
    -131, 100, 33, -186, 57, -24, -97, -71, -37,
    -- filter=55 channel=26
    129, 56, 119, 33, -20, -137, 80, -4, 15,
    -- filter=55 channel=27
    -38, -82, 52, -313, 68, -206, 31, -48, -15,
    -- filter=55 channel=28
    206, -48, 23, 75, 162, -459, 33, -53, 95,
    -- filter=55 channel=29
    -54, 30, -5, -165, -165, 216, -265, -79, -4,
    -- filter=55 channel=30
    35, 64, -219, -249, 314, 22, -33, 166, -54,
    -- filter=55 channel=31
    44, 127, 122, 159, -156, 77, -72, -91, -31,
    -- filter=56 channel=0
    -197, -65, -7, -152, -173, 65, 60, -30, -113,
    -- filter=56 channel=1
    185, 128, 91, -77, 181, 22, -34, 128, -68,
    -- filter=56 channel=2
    -130, 37, 14, 30, -28, -147, -98, -205, -102,
    -- filter=56 channel=3
    -470, -266, -10, -184, 75, -169, -23, -46, -104,
    -- filter=56 channel=4
    -23, -169, -86, -31, -434, -453, -38, 71, 0,
    -- filter=56 channel=5
    -56, 165, 115, -62, -67, 103, 71, 19, -43,
    -- filter=56 channel=6
    10, -41, 175, -15, 124, 56, -43, 100, -79,
    -- filter=56 channel=7
    46, 92, -54, 46, -94, -129, -128, -231, -108,
    -- filter=56 channel=8
    152, -52, 24, 63, 77, -89, -135, -17, 85,
    -- filter=56 channel=9
    18, -116, 82, 46, -126, 60, 76, -185, 69,
    -- filter=56 channel=10
    1, -174, -36, 65, 72, -44, -75, 110, -6,
    -- filter=56 channel=11
    21, 31, -177, -143, 187, 30, -126, 20, -237,
    -- filter=56 channel=12
    -34, -156, -409, -18, -209, -213, 53, 112, 204,
    -- filter=56 channel=13
    -12, -3, -8, -20, -7, -6, -11, 21, -9,
    -- filter=56 channel=14
    176, -156, -79, -89, -189, 144, -16, 69, -136,
    -- filter=56 channel=15
    40, -265, -211, -51, 79, -68, -39, -306, 46,
    -- filter=56 channel=16
    38, -6, 28, -31, 81, -53, 90, -245, -88,
    -- filter=56 channel=17
    -200, 49, 14, -34, 171, 167, -52, -50, -11,
    -- filter=56 channel=18
    -60, 10, -228, 2, 199, -178, 0, 46, -261,
    -- filter=56 channel=19
    21, 114, -26, -92, 184, 61, 29, 33, 43,
    -- filter=56 channel=20
    -18, -98, 124, -90, 209, 60, 250, -115, 145,
    -- filter=56 channel=21
    41, -117, 99, 20, 79, -152, 68, 224, -148,
    -- filter=56 channel=22
    -206, 216, 119, 146, -112, 199, 90, 175, 18,
    -- filter=56 channel=23
    49, 66, 2, 221, -152, -4, 10, -3, -287,
    -- filter=56 channel=24
    -98, -232, -20, 25, 14, -160, 71, -113, -204,
    -- filter=56 channel=25
    -317, 59, 53, -67, 13, 187, -530, -207, -38,
    -- filter=56 channel=26
    -259, 86, 152, -36, -83, 101, 241, -67, 56,
    -- filter=56 channel=27
    95, 53, -265, 75, 85, 90, -7, -167, -58,
    -- filter=56 channel=28
    -102, -23, 37, 255, -56, 3, 186, -33, -97,
    -- filter=56 channel=29
    119, 82, 30, -17, -69, 168, 49, 117, 204,
    -- filter=56 channel=30
    -12, 229, 80, 80, -10, 201, -93, 144, -30,
    -- filter=56 channel=31
    -45, 54, -51, 30, -30, -66, -33, -81, 44,
    -- filter=57 channel=0
    23, 11, 54, -70, -75, -79, -19, 54, 88,
    -- filter=57 channel=1
    -269, 152, -222, -68, 221, 21, 45, 80, 38,
    -- filter=57 channel=2
    1, -96, -1, -9, -2, -9, -285, 135, 62,
    -- filter=57 channel=3
    -23, -219, 21, 155, -200, -34, 126, 50, 16,
    -- filter=57 channel=4
    126, -57, -203, 25, -61, -142, 226, -223, 7,
    -- filter=57 channel=5
    86, 146, -52, -134, -68, 38, 20, 0, 48,
    -- filter=57 channel=6
    -13, 202, 22, -40, 160, 47, 41, -111, 26,
    -- filter=57 channel=7
    28, 185, -104, 0, 57, 77, -65, -333, -104,
    -- filter=57 channel=8
    -210, 40, 98, -167, 36, -45, -276, 49, 66,
    -- filter=57 channel=9
    157, 31, -135, 177, -57, 43, 80, 167, -177,
    -- filter=57 channel=10
    71, -124, 76, -160, -43, 222, -158, -28, 171,
    -- filter=57 channel=11
    -22, 67, 159, 165, 9, -67, -195, -144, 46,
    -- filter=57 channel=12
    -66, -14, 243, -242, 4, 50, -160, 180, -127,
    -- filter=57 channel=13
    -3, -8, 10, 8, -13, -12, -9, -8, 21,
    -- filter=57 channel=14
    5, -46, -195, 120, -90, -140, 307, -17, 3,
    -- filter=57 channel=15
    -25, -170, -240, -38, 82, -89, 18, 138, 220,
    -- filter=57 channel=16
    -40, -26, 57, -8, 60, 143, -51, -121, 94,
    -- filter=57 channel=17
    31, -1, -46, -43, -39, 42, 310, -119, 174,
    -- filter=57 channel=18
    98, 186, -68, -48, -101, -109, -142, 8, -25,
    -- filter=57 channel=19
    -24, -49, 78, -3, 94, 55, -111, 250, 88,
    -- filter=57 channel=20
    -174, -73, 188, -17, 91, 107, 70, -153, 103,
    -- filter=57 channel=21
    -425, -89, 140, -40, 10, -33, 16, 207, 105,
    -- filter=57 channel=22
    52, 56, -236, -59, 13, 0, 124, 60, 123,
    -- filter=57 channel=23
    85, -76, -37, 64, -174, -36, 54, 142, 19,
    -- filter=57 channel=24
    -100, -9, 49, 80, -164, 141, -88, -8, -8,
    -- filter=57 channel=25
    -161, 109, -6, 47, 52, -49, -95, 166, -195,
    -- filter=57 channel=26
    -188, 243, 111, -142, 110, -58, 28, 111, 26,
    -- filter=57 channel=27
    -164, -32, 168, -3, -36, 150, 76, -245, 194,
    -- filter=57 channel=28
    -182, -7, 85, -331, -203, 240, -109, 230, 98,
    -- filter=57 channel=29
    -90, 118, -10, -93, -38, -163, -266, 54, 0,
    -- filter=57 channel=30
    -59, -108, 80, -142, 201, -115, -159, -119, 18,
    -- filter=57 channel=31
    9, -115, -227, 35, 50, -110, -21, 26, -121,
    -- filter=58 channel=0
    70, 36, -85, 136, -41, -50, 83, -19, -23,
    -- filter=58 channel=1
    28, 38, -49, 39, -25, -93, 229, 121, -120,
    -- filter=58 channel=2
    -84, -49, 41, 255, 70, -87, 123, -110, 116,
    -- filter=58 channel=3
    -202, -140, 153, -12, -181, 18, 12, 151, 39,
    -- filter=58 channel=4
    -134, -52, -329, -144, -117, -32, -192, -446, -296,
    -- filter=58 channel=5
    22, -111, -14, 89, -133, -143, -13, -77, 22,
    -- filter=58 channel=6
    -78, 65, 110, -51, 132, -90, 76, 92, -48,
    -- filter=58 channel=7
    -88, 24, 0, 34, 111, 19, 64, 28, 122,
    -- filter=58 channel=8
    114, -140, 61, -150, 66, 35, -124, -191, 96,
    -- filter=58 channel=9
    171, 27, -7, 132, 9, -89, -125, -115, -774,
    -- filter=58 channel=10
    -23, 7, -134, 39, 281, -48, 119, -250, -42,
    -- filter=58 channel=11
    67, -50, 68, 52, -182, -142, 102, 62, -149,
    -- filter=58 channel=12
    -131, -72, 191, 224, 168, 146, 35, 61, -134,
    -- filter=58 channel=13
    -16, 22, 19, -16, 16, 0, -6, -22, -21,
    -- filter=58 channel=14
    -13, 59, -43, 40, -106, -18, 49, 66, 79,
    -- filter=58 channel=15
    47, -131, 0, 35, -30, 41, 234, 62, -96,
    -- filter=58 channel=16
    0, 5, -269, 114, -35, 40, 140, -16, 118,
    -- filter=58 channel=17
    -15, 82, -38, -50, 118, 224, -44, -216, 53,
    -- filter=58 channel=18
    -191, -149, 134, -81, -11, 42, 31, -11, 14,
    -- filter=58 channel=19
    -136, -198, 15, -184, 245, 129, 51, 140, -100,
    -- filter=58 channel=20
    171, 25, 55, 71, -208, -95, 0, 170, 9,
    -- filter=58 channel=21
    -104, 372, -13, 54, 20, -57, 311, -113, -727,
    -- filter=58 channel=22
    3, 7, 56, -65, 27, -45, 50, -187, -105,
    -- filter=58 channel=23
    -37, -16, 142, -16, -56, -64, -70, 94, 51,
    -- filter=58 channel=24
    -217, 225, 14, -213, 157, -2, -157, 39, -81,
    -- filter=58 channel=25
    4, 4, 141, 9, 41, -54, -60, -1, -63,
    -- filter=58 channel=26
    -9, -52, 88, 143, 58, 58, -47, 82, 130,
    -- filter=58 channel=27
    176, 64, 150, 139, 14, 91, -114, -3, -63,
    -- filter=58 channel=28
    -126, 159, -96, 83, -716, -231, -372, -38, -559,
    -- filter=58 channel=29
    119, -126, 40, 10, -170, 52, 74, -14, 84,
    -- filter=58 channel=30
    0, -131, -172, -244, 37, -48, -15, 263, 4,
    -- filter=58 channel=31
    -112, -135, 154, 36, -112, -51, 55, -140, 44,
    -- filter=59 channel=0
    -455, -162, -32, -323, -260, -126, -330, -52, -106,
    -- filter=59 channel=1
    151, -46, 131, 425, -41, -50, 60, 31, 0,
    -- filter=59 channel=2
    28, 30, -112, 119, 120, 45, 57, 149, -7,
    -- filter=59 channel=3
    16, -196, -207, 51, 34, 178, 61, 169, -80,
    -- filter=59 channel=4
    -364, -502, -174, -373, -718, -167, -209, -322, -210,
    -- filter=59 channel=5
    36, 19, -57, 59, 42, 89, -284, -14, -382,
    -- filter=59 channel=6
    163, -108, 21, 206, 129, 22, -79, -258, 225,
    -- filter=59 channel=7
    -99, -208, 55, 72, 151, 118, 139, 63, 84,
    -- filter=59 channel=8
    61, 138, -103, 260, -189, -355, 69, -104, -132,
    -- filter=59 channel=9
    20, 121, 133, 26, -189, 12, 119, -10, 69,
    -- filter=59 channel=10
    26, 30, -78, 32, -85, 151, 136, -116, 70,
    -- filter=59 channel=11
    5, -228, 17, 35, 50, -107, 112, -95, 70,
    -- filter=59 channel=12
    -48, -62, -274, -173, 21, -59, 47, -195, -82,
    -- filter=59 channel=13
    3, -19, -11, 15, 5, -2, 10, -21, 17,
    -- filter=59 channel=14
    -295, -175, -206, -296, -607, -82, -312, -180, 79,
    -- filter=59 channel=15
    -209, -175, -190, 38, 88, 20, 248, 141, -37,
    -- filter=59 channel=16
    239, -63, -43, 131, 61, 9, 200, 40, -554,
    -- filter=59 channel=17
    -27, 255, -151, 106, -240, 14, 26, -53, -463,
    -- filter=59 channel=18
    -90, -44, 47, -64, -135, 108, 22, 0, -7,
    -- filter=59 channel=19
    -192, 165, -60, 132, 194, 45, 107, 56, -37,
    -- filter=59 channel=20
    68, 143, 41, -146, 94, -243, -16, -391, 136,
    -- filter=59 channel=21
    143, 111, -163, -19, -53, -143, -54, 63, 118,
    -- filter=59 channel=22
    29, -89, 11, -40, 80, -34, -310, -10, 122,
    -- filter=59 channel=23
    -137, 94, -11, -210, 64, 2, -455, 69, 209,
    -- filter=59 channel=24
    -123, 45, 72, -66, -119, 54, 105, 0, 106,
    -- filter=59 channel=25
    -133, -73, 27, -309, 73, -118, -84, 99, 98,
    -- filter=59 channel=26
    -125, 246, 37, -4, 36, -13, -126, 2, -97,
    -- filter=59 channel=27
    166, 0, 88, 106, -53, 21, -238, 100, 39,
    -- filter=59 channel=28
    233, -241, -46, 96, -158, -86, 122, 56, 0,
    -- filter=59 channel=29
    48, -60, 69, 144, -172, -154, -37, -14, -259,
    -- filter=59 channel=30
    -115, -45, 138, -126, -32, 32, -257, 95, -131,
    -- filter=59 channel=31
    223, 145, -109, 14, -217, -124, -190, -51, 180,
    -- filter=60 channel=0
    -64, 15, 67, 20, 224, 162, 198, 71, 125,
    -- filter=60 channel=1
    -99, 0, 44, 17, -93, 73, 110, 100, 328,
    -- filter=60 channel=2
    111, 4, -45, 205, -56, 167, -163, -13, -22,
    -- filter=60 channel=3
    -173, -47, -149, -374, 20, -104, 22, -157, -102,
    -- filter=60 channel=4
    44, 72, -34, -33, 95, 5, 48, 63, 0,
    -- filter=60 channel=5
    45, 40, -66, 13, 62, 81, -112, -85, -76,
    -- filter=60 channel=6
    174, 178, -173, 17, -41, 41, -272, -58, 248,
    -- filter=60 channel=7
    184, 160, -57, -158, -89, -483, -272, -18, -168,
    -- filter=60 channel=8
    151, -163, -92, 25, -62, -210, 202, -120, -419,
    -- filter=60 channel=9
    -83, -261, 58, -23, 166, 120, -77, -32, -135,
    -- filter=60 channel=10
    -28, 28, 158, -232, -170, -142, 6, -29, -73,
    -- filter=60 channel=11
    -104, 120, 139, -10, 21, -80, 98, 132, 102,
    -- filter=60 channel=12
    100, 66, 84, -28, 128, 49, -102, -2, 106,
    -- filter=60 channel=13
    -21, 5, 0, -13, 7, -6, -9, 13, 13,
    -- filter=60 channel=14
    -107, 0, -1, 67, 108, 147, 122, 33, -43,
    -- filter=60 channel=15
    193, 84, -27, -28, -37, -139, 73, -270, -271,
    -- filter=60 channel=16
    12, -45, 56, -128, -49, -42, 19, 61, 0,
    -- filter=60 channel=17
    -40, 123, 74, -5, 173, 32, -48, -45, -103,
    -- filter=60 channel=18
    -12, 25, 98, -308, 151, 142, -193, -62, -33,
    -- filter=60 channel=19
    75, -39, 153, -76, 30, -302, 150, -53, 133,
    -- filter=60 channel=20
    -131, 133, 16, 5, -39, 91, 100, -6, -76,
    -- filter=60 channel=21
    -55, 148, -9, 123, -149, -145, 56, -293, -84,
    -- filter=60 channel=22
    -32, -3, 392, -53, -87, 125, -235, 73, 84,
    -- filter=60 channel=23
    -32, -58, 29, 95, 125, -37, 11, -78, -242,
    -- filter=60 channel=24
    -68, -147, -170, 97, 139, 27, 88, 142, 81,
    -- filter=60 channel=25
    195, 56, 8, -133, 94, 6, -175, -48, 204,
    -- filter=60 channel=26
    -115, -208, -13, 61, 76, 4, -62, -116, -51,
    -- filter=60 channel=27
    52, -29, -147, 78, -155, -75, -109, -46, -124,
    -- filter=60 channel=28
    169, -262, 25, 32, 112, -111, 122, -90, 99,
    -- filter=60 channel=29
    -56, -91, -31, -46, 5, 13, 53, -99, -276,
    -- filter=60 channel=30
    -243, 79, 20, -319, 102, -118, 27, -31, 154,
    -- filter=60 channel=31
    -51, -38, -103, -83, -167, 14, -88, 164, 15,
    -- filter=61 channel=0
    56, -29, 52, -66, -53, 14, -37, -3, -184,
    -- filter=61 channel=1
    -7, -36, 76, 143, -17, 267, -27, 92, 193,
    -- filter=61 channel=2
    -163, 4, 235, -85, -117, 92, -92, -184, 390,
    -- filter=61 channel=3
    8, -124, -105, 59, -40, -89, -180, 68, -49,
    -- filter=61 channel=4
    137, 58, 0, 7, -2, 126, -40, -180, -166,
    -- filter=61 channel=5
    105, 159, -205, -80, 61, -38, 6, 6, 134,
    -- filter=61 channel=6
    66, -124, 37, 71, -175, -12, -167, -22, 55,
    -- filter=61 channel=7
    -72, -130, -216, -33, -265, -83, 57, -148, -8,
    -- filter=61 channel=8
    -31, 9, -21, -82, 25, -230, 31, -6, -35,
    -- filter=61 channel=9
    43, -78, -59, 23, -205, -21, 30, -18, -80,
    -- filter=61 channel=10
    57, -64, 117, 103, 46, -9, 270, 130, 92,
    -- filter=61 channel=11
    -62, 11, 19, -116, -52, -140, 148, 65, -70,
    -- filter=61 channel=12
    16, 170, 117, 139, 8, -8, 44, 105, 100,
    -- filter=61 channel=13
    7, 10, -3, -13, -11, -2, 3, 5, -3,
    -- filter=61 channel=14
    31, 4, -38, -9, -45, 7, -32, -208, -259,
    -- filter=61 channel=15
    -6, 24, -74, -98, -267, -5, 35, 380, -189,
    -- filter=61 channel=16
    37, -38, -43, 97, -64, -238, -15, 138, 178,
    -- filter=61 channel=17
    -385, 53, 87, -91, 182, 145, -209, 224, 130,
    -- filter=61 channel=18
    -72, -74, 260, 44, 71, -303, 111, -96, -172,
    -- filter=61 channel=19
    -64, -383, -13, 3, -127, 198, 109, -30, 71,
    -- filter=61 channel=20
    -68, -15, -63, 42, -191, -63, 60, -116, 53,
    -- filter=61 channel=21
    -126, -33, -60, 386, -9, 74, 236, 3, -209,
    -- filter=61 channel=22
    -42, -89, 79, -181, -74, 276, -81, -101, -120,
    -- filter=61 channel=23
    -84, -231, 7, -6, 102, 42, 44, 266, -59,
    -- filter=61 channel=24
    52, -10, 42, 14, -3, -219, 27, 90, -72,
    -- filter=61 channel=25
    133, 24, 19, 81, 186, -15, -72, 114, -149,
    -- filter=61 channel=26
    -43, -151, 157, 120, 215, -97, 18, -358, -164,
    -- filter=61 channel=27
    -308, -242, -83, -15, -80, -343, 107, 93, -89,
    -- filter=61 channel=28
    18, 8, 104, -304, -8, 138, 158, -101, -194,
    -- filter=61 channel=29
    -5, -113, -80, 173, 43, -129, -128, -47, 201,
    -- filter=61 channel=30
    35, -204, -265, 128, 165, -155, 32, 161, -30,
    -- filter=61 channel=31
    -141, -128, -65, 57, -38, -158, 96, 14, 15,
    -- filter=62 channel=0
    113, 133, -52, 69, 30, 34, -41, 225, 66,
    -- filter=62 channel=1
    -21, 75, -47, -31, -71, 167, -130, 70, 16,
    -- filter=62 channel=2
    6, 37, -3, -165, 58, 100, -190, -18, -8,
    -- filter=62 channel=3
    -104, 24, -213, 68, 89, -31, -167, 104, -160,
    -- filter=62 channel=4
    51, -19, 7, -1, 29, -187, 47, -43, 121,
    -- filter=62 channel=5
    0, 9, 41, 83, -129, -19, -159, -114, -206,
    -- filter=62 channel=6
    -3, -88, -57, 125, 98, -63, 76, -91, 20,
    -- filter=62 channel=7
    -41, -105, 127, 87, -69, 16, -47, -54, 71,
    -- filter=62 channel=8
    99, 44, 56, -65, 133, -7, -132, 11, 20,
    -- filter=62 channel=9
    34, 82, -19, 0, 211, 19, 138, 71, -71,
    -- filter=62 channel=10
    40, 69, 13, -55, 41, -154, -59, 65, -146,
    -- filter=62 channel=11
    -31, 103, 24, -34, -32, 219, 23, 76, 107,
    -- filter=62 channel=12
    -6, 46, 112, -47, -22, -257, -80, -411, -210,
    -- filter=62 channel=13
    -11, 15, 3, -25, 22, 3, 12, -12, 18,
    -- filter=62 channel=14
    -119, 4, -96, 87, 56, 73, 126, 114, 208,
    -- filter=62 channel=15
    -46, -53, -150, -127, -40, 10, -54, 151, 3,
    -- filter=62 channel=16
    -41, -112, -49, -181, -80, -190, 11, -84, -61,
    -- filter=62 channel=17
    14, -16, 113, 40, -138, -14, 60, -129, -48,
    -- filter=62 channel=18
    24, 14, -128, -26, 61, -64, -319, 247, 45,
    -- filter=62 channel=19
    29, -161, 154, -172, 98, 2, -21, 135, -34,
    -- filter=62 channel=20
    -11, -53, 2, -81, 155, 70, -138, 0, 73,
    -- filter=62 channel=21
    15, -17, 153, -267, -59, 6, -77, -33, 2,
    -- filter=62 channel=22
    -73, -54, -26, -45, -29, 150, 101, 6, -57,
    -- filter=62 channel=23
    30, -33, -60, 22, 27, 48, 52, -2, 125,
    -- filter=62 channel=24
    -3, -97, 3, 45, -162, 3, -145, -152, -104,
    -- filter=62 channel=25
    112, -121, -84, -68, -96, -94, -402, 13, -303,
    -- filter=62 channel=26
    -2, -378, 71, -36, 2, -69, 28, 22, -114,
    -- filter=62 channel=27
    -70, -9, -29, 81, 93, -131, 106, 45, 106,
    -- filter=62 channel=28
    -47, -17, 201, -41, 69, -99, 111, 48, 108,
    -- filter=62 channel=29
    -64, 88, -172, 52, 2, 208, 14, -21, 30,
    -- filter=62 channel=30
    -246, -18, 69, -54, 61, -16, -50, 20, 7,
    -- filter=62 channel=31
    -29, 157, -73, 217, -59, -183, 87, -52, -127,
    -- filter=63 channel=0
    46, 117, -11, 44, 68, -201, 131, 56, 50,
    -- filter=63 channel=1
    46, -7, 95, -149, 32, 58, 16, -103, -77,
    -- filter=63 channel=2
    -109, 13, -95, -41, 36, 42, 120, 122, -58,
    -- filter=63 channel=3
    52, -48, 150, 6, 12, -93, -171, 42, -86,
    -- filter=63 channel=4
    18, 3, 73, 81, 84, 47, 2, 144, -157,
    -- filter=63 channel=5
    133, -44, 119, -42, -82, -130, 7, -55, 36,
    -- filter=63 channel=6
    50, -105, 245, 18, -43, 309, -74, -74, 5,
    -- filter=63 channel=7
    11, -68, 3, 5, -49, 8, 0, -115, -23,
    -- filter=63 channel=8
    110, -30, 42, 22, -161, 63, -92, -15, 17,
    -- filter=63 channel=9
    252, 112, 32, -2, 145, 160, 35, -97, -78,
    -- filter=63 channel=10
    -164, 51, 50, 84, 45, -33, 100, -82, 134,
    -- filter=63 channel=11
    24, 46, 8, 14, -12, 44, 55, -125, 42,
    -- filter=63 channel=12
    81, 216, 231, 1, 59, -59, -6, 38, -103,
    -- filter=63 channel=13
    13, 0, 11, 22, -7, -8, 28, -2, -2,
    -- filter=63 channel=14
    45, 70, 3, 66, 71, -34, 141, 64, 32,
    -- filter=63 channel=15
    -170, -210, 45, -36, -138, -9, -113, 29, 190,
    -- filter=63 channel=16
    -3, -57, -103, 21, 22, 140, 29, 26, -75,
    -- filter=63 channel=17
    125, -88, 188, -18, 137, 1, -117, 84, 155,
    -- filter=63 channel=18
    83, 218, 21, 71, 6, -99, -68, 82, -40,
    -- filter=63 channel=19
    110, 183, 135, -178, -23, 140, -358, -144, 118,
    -- filter=63 channel=20
    -132, -217, -49, -86, -290, -29, 143, -220, -53,
    -- filter=63 channel=21
    -7, 1, 70, -53, -26, 46, -51, 3, 61,
    -- filter=63 channel=22
    -74, -143, -126, -52, 126, 221, -78, 0, 48,
    -- filter=63 channel=23
    -33, -2, 30, 50, -77, -137, 105, -67, -7,
    -- filter=63 channel=24
    123, -40, 25, 2, 76, 74, 89, 15, 58,
    -- filter=63 channel=25
    -7, -19, -21, -51, 107, 112, 22, 0, 93,
    -- filter=63 channel=26
    3, 151, -194, -76, -147, 131, 3, -78, 80,
    -- filter=63 channel=27
    22, 11, 19, 53, 174, 76, -116, 18, 40,
    -- filter=63 channel=28
    24, -29, 66, 24, 12, -10, -103, 100, 20,
    -- filter=63 channel=29
    7, 79, -117, -136, 92, 63, -124, -52, -23,
    -- filter=63 channel=30
    75, 83, 62, 48, 26, 39, -176, 45, -9,
    -- filter=63 channel=31
    -178, -59, -13, 6, 151, -83, 62, -86, -32,

    -- ifmap
    -- channel=0
    0, 0, 0, 0, 278, 0, 85, 
    407, 0, 183, 82, 0, 0, 0, 
    0, 0, 204, 71, 38, 242, 39, 
    0, 23, 0, 94, 0, 0, 36, 
    0, 127, 107, 0, 0, 452, 0, 
    0, 0, 381, 89, 55, 0, 0, 
    23, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 144, 155, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 31, 24, 
    0, 0, 0, 15, 0, 132, 0, 
    0, 0, 0, 0, 0, 210, 0, 
    116, 0, 0, 425, 204, 5, 24, 
    0, 563, 70, 39, 21, 18, 3, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 80, 0, 0, 
    135, 0, 306, 251, 136, 245, 163, 
    0, 317, 350, 245, 218, 211, 181, 
    
    -- channel=3
    219, 336, 63, 0, 0, 0, 109, 
    0, 31, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 16, 
    117, 0, 0, 101, 0, 0, 173, 
    0, 0, 0, 0, 0, 185, 0, 
    0, 0, 0, 27, 103, 45, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 193, 0, 0, 283, 
    0, 0, 0, 83, 0, 218, 46, 
    27, 88, 0, 0, 0, 170, 0, 
    0, 0, 0, 0, 0, 82, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    265, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 323, 0, 33, 0, 
    55, 0, 0, 0, 38, 0, 4, 
    0, 0, 0, 0, 0, 9, 0, 
    10, 0, 0, 46, 0, 30, 43, 
    0, 57, 0, 0, 395, 0, 0, 
    57, 0, 155, 158, 0, 0, 0, 
    0, 281, 0, 1, 0, 0, 0, 
    
    -- channel=6
    0, 0, 83, 600, 540, 484, 284, 
    167, 0, 131, 16, 0, 0, 127, 
    0, 0, 0, 0, 0, 87, 0, 
    0, 217, 124, 86, 0, 131, 0, 
    0, 0, 59, 38, 277, 284, 0, 
    7, 27, 527, 162, 11, 0, 0, 
    34, 247, 8, 0, 0, 0, 0, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 
    120, 0, 0, 0, 0, 0, 0, 
    66, 0, 0, 0, 110, 0, 18, 
    0, 0, 0, 0, 0, 0, 87, 
    0, 66, 25, 189, 0, 4, 66, 
    0, 443, 0, 0, 32, 1, 0, 
    0, 0, 0, 0, 0, 0, 73, 
    
    -- channel=8
    15, 0, 41, 66, 10, 151, 0, 
    79, 0, 274, 225, 0, 0, 20, 
    57, 0, 0, 0, 162, 0, 0, 
    0, 0, 0, 0, 97, 0, 0, 
    0, 204, 116, 238, 115, 0, 0, 
    0, 391, 273, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 
    99, 84, 21, 0, 145, 0, 0, 
    0, 0, 0, 0, 603, 0, 0, 
    0, 0, 0, 0, 216, 0, 0, 
    0, 418, 2, 0, 0, 0, 113, 
    0, 143, 0, 0, 32, 60, 0, 
    0, 0, 148, 0, 0, 0, 0, 
    
    -- channel=10
    0, 47, 295, 478, 325, 224, 47, 
    124, 166, 153, 278, 0, 155, 0, 
    89, 0, 0, 48, 39, 95, 0, 
    124, 0, 0, 110, 0, 0, 0, 
    0, 0, 46, 229, 209, 49, 151, 
    0, 489, 118, 249, 220, 204, 156, 
    0, 60, 95, 0, 44, 2, 242, 
    
    -- channel=11
    71, 105, 54, 106, 0, 159, 228, 
    159, 84, 0, 13, 54, 0, 0, 
    170, 244, 144, 0, 0, 0, 133, 
    106, 212, 163, 34, 229, 0, 173, 
    0, 0, 354, 251, 226, 60, 180, 
    201, 79, 0, 248, 123, 103, 57, 
    49, 142, 0, 5, 4, 0, 0, 
    
    -- channel=12
    0, 0, 0, 28, 67, 265, 104, 
    0, 0, 0, 227, 0, 155, 0, 
    170, 0, 0, 433, 0, 218, 78, 
    293, 95, 0, 280, 0, 139, 0, 
    169, 138, 0, 214, 76, 54, 0, 
    0, 0, 501, 0, 226, 0, 33, 
    0, 154, 78, 59, 26, 8, 0, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    29, 0, 340, 0, 134, 0, 43, 
    26, 75, 0, 0, 126, 0, 0, 
    451, 0, 29, 0, 172, 0, 157, 
    315, 324, 391, 76, 249, 0, 168, 
    118, 0, 0, 328, 44, 0, 168, 
    50, 576, 0, 0, 47, 34, 0, 
    0, 763, 32, 12, 32, 54, 96, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 43, 88, 110, 0, 
    0, 0, 0, 83, 226, 79, 126, 
    107, 153, 0, 31, 0, 0, 23, 
    152, 88, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 200, 258, 254, 
    0, 45, 71, 165, 301, 259, 180, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 
    79, 0, 0, 0, 0, 72, 142, 
    289, 0, 0, 0, 0, 9, 30, 
    0, 0, 0, 113, 0, 0, 337, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 202, 119, 106, 0, 122, 
    240, 0, 0, 49, 29, 96, 115, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 53, 0, 0, 0, 0, 
    0, 111, 0, 0, 0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 175, 
    0, 0, 0, 0, 0, 0, 0, 
    103, 0, 0, 0, 0, 1, 79, 
    277, 0, 0, 137, 134, 177, 199, 
    
    -- channel=20
    121, 26, 128, 269, 162, 50, 126, 
    59, 279, 179, 0, 0, 40, 93, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 147, 0, 123, 0, 0, 0, 
    33, 0, 0, 0, 0, 67, 249, 
    0, 39, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    0, 66, 0, 0, 0, 0, 121, 
    115, 42, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 134, 0, 
    0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 337, 230, 230, 188, 
    213, 0, 0, 0, 176, 166, 189, 
    
    -- channel=23
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 111, 0, 56, 70, 
    0, 264, 197, 20, 0, 51, 0, 
    0, 0, 142, 32, 57, 126, 102, 
    0, 0, 0, 0, 115, 0, 0, 
    199, 50, 26, 123, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 201, 0, 130, 0, 
    0, 0, 0, 0, 0, 0, 64, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 49, 331, 160, 177, 
    18, 0, 0, 0, 191, 115, 0, 
    
    -- channel=25
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 41, 0, 
    0, 0, 5, 0, 0, 0, 0, 
    0, 0, 82, 0, 0, 0, 0, 
    183, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 235, 0, 0, 0, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 40, 0, 0, 
    80, 0, 0, 0, 15, 0, 0, 
    149, 0, 0, 0, 70, 0, 0, 
    21, 16, 0, 164, 115, 0, 0, 
    339, 385, 0, 387, 277, 325, 330, 
    453, 283, 208, 151, 193, 222, 303, 
    
    -- channel=27
    264, 0, 0, 160, 0, 8, 433, 
    12, 153, 0, 0, 251, 0, 64, 
    0, 0, 0, 0, 7, 0, 0, 
    0, 185, 46, 0, 0, 0, 143, 
    0, 0, 0, 0, 0, 62, 239, 
    283, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    271, 475, 529, 311, 60, 0, 56, 
    0, 330, 0, 0, 9, 90, 0, 
    0, 296, 0, 103, 125, 194, 0, 
    0, 0, 337, 136, 233, 219, 4, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    0, 0, 203, 0, 0, 0, 0, 
    0, 0, 48, 148, 0, 31, 0, 
    0, 380, 35, 231, 119, 46, 0, 
    0, 0, 61, 0, 124, 179, 0, 
    0, 0, 83, 83, 0, 0, 0, 
    0, 0, 264, 0, 0, 0, 0, 
    0, 0, 103, 0, 0, 0, 0, 
    
    -- channel=30
    93, 231, 0, 0, 0, 0, 0, 
    0, 80, 0, 0, 0, 0, 0, 
    49, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 47, 
    0, 0, 0, 0, 0, 0, 48, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    20, 18, 176, 92, 113, 80, 0, 
    44, 123, 78, 122, 8, 0, 0, 
    0, 102, 0, 7, 137, 0, 55, 
    134, 170, 0, 36, 67, 2, 77, 
    16, 208, 160, 98, 52, 42, 0, 
    0, 130, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end inmem_package;
