library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package inmem_package is
  type mem is array(0 to 4000000) of integer;

  constant input_mem : mem := (

    -- ifmap
    -- channel=0
    146, 118, 122, 126, 125, 121, 126, 124, 125, 123, 123, 123, 123, 125, 125, 127, 129, 126, 124, 125, 123, 120, 122, 122, 128, 124, 124, 123, 126, 126, 126, 165, 
    93, 103, 101, 113, 115, 108, 111, 112, 116, 112, 106, 104, 108, 113, 115, 121, 126, 118, 107, 102, 103, 98, 103, 102, 111, 113, 114, 113, 120, 122, 121, 213, 
    99, 111, 103, 115, 112, 110, 112, 112, 116, 116, 107, 107, 105, 112, 122, 121, 120, 110, 99, 101, 104, 97, 91, 92, 93, 97, 116, 117, 121, 123, 121, 214, 
    103, 119, 107, 117, 110, 106, 111, 113, 111, 106, 89, 120, 104, 101, 109, 105, 92, 107, 102, 104, 93, 96, 88, 84, 89, 81, 97, 110, 116, 118, 120, 218, 
    96, 108, 101, 111, 114, 105, 112, 115, 112, 97, 15, 91, 120, 99, 83, 97, 107, 107, 82, 67, 58, 74, 85, 86, 86, 84, 67, 86, 108, 120, 117, 222, 
    83, 90, 74, 107, 123, 111, 112, 121, 114, 102, 9, 68, 144, 129, 103, 104, 131, 78, 29, 40, 44, 49, 69, 80, 82, 94, 87, 67, 83, 119, 116, 220, 
    78, 120, 68, 82, 118, 116, 112, 119, 118, 110, 87, 90, 109, 129, 125, 85, 90, 57, 5, 31, 60, 57, 65, 62, 80, 105, 111, 70, 52, 103, 121, 222, 
    85, 138, 91, 54, 86, 114, 114, 112, 117, 116, 103, 96, 75, 92, 99, 63, 73, 77, 5, 0, 78, 98, 62, 53, 87, 109, 108, 97, 46, 78, 123, 225, 
    89, 128, 55, 57, 80, 105, 110, 102, 105, 137, 94, 48, 41, 70, 98, 69, 67, 81, 48, 0, 59, 107, 89, 70, 79, 104, 106, 112, 64, 46, 109, 231, 
    61, 108, 11, 31, 106, 103, 101, 41, 43, 88, 82, 0, 40, 72, 105, 86, 67, 87, 77, 21, 38, 70, 105, 84, 67, 83, 94, 122, 103, 38, 71, 231, 
    50, 34, 6, 26, 120, 109, 117, 0, 0, 27, 92, 23, 56, 86, 75, 98, 76, 112, 56, 2, 40, 31, 91, 85, 63, 78, 85, 108, 130, 76, 48, 202, 
    74, 0, 0, 38, 120, 109, 135, 12, 0, 27, 81, 25, 41, 105, 64, 88, 93, 128, 17, 0, 33, 34, 96, 95, 56, 61, 90, 91, 117, 96, 78, 175, 
    87, 4, 0, 29, 93, 112, 134, 126, 0, 10, 78, 23, 2, 97, 91, 64, 72, 143, 0, 0, 38, 70, 98, 92, 63, 47, 78, 85, 98, 89, 111, 177, 
    97, 2, 0, 58, 78, 93, 123, 157, 0, 26, 71, 25, 0, 50, 95, 73, 53, 121, 0, 0, 49, 82, 103, 85, 74, 65, 62, 69, 82, 78, 115, 197, 
    93, 0, 0, 101, 100, 52, 103, 159, 40, 38, 9, 25, 0, 15, 70, 69, 72, 105, 0, 0, 59, 76, 84, 82, 67, 70, 45, 44, 80, 85, 106, 214, 
    72, 0, 0, 87, 125, 29, 77, 139, 68, 23, 0, 0, 56, 40, 43, 52, 82, 109, 0, 0, 51, 82, 78, 92, 60, 51, 48, 44, 92, 107, 104, 218, 
    45, 0, 0, 43, 133, 18, 41, 107, 97, 1, 0, 0, 80, 102, 60, 76, 66, 94, 27, 11, 24, 91, 99, 87, 60, 37, 55, 77, 104, 103, 101, 224, 
    20, 4, 0, 3, 126, 46, 0, 77, 132, 25, 0, 40, 84, 99, 74, 84, 47, 63, 71, 75, 33, 50, 97, 105, 87, 63, 61, 99, 92, 83, 99, 231, 
    0, 15, 0, 0, 96, 93, 0, 25, 99, 84, 76, 34, 82, 68, 51, 96, 45, 4, 95, 124, 53, 36, 104, 130, 85, 89, 57, 85, 88, 94, 109, 237, 
    0, 24, 0, 0, 61, 108, 0, 15, 50, 63, 132, 11, 58, 48, 15, 94, 90, 0, 46, 65, 82, 111, 101, 103, 59, 72, 61, 74, 95, 105, 111, 232, 
    0, 33, 2, 0, 42, 97, 13, 7, 81, 47, 110, 64, 43, 11, 0, 57, 118, 57, 44, 60, 95, 128, 114, 77, 41, 39, 51, 66, 95, 88, 93, 216, 
    0, 22, 13, 0, 41, 97, 0, 0, 48, 106, 51, 14, 0, 0, 0, 23, 77, 80, 99, 95, 90, 75, 76, 51, 33, 19, 23, 39, 67, 57, 55, 187, 
    0, 0, 19, 0, 48, 102, 0, 0, 0, 46, 45, 0, 0, 0, 0, 16, 61, 66, 94, 86, 57, 35, 21, 22, 29, 18, 12, 17, 33, 32, 29, 163, 
    0, 0, 0, 0, 31, 47, 0, 0, 0, 14, 69, 64, 26, 26, 32, 32, 53, 52, 44, 33, 28, 28, 20, 18, 19, 21, 10, 9, 24, 21, 21, 166, 
    0, 0, 0, 0, 34, 0, 0, 0, 4, 70, 95, 58, 41, 37, 37, 33, 29, 33, 35, 27, 21, 25, 23, 19, 10, 12, 15, 13, 16, 15, 18, 171, 
    11, 7, 0, 0, 34, 0, 0, 0, 71, 81, 61, 33, 26, 29, 33, 34, 36, 37, 36, 29, 20, 21, 18, 7, 0, 2, 10, 6, 13, 6, 0, 172, 
    2, 27, 6, 0, 0, 0, 0, 42, 102, 70, 23, 25, 32, 30, 33, 35, 36, 33, 27, 22, 15, 4, 4, 1, 3, 7, 11, 1, 0, 0, 0, 183, 
    0, 24, 22, 13, 0, 0, 0, 102, 83, 52, 23, 17, 40, 38, 28, 27, 27, 24, 22, 15, 14, 2, 0, 7, 19, 23, 10, 0, 0, 0, 0, 191, 
    1, 15, 15, 16, 6, 0, 0, 107, 74, 35, 27, 15, 26, 36, 35, 27, 28, 22, 19, 13, 15, 16, 5, 8, 19, 24, 0, 0, 0, 38, 9, 174, 
    3, 18, 7, 15, 18, 0, 0, 60, 82, 32, 22, 13, 13, 20, 35, 32, 26, 18, 16, 20, 17, 16, 22, 17, 9, 0, 0, 0, 21, 55, 6, 146, 
    0, 36, 7, 13, 16, 31, 18, 29, 59, 46, 27, 24, 19, 19, 23, 20, 15, 14, 12, 19, 24, 24, 29, 8, 0, 0, 0, 8, 28, 42, 37, 140, 
    0, 31, 14, 11, 14, 23, 35, 32, 45, 48, 31, 37, 34, 36, 32, 22, 14, 3, 0, 5, 29, 29, 26, 0, 0, 0, 0, 27, 51, 28, 44, 149, 
    
    -- channel=1
    33, 94, 95, 98, 98, 97, 97, 98, 96, 97, 93, 95, 98, 101, 103, 100, 96, 93, 92, 92, 90, 87, 84, 84, 82, 81, 77, 75, 69, 63, 57, 0, 
    48, 156, 157, 159, 161, 159, 163, 165, 163, 161, 160, 161, 163, 166, 167, 168, 166, 163, 155, 146, 130, 123, 116, 120, 127, 130, 132, 133, 127, 122, 116, 44, 
    48, 155, 157, 155, 162, 164, 169, 171, 168, 167, 171, 177, 189, 178, 168, 171, 167, 152, 138, 116, 118, 113, 107, 99, 92, 107, 109, 126, 132, 130, 121, 47, 
    50, 159, 164, 161, 161, 164, 167, 169, 166, 168, 201, 214, 238, 191, 165, 153, 134, 103, 91, 112, 127, 124, 113, 99, 96, 89, 108, 116, 124, 129, 125, 47, 
    49, 155, 156, 153, 161, 164, 167, 166, 166, 165, 194, 199, 193, 159, 122, 94, 66, 72, 96, 114, 136, 139, 131, 113, 92, 92, 82, 86, 107, 126, 132, 52, 
    37, 119, 121, 109, 142, 168, 168, 168, 168, 167, 170, 167, 185, 144, 109, 89, 75, 79, 90, 122, 161, 160, 136, 120, 114, 92, 68, 70, 86, 110, 129, 51, 
    29, 107, 92, 104, 143, 167, 166, 167, 169, 167, 156, 143, 150, 146, 126, 97, 78, 84, 102, 136, 170, 170, 142, 123, 107, 84, 64, 42, 65, 93, 122, 53, 
    39, 130, 106, 100, 166, 176, 169, 172, 180, 167, 163, 145, 166, 171, 144, 107, 81, 84, 92, 123, 148, 165, 144, 111, 91, 81, 62, 46, 44, 69, 110, 59, 
    59, 167, 159, 151, 185, 189, 170, 187, 216, 246, 239, 222, 187, 184, 149, 114, 87, 81, 73, 91, 141, 181, 153, 118, 102, 85, 74, 50, 40, 53, 84, 45, 
    64, 215, 178, 203, 221, 197, 156, 197, 232, 293, 276, 226, 194, 197, 165, 117, 98, 60, 71, 98, 147, 211, 180, 141, 100, 89, 94, 65, 39, 33, 60, 26, 
    61, 233, 202, 224, 244, 218, 155, 167, 200, 243, 279, 251, 217, 212, 187, 131, 101, 72, 78, 117, 187, 240, 181, 140, 102, 96, 97, 89, 59, 43, 39, 10, 
    56, 232, 184, 241, 256, 219, 160, 136, 152, 207, 247, 233, 217, 241, 219, 160, 134, 87, 119, 138, 213, 238, 175, 135, 100, 97, 102, 92, 73, 63, 48, 4, 
    52, 235, 187, 237, 246, 193, 163, 134, 136, 143, 211, 223, 263, 273, 261, 192, 155, 111, 135, 151, 224, 241, 166, 126, 86, 84, 91, 100, 99, 92, 72, 20, 
    56, 250, 198, 224, 224, 183, 160, 136, 133, 115, 197, 231, 268, 269, 248, 198, 168, 132, 144, 152, 228, 230, 167, 135, 105, 93, 108, 121, 118, 115, 97, 31, 
    67, 263, 214, 232, 216, 175, 156, 151, 143, 129, 220, 260, 298, 281, 228, 197, 155, 120, 145, 158, 212, 215, 171, 113, 87, 89, 107, 125, 125, 120, 109, 50, 
    81, 278, 229, 249, 222, 189, 153, 171, 151, 143, 177, 247, 249, 203, 181, 149, 143, 129, 140, 146, 209, 201, 164, 134, 107, 93, 106, 116, 116, 120, 127, 58, 
    94, 292, 251, 264, 229, 193, 150, 169, 177, 155, 161, 177, 194, 184, 144, 129, 137, 133, 148, 143, 143, 141, 154, 112, 60, 56, 78, 101, 125, 140, 142, 64, 
    103, 297, 266, 273, 244, 205, 159, 174, 189, 174, 127, 137, 139, 167, 160, 139, 147, 142, 149, 143, 153, 148, 115, 67, 53, 41, 77, 106, 139, 149, 147, 70, 
    105, 295, 275, 273, 257, 214, 166, 151, 192, 178, 129, 148, 112, 151, 166, 164, 166, 146, 136, 163, 141, 97, 77, 50, 42, 58, 107, 132, 161, 160, 158, 74, 
    99, 276, 284, 275, 260, 222, 182, 161, 196, 206, 122, 101, 102, 160, 208, 223, 195, 149, 125, 118, 91, 54, 35, 22, 30, 68, 111, 140, 163, 163, 151, 69, 
    90, 254, 291, 274, 255, 216, 185, 185, 247, 264, 228, 184, 174, 239, 262, 264, 242, 184, 120, 101, 61, 56, 45, 46, 66, 91, 131, 148, 153, 151, 140, 66, 
    80, 236, 296, 279, 252, 218, 217, 246, 337, 341, 270, 232, 185, 194, 214, 219, 194, 156, 100, 69, 65, 65, 67, 71, 70, 89, 106, 125, 136, 131, 115, 69, 
    50, 192, 258, 270, 260, 248, 270, 297, 371, 365, 281, 159, 132, 133, 141, 142, 127, 120, 101, 87, 70, 68, 74, 81, 85, 88, 97, 110, 108, 105, 99, 60, 
    11, 138, 201, 224, 243, 262, 276, 327, 374, 314, 210, 148, 108, 101, 105, 98, 96, 94, 77, 72, 74, 78, 79, 80, 90, 97, 105, 108, 107, 105, 98, 59, 
    0, 111, 145, 186, 202, 258, 305, 350, 335, 235, 147, 106, 85, 80, 76, 71, 67, 69, 68, 69, 75, 80, 86, 93, 101, 113, 114, 111, 109, 113, 119, 88, 
    0, 103, 101, 121, 164, 239, 303, 337, 285, 180, 116, 89, 86, 81, 75, 75, 75, 75, 75, 78, 80, 88, 98, 107, 111, 108, 103, 105, 111, 134, 152, 100, 
    0, 107, 92, 91, 123, 214, 269, 310, 259, 155, 97, 93, 84, 84, 78, 73, 75, 77, 80, 83, 85, 93, 97, 100, 102, 101, 97, 106, 130, 147, 136, 76, 
    0, 107, 91, 86, 94, 153, 223, 236, 229, 119, 92, 94, 97, 96, 86, 81, 73, 74, 77, 85, 87, 88, 95, 98, 96, 92, 100, 118, 127, 106, 100, 55, 
    1, 115, 92, 82, 87, 103, 146, 164, 152, 94, 77, 78, 88, 99, 94, 88, 84, 89, 95, 94, 91, 91, 86, 83, 91, 107, 128, 135, 125, 106, 94, 37, 
    4, 108, 92, 81, 85, 89, 96, 107, 117, 70, 63, 65, 72, 77, 79, 83, 87, 95, 103, 111, 112, 100, 86, 87, 105, 135, 157, 160, 139, 97, 66, 28, 
    4, 113, 95, 80, 83, 84, 84, 74, 75, 58, 49, 46, 56, 58, 63, 62, 64, 84, 108, 120, 116, 102, 89, 95, 109, 147, 168, 162, 126, 90, 65, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 16, 11, 0, 0, 0, 0, 
    
    -- channel=2
    41, 13, 19, 13, 8, 16, 14, 12, 11, 13, 18, 19, 13, 10, 12, 10, 12, 17, 21, 18, 15, 16, 14, 16, 13, 12, 12, 12, 12, 12, 13, 0, 
    66, 23, 32, 23, 20, 30, 26, 23, 21, 26, 31, 29, 23, 23, 28, 29, 30, 33, 31, 26, 25, 26, 29, 32, 29, 29, 20, 20, 23, 23, 21, 0, 
    64, 21, 34, 28, 27, 31, 26, 23, 22, 27, 41, 29, 5, 16, 32, 35, 36, 27, 25, 33, 23, 16, 13, 25, 30, 32, 30, 25, 23, 22, 20, 0, 
    69, 29, 34, 27, 30, 33, 27, 21, 25, 34, 71, 24, 0, 3, 33, 27, 20, 24, 46, 34, 12, 0, 0, 1, 11, 28, 22, 28, 27, 21, 17, 0, 
    76, 32, 33, 30, 27, 32, 27, 21, 26, 36, 80, 13, 0, 0, 19, 21, 24, 31, 52, 32, 2, 0, 0, 0, 0, 0, 10, 35, 37, 20, 14, 0, 
    79, 14, 19, 49, 34, 27, 28, 24, 27, 33, 75, 22, 0, 0, 1, 13, 5, 25, 62, 36, 0, 0, 0, 0, 0, 0, 0, 22, 45, 24, 11, 0, 
    79, 0, 11, 58, 32, 18, 28, 30, 31, 33, 37, 34, 28, 0, 0, 7, 7, 10, 49, 40, 0, 0, 0, 0, 0, 0, 0, 12, 48, 36, 12, 0, 
    72, 0, 5, 65, 8, 6, 32, 37, 39, 20, 16, 47, 42, 0, 0, 0, 1, 0, 27, 46, 0, 0, 0, 0, 0, 0, 0, 0, 37, 55, 22, 0, 
    70, 0, 3, 27, 0, 0, 31, 62, 71, 0, 0, 16, 22, 0, 0, 0, 0, 0, 7, 67, 25, 0, 0, 0, 0, 0, 0, 0, 7, 56, 44, 0, 
    67, 0, 23, 0, 0, 0, 23, 91, 97, 0, 0, 2, 0, 0, 0, 0, 0, 0, 1, 85, 43, 0, 0, 0, 2, 0, 0, 0, 0, 44, 54, 0, 
    66, 0, 18, 0, 0, 0, 4, 88, 111, 3, 0, 0, 0, 0, 0, 0, 0, 0, 26, 114, 16, 0, 0, 0, 3, 3, 0, 0, 0, 11, 45, 0, 
    46, 0, 36, 0, 0, 0, 0, 49, 123, 21, 0, 0, 21, 0, 0, 0, 0, 0, 42, 122, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 7, 0, 
    36, 0, 50, 0, 0, 0, 3, 0, 108, 50, 0, 23, 38, 0, 0, 0, 0, 0, 57, 108, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 
    34, 0, 48, 0, 0, 0, 12, 0, 78, 57, 10, 36, 25, 0, 0, 0, 0, 0, 58, 85, 0, 0, 0, 0, 0, 5, 8, 2, 0, 0, 0, 0, 
    45, 0, 33, 0, 0, 0, 21, 0, 50, 54, 62, 43, 0, 0, 0, 0, 0, 0, 46, 61, 0, 0, 0, 0, 0, 10, 13, 0, 0, 0, 0, 0, 
    63, 0, 16, 0, 0, 0, 25, 0, 1, 46, 97, 15, 0, 0, 0, 0, 0, 0, 39, 48, 0, 0, 0, 0, 0, 15, 7, 0, 0, 0, 7, 0, 
    82, 0, 0, 0, 0, 0, 19, 0, 0, 36, 67, 12, 0, 0, 0, 0, 0, 0, 18, 3, 19, 1, 0, 0, 0, 24, 16, 0, 0, 10, 13, 0, 
    96, 0, 0, 0, 0, 0, 17, 0, 0, 0, 12, 7, 0, 0, 4, 0, 0, 10, 2, 0, 26, 0, 0, 0, 2, 23, 15, 0, 0, 10, 8, 0, 
    109, 0, 0, 0, 0, 0, 8, 13, 0, 0, 0, 8, 16, 0, 37, 0, 0, 14, 0, 0, 3, 0, 0, 0, 28, 25, 22, 19, 7, 10, 12, 0, 
    128, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 31, 29, 36, 42, 0, 0, 0, 0, 0, 0, 0, 0, 10, 44, 24, 28, 30, 9, 14, 22, 0, 
    154, 0, 0, 0, 0, 0, 0, 60, 0, 0, 0, 2, 26, 30, 16, 0, 0, 0, 0, 0, 0, 0, 3, 19, 27, 22, 23, 25, 13, 20, 25, 0, 
    180, 3, 0, 0, 0, 0, 14, 83, 0, 0, 0, 0, 7, 17, 0, 0, 0, 0, 0, 0, 1, 1, 0, 4, 1, 0, 3, 0, 0, 0, 0, 0, 
    175, 11, 0, 0, 0, 0, 34, 69, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    141, 1, 0, 0, 0, 0, 58, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    100, 0, 0, 2, 0, 0, 57, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    78, 0, 0, 7, 0, 42, 52, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    79, 0, 0, 0, 0, 72, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    82, 0, 0, 0, 0, 67, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    82, 0, 0, 0, 0, 23, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    79, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    83, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    163, 153, 154, 144, 139, 140, 144, 142, 145, 146, 144, 134, 138, 151, 155, 160, 158, 151, 147, 149, 143, 142, 142, 139, 137, 126, 123, 132, 139, 137, 132, 105, 
    165, 155, 154, 144, 140, 145, 144, 144, 145, 143, 126, 104, 125, 154, 155, 150, 144, 133, 143, 137, 134, 127, 139, 149, 144, 150, 139, 134, 137, 135, 129, 101, 
    163, 147, 144, 141, 137, 145, 145, 146, 147, 145, 118, 57, 80, 128, 144, 136, 143, 152, 124, 101, 70, 57, 66, 90, 122, 130, 158, 150, 138, 132, 132, 101, 
    156, 139, 141, 142, 147, 151, 156, 152, 154, 153, 142, 126, 88, 120, 149, 159, 150, 144, 112, 63, 35, 28, 25, 38, 42, 77, 118, 153, 147, 131, 130, 105, 
    153, 132, 176, 179, 158, 152, 153, 151, 150, 159, 175, 201, 188, 140, 134, 141, 123, 89, 75, 53, 43, 53, 62, 49, 47, 62, 89, 138, 153, 131, 119, 98, 
    125, 113, 147, 197, 178, 154, 152, 150, 143, 147, 156, 155, 133, 91, 58, 48, 51, 55, 77, 75, 46, 58, 82, 79, 74, 69, 81, 93, 140, 147, 128, 101, 
    74, 49, 68, 84, 139, 157, 155, 150, 138, 122, 138, 114, 80, 55, 41, 52, 62, 63, 81, 120, 92, 54, 66, 96, 95, 83, 67, 84, 117, 150, 137, 101, 
    60, 0, 16, 33, 70, 138, 152, 138, 77, 39, 24, 63, 46, 48, 53, 67, 81, 86, 99, 119, 123, 78, 50, 70, 91, 76, 54, 56, 93, 150, 157, 101, 
    74, 23, 0, 28, 78, 127, 145, 135, 48, 0, 0, 0, 38, 50, 61, 46, 71, 77, 99, 89, 64, 58, 40, 44, 58, 59, 59, 50, 59, 111, 167, 128, 
    84, 50, 48, 34, 87, 126, 138, 133, 153, 68, 48, 39, 49, 31, 48, 57, 46, 72, 77, 57, 25, 30, 51, 59, 70, 69, 54, 60, 50, 67, 115, 135, 
    77, 55, 74, 65, 92, 114, 121, 121, 165, 166, 113, 92, 58, 27, 29, 60, 49, 35, 60, 53, 44, 47, 83, 78, 83, 85, 76, 53, 40, 39, 71, 100, 
    78, 50, 59, 67, 119, 140, 130, 107, 101, 129, 125, 96, 88, 41, 21, 40, 50, 33, 32, 68, 70, 81, 83, 81, 76, 89, 96, 66, 46, 42, 60, 73, 
    73, 33, 41, 53, 105, 166, 153, 117, 99, 120, 104, 58, 56, 85, 57, 38, 48, 63, 60, 72, 74, 75, 61, 60, 71, 73, 79, 65, 42, 56, 80, 68, 
    68, 21, 46, 49, 54, 120, 147, 124, 98, 104, 95, 40, 26, 106, 110, 89, 69, 61, 77, 97, 84, 62, 69, 58, 57, 58, 50, 60, 66, 85, 100, 88, 
    66, 19, 42, 39, 20, 65, 111, 100, 79, 104, 72, 79, 66, 53, 110, 111, 107, 84, 79, 94, 106, 78, 63, 83, 89, 86, 78, 85, 106, 105, 109, 91, 
    63, 15, 35, 37, 14, 34, 96, 66, 79, 99, 138, 155, 178, 143, 110, 108, 99, 86, 78, 130, 146, 104, 62, 65, 72, 93, 104, 102, 111, 110, 111, 91, 
    72, 11, 30, 49, 33, 25, 74, 83, 52, 60, 116, 155, 134, 119, 88, 66, 72, 85, 84, 107, 137, 157, 128, 102, 115, 103, 114, 106, 93, 108, 121, 100, 
    98, 35, 35, 51, 43, 21, 49, 89, 75, 45, 50, 109, 96, 65, 44, 15, 28, 93, 99, 52, 35, 82, 130, 117, 77, 63, 75, 93, 99, 118, 133, 110, 
    123, 60, 48, 58, 50, 31, 37, 65, 54, 79, 62, 48, 104, 68, 44, 20, 2, 58, 135, 118, 104, 92, 95, 94, 60, 63, 73, 100, 120, 137, 138, 109, 
    133, 76, 52, 61, 56, 47, 46, 21, 0, 0, 62, 49, 30, 25, 15, 14, 1, 14, 79, 149, 148, 122, 74, 44, 54, 66, 105, 121, 125, 127, 129, 99, 
    113, 83, 48, 58, 58, 55, 53, 19, 0, 0, 0, 0, 0, 8, 42, 64, 46, 35, 45, 44, 52, 41, 21, 0, 0, 30, 74, 96, 104, 98, 93, 73, 
    91, 105, 62, 49, 43, 23, 3, 9, 22, 27, 28, 41, 109, 140, 154, 164, 135, 105, 88, 46, 9, 5, 15, 26, 25, 27, 36, 47, 45, 37, 31, 30, 
    74, 132, 137, 77, 46, 42, 8, 21, 52, 118, 127, 130, 113, 111, 116, 112, 96, 70, 56, 48, 38, 35, 32, 32, 30, 20, 18, 26, 29, 24, 20, 19, 
    32, 80, 135, 137, 94, 75, 67, 54, 94, 119, 90, 52, 27, 20, 21, 26, 28, 35, 39, 36, 35, 33, 27, 22, 10, 9, 9, 10, 12, 11, 0, 0, 
    9, 11, 57, 110, 125, 70, 52, 61, 105, 91, 67, 24, 22, 27, 29, 34, 36, 36, 30, 26, 21, 15, 10, 5, 13, 19, 28, 27, 13, 0, 0, 0, 
    21, 12, 28, 61, 95, 105, 66, 69, 77, 59, 30, 31, 23, 29, 35, 31, 26, 22, 19, 17, 13, 16, 17, 13, 22, 38, 48, 32, 11, 6, 25, 36, 
    24, 16, 16, 23, 47, 102, 148, 88, 68, 46, 25, 26, 26, 16, 20, 31, 30, 26, 19, 16, 20, 21, 35, 42, 35, 27, 15, 1, 13, 40, 73, 66, 
    11, 10, 16, 10, 24, 72, 161, 171, 80, 73, 53, 38, 30, 18, 11, 15, 21, 20, 20, 19, 20, 22, 26, 36, 32, 11, 0, 0, 12, 47, 63, 57, 
    14, 0, 14, 13, 13, 40, 92, 142, 102, 64, 67, 65, 63, 56, 41, 24, 13, 6, 2, 1, 8, 20, 27, 27, 16, 0, 0, 0, 0, 13, 13, 48, 
    29, 14, 11, 16, 16, 24, 38, 51, 58, 41, 42, 48, 59, 69, 75, 71, 55, 41, 24, 9, 5, 13, 20, 21, 12, 3, 0, 0, 13, 21, 24, 31, 
    108, 100, 87, 90, 96, 100, 101, 101, 98, 92, 89, 93, 91, 96, 101, 117, 129, 128, 125, 123, 113, 102, 98, 97, 114, 128, 139, 130, 105, 93, 90, 76, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 3, 13, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 68, 12, 0, 0, 0, 0, 0, 10, 37, 52, 48, 26, 15, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 80, 27, 0, 0, 0, 0, 2, 25, 67, 86, 85, 65, 38, 23, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 38, 16, 11, 9, 1, 0, 34, 91, 104, 94, 75, 62, 52, 22, 0, 0, 0, 0, 0, 
    0, 40, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 39, 51, 24, 8, 15, 6, 35, 96, 114, 87, 61, 61, 60, 37, 0, 0, 0, 0, 0, 
    0, 92, 47, 0, 0, 0, 0, 0, 0, 0, 7, 0, 19, 64, 82, 48, 25, 34, 16, 19, 74, 116, 85, 49, 47, 50, 36, 10, 0, 0, 0, 2, 
    0, 141, 82, 23, 42, 8, 0, 0, 12, 85, 103, 64, 56, 105, 107, 67, 36, 41, 27, 0, 42, 115, 101, 63, 44, 37, 37, 22, 0, 0, 0, 0, 
    0, 180, 98, 88, 111, 37, 0, 0, 27, 159, 198, 125, 103, 143, 124, 76, 48, 33, 29, 0, 30, 121, 121, 92, 44, 32, 46, 37, 13, 0, 0, 0, 
    0, 184, 115, 133, 148, 66, 0, 0, 17, 160, 243, 181, 135, 161, 132, 85, 57, 45, 22, 0, 63, 150, 130, 107, 47, 36, 48, 51, 41, 0, 0, 0, 
    0, 187, 97, 156, 169, 76, 0, 0, 0, 112, 208, 157, 116, 169, 154, 95, 74, 63, 33, 0, 104, 176, 138, 106, 44, 34, 50, 51, 50, 32, 0, 0, 
    0, 195, 88, 160, 176, 69, 1, 4, 0, 35, 149, 112, 107, 172, 193, 115, 80, 87, 42, 0, 135, 192, 133, 90, 39, 28, 36, 49, 60, 51, 18, 0, 
    0, 197, 89, 177, 180, 61, 0, 4, 0, 4, 97, 91, 113, 173, 197, 133, 96, 102, 53, 18, 150, 183, 127, 89, 55, 37, 36, 48, 66, 59, 25, 1, 
    0, 200, 107, 200, 192, 67, 2, 20, 4, 0, 66, 103, 181, 204, 173, 132, 104, 94, 49, 29, 138, 165, 123, 81, 48, 35, 37, 50, 69, 54, 6, 0, 
    0, 214, 138, 205, 210, 108, 24, 54, 27, 4, 21, 107, 201, 180, 124, 90, 89, 85, 36, 14, 110, 139, 117, 92, 56, 31, 46, 54, 56, 29, 0, 0, 
    0, 233, 170, 203, 224, 151, 55, 74, 73, 22, 20, 92, 155, 147, 84, 63, 69, 61, 31, 21, 53, 74, 108, 84, 30, 10, 27, 42, 36, 7, 0, 8, 
    0, 244, 196, 204, 231, 184, 79, 90, 116, 65, 33, 77, 75, 92, 67, 59, 80, 53, 45, 52, 41, 45, 82, 60, 23, 0, 7, 12, 10, 0, 0, 8, 
    0, 233, 207, 202, 223, 202, 102, 76, 133, 111, 80, 65, 30, 71, 57, 90, 117, 56, 48, 80, 50, 38, 54, 33, 3, 0, 3, 0, 4, 0, 0, 8, 
    0, 200, 209, 196, 206, 209, 134, 88, 138, 148, 107, 45, 21, 71, 77, 145, 168, 81, 41, 52, 53, 52, 24, 1, 0, 5, 4, 0, 7, 2, 0, 15, 
    0, 164, 212, 188, 192, 204, 141, 87, 173, 207, 167, 103, 71, 110, 132, 190, 212, 143, 64, 52, 41, 45, 29, 17, 24, 38, 40, 37, 49, 41, 30, 59, 
    0, 145, 225, 194, 193, 204, 138, 87, 213, 284, 215, 154, 110, 120, 159, 190, 196, 162, 98, 60, 45, 41, 46, 54, 63, 77, 74, 81, 93, 88, 78, 103, 
    0, 129, 215, 201, 205, 213, 141, 110, 231, 300, 277, 169, 119, 128, 149, 152, 158, 148, 113, 88, 70, 69, 74, 90, 105, 111, 112, 116, 119, 119, 114, 139, 
    0, 114, 173, 178, 200, 206, 134, 156, 264, 294, 257, 177, 116, 114, 122, 112, 117, 116, 95, 87, 90, 97, 101, 106, 117, 123, 128, 125, 130, 132, 129, 156, 
    0, 124, 123, 139, 178, 182, 142, 206, 292, 273, 195, 130, 103, 103, 102, 92, 88, 93, 91, 88, 95, 104, 111, 116, 121, 132, 137, 135, 139, 143, 142, 178, 
    0, 145, 110, 98, 143, 148, 142, 243, 301, 225, 140, 113, 111, 111, 106, 98, 95, 95, 94, 95, 100, 110, 121, 125, 131, 136, 135, 136, 142, 153, 159, 201, 
    0, 161, 130, 106, 108, 115, 144, 273, 289, 174, 108, 114, 114, 116, 107, 99, 99, 99, 102, 105, 109, 119, 124, 131, 139, 141, 134, 132, 147, 166, 166, 197, 
    0, 163, 140, 126, 110, 87, 131, 249, 257, 129, 107, 111, 119, 123, 110, 105, 102, 102, 107, 114, 119, 124, 126, 133, 139, 136, 131, 134, 154, 167, 155, 164, 
    0, 167, 142, 133, 130, 97, 94, 187, 194, 104, 97, 98, 107, 121, 120, 114, 109, 111, 118, 123, 124, 128, 123, 121, 125, 131, 139, 157, 176, 176, 137, 128, 
    0, 169, 141, 133, 136, 121, 93, 121, 144, 90, 81, 83, 93, 102, 110, 111, 107, 112, 121, 132, 137, 133, 123, 116, 115, 130, 158, 190, 196, 169, 113, 114, 
    0, 172, 141, 127, 131, 124, 110, 93, 99, 88, 72, 71, 81, 83, 91, 87, 84, 98, 116, 133, 144, 135, 119, 111, 106, 131, 172, 204, 194, 156, 117, 119, 
    0, 66, 50, 39, 43, 38, 34, 24, 20, 20, 8, 8, 12, 11, 12, 7, 7, 16, 28, 44, 58, 50, 36, 26, 23, 40, 70, 98, 90, 56, 36, 48, 
    
    -- channel=5
    66, 97, 98, 97, 95, 97, 95, 97, 96, 96, 96, 93, 97, 102, 102, 104, 104, 100, 98, 94, 89, 86, 84, 86, 85, 83, 79, 79, 80, 78, 74, 30, 
    145, 165, 165, 158, 158, 167, 165, 165, 162, 165, 160, 154, 159, 170, 173, 171, 167, 160, 154, 147, 143, 136, 138, 141, 138, 143, 139, 137, 136, 132, 123, 40, 
    142, 165, 167, 158, 157, 164, 168, 166, 163, 164, 168, 162, 149, 159, 166, 162, 157, 150, 138, 142, 122, 110, 100, 108, 119, 123, 140, 143, 138, 134, 129, 44, 
    140, 161, 165, 155, 160, 167, 173, 168, 169, 172, 189, 184, 150, 156, 155, 150, 138, 129, 134, 111, 101, 91, 90, 85, 82, 105, 105, 130, 141, 138, 130, 48, 
    136, 149, 163, 167, 164, 170, 170, 169, 167, 177, 210, 193, 195, 164, 139, 129, 126, 95, 94, 109, 119, 107, 94, 87, 89, 77, 97, 117, 136, 139, 131, 43, 
    129, 132, 132, 170, 176, 170, 168, 167, 167, 176, 229, 190, 150, 136, 112, 83, 58, 70, 111, 140, 137, 122, 116, 110, 95, 79, 83, 88, 118, 134, 133, 44, 
    122, 89, 102, 123, 156, 170, 171, 168, 167, 166, 174, 159, 140, 110, 79, 76, 73, 90, 122, 152, 159, 135, 114, 115, 105, 82, 56, 80, 103, 125, 136, 44, 
    123, 53, 71, 129, 141, 164, 173, 169, 162, 155, 136, 147, 143, 121, 98, 94, 95, 99, 128, 152, 165, 142, 116, 108, 102, 82, 56, 47, 86, 118, 136, 45, 
    132, 89, 86, 127, 162, 161, 168, 178, 188, 147, 125, 118, 156, 141, 115, 101, 93, 80, 105, 157, 148, 127, 120, 100, 84, 74, 66, 49, 60, 92, 128, 56, 
    147, 110, 165, 156, 163, 168, 164, 184, 223, 188, 167, 185, 175, 144, 105, 99, 81, 80, 70, 135, 158, 136, 114, 92, 98, 92, 72, 52, 48, 79, 101, 42, 
    161, 143, 174, 201, 171, 165, 153, 198, 230, 268, 199, 196, 173, 151, 109, 98, 99, 52, 77, 153, 168, 163, 131, 108, 103, 102, 102, 64, 37, 54, 87, 18, 
    145, 163, 192, 198, 168, 176, 149, 185, 218, 209, 182, 193, 204, 165, 140, 103, 101, 62, 90, 183, 189, 191, 130, 106, 103, 103, 99, 88, 56, 52, 69, 15, 
    138, 159, 194, 184, 158, 182, 163, 132, 180, 178, 177, 199, 205, 189, 158, 131, 112, 70, 135, 206, 201, 168, 119, 94, 96, 105, 105, 102, 73, 71, 69, 20, 
    135, 159, 198, 177, 150, 147, 166, 127, 158, 157, 171, 202, 232, 199, 183, 166, 138, 76, 151, 208, 191, 156, 123, 93, 84, 97, 99, 104, 99, 93, 86, 34, 
    140, 179, 203, 158, 128, 131, 159, 128, 149, 144, 185, 227, 239, 183, 168, 149, 145, 110, 150, 193, 190, 157, 109, 104, 100, 100, 121, 125, 116, 115, 116, 35, 
    154, 187, 206, 169, 116, 124, 148, 131, 140, 142, 231, 225, 226, 212, 156, 158, 129, 103, 160, 199, 172, 163, 138, 91, 87, 99, 120, 132, 120, 124, 126, 43, 
    176, 193, 204, 190, 127, 131, 138, 156, 139, 160, 193, 236, 183, 150, 144, 127, 116, 118, 155, 151, 180, 171, 122, 88, 99, 104, 115, 127, 115, 124, 136, 53, 
    195, 208, 209, 208, 144, 136, 136, 146, 137, 159, 144, 155, 152, 115, 130, 113, 105, 121, 158, 152, 142, 108, 112, 98, 67, 88, 98, 112, 130, 145, 153, 56, 
    210, 220, 217, 219, 163, 126, 146, 149, 139, 156, 122, 98, 117, 128, 157, 129, 110, 128, 141, 122, 131, 121, 78, 50, 59, 72, 106, 125, 147, 158, 156, 51, 
    214, 232, 218, 218, 185, 129, 144, 156, 149, 105, 98, 142, 114, 158, 176, 139, 124, 131, 118, 135, 119, 97, 62, 36, 66, 77, 141, 161, 164, 160, 157, 55, 
    207, 229, 218, 219, 193, 131, 145, 182, 180, 155, 65, 106, 120, 149, 194, 180, 125, 122, 115, 92, 76, 45, 41, 44, 56, 82, 118, 139, 141, 135, 124, 42, 
    195, 217, 219, 215, 191, 139, 164, 223, 197, 189, 158, 113, 162, 208, 225, 205, 154, 120, 102, 81, 47, 39, 39, 61, 75, 88, 113, 129, 114, 112, 108, 26, 
    172, 203, 229, 221, 188, 144, 198, 275, 296, 227, 180, 198, 180, 181, 181, 162, 133, 109, 71, 58, 63, 76, 81, 83, 84, 90, 94, 99, 98, 94, 87, 11, 
    140, 170, 194, 226, 196, 172, 270, 307, 303, 232, 170, 117, 108, 100, 93, 94, 73, 69, 75, 77, 79, 82, 86, 88, 86, 87, 93, 98, 93, 89, 87, 11, 
    96, 128, 152, 181, 196, 218, 278, 298, 250, 170, 107, 74, 74, 71, 68, 74, 77, 75, 75, 78, 78, 80, 81, 83, 92, 91, 96, 97, 94, 95, 98, 5, 
    72, 92, 123, 153, 149, 231, 289, 280, 189, 124, 73, 82, 78, 76, 77, 76, 75, 73, 73, 74, 80, 83, 87, 90, 95, 103, 103, 103, 107, 109, 109, 16, 
    78, 83, 91, 115, 127, 213, 303, 246, 144, 97, 81, 82, 87, 76, 70, 73, 75, 75, 76, 81, 85, 86, 95, 107, 106, 98, 94, 106, 107, 115, 132, 33, 
    81, 82, 78, 80, 113, 198, 255, 216, 129, 103, 95, 93, 81, 80, 75, 69, 73, 78, 83, 85, 86, 96, 97, 94, 92, 90, 91, 100, 110, 122, 119, 16, 
    83, 79, 76, 77, 84, 160, 199, 146, 137, 92, 89, 98, 95, 91, 84, 80, 77, 78, 77, 84, 85, 83, 89, 90, 91, 90, 102, 112, 115, 78, 74, 0, 
    82, 92, 80, 77, 76, 100, 148, 95, 83, 82, 79, 84, 88, 94, 92, 90, 86, 92, 98, 95, 86, 80, 82, 85, 94, 113, 131, 118, 88, 61, 80, 0, 
    86, 87, 82, 75, 80, 77, 89, 85, 65, 63, 67, 73, 78, 79, 73, 83, 98, 106, 110, 108, 100, 92, 81, 87, 116, 144, 149, 131, 96, 70, 64, 0, 
    58, 93, 94, 85, 84, 85, 81, 80, 70, 63, 64, 61, 65, 65, 71, 73, 76, 91, 109, 115, 107, 96, 89, 103, 120, 151, 154, 133, 99, 80, 61, 14, 
    
    -- channel=6
    58, 50, 53, 60, 56, 51, 57, 56, 57, 53, 54, 55, 54, 56, 58, 59, 59, 56, 52, 53, 53, 50, 51, 50, 56, 54, 53, 52, 54, 54, 53, 93, 
    36, 52, 53, 60, 56, 56, 58, 58, 60, 58, 56, 54, 53, 57, 60, 60, 62, 58, 55, 50, 50, 45, 43, 45, 47, 52, 55, 52, 57, 59, 57, 110, 
    37, 56, 53, 60, 53, 55, 58, 60, 58, 58, 52, 61, 57, 52, 59, 60, 60, 63, 47, 46, 43, 41, 34, 32, 36, 33, 48, 53, 57, 60, 60, 112, 
    34, 57, 55, 58, 56, 53, 59, 60, 58, 53, 27, 82, 68, 50, 53, 59, 51, 48, 36, 42, 38, 43, 40, 36, 31, 29, 30, 43, 53, 59, 58, 115, 
    32, 52, 48, 54, 59, 55, 59, 61, 57, 53, 12, 60, 73, 57, 45, 42, 49, 29, 22, 29, 29, 34, 40, 38, 36, 41, 24, 25, 41, 59, 56, 115, 
    27, 57, 20, 37, 62, 61, 58, 62, 60, 56, 32, 30, 49, 61, 52, 28, 44, 27, 4, 19, 29, 25, 26, 25, 40, 39, 35, 15, 21, 53, 57, 115, 
    31, 67, 15, 12, 51, 61, 58, 60, 63, 57, 53, 37, 37, 61, 59, 34, 39, 30, 0, 6, 39, 33, 16, 21, 33, 39, 39, 25, 5, 34, 56, 116, 
    50, 66, 19, 24, 42, 55, 56, 55, 55, 71, 47, 37, 38, 54, 52, 28, 27, 33, 5, 0, 29, 50, 29, 19, 26, 42, 37, 35, 5, 13, 53, 118, 
    50, 65, 3, 32, 52, 51, 54, 38, 48, 86, 62, 21, 37, 42, 50, 27, 23, 28, 17, 0, 12, 43, 48, 30, 22, 35, 41, 44, 22, 0, 35, 122, 
    38, 35, 10, 19, 60, 51, 59, 0, 29, 67, 80, 14, 35, 39, 40, 43, 22, 38, 8, 0, 23, 27, 55, 40, 21, 34, 34, 47, 44, 4, 8, 110, 
    44, 0, 1, 19, 63, 53, 71, 0, 0, 30, 55, 16, 27, 54, 29, 45, 32, 50, 0, 0, 40, 23, 53, 36, 18, 28, 37, 38, 49, 27, 13, 83, 
    53, 0, 0, 19, 56, 54, 72, 45, 0, 5, 33, 1, 12, 65, 42, 31, 40, 64, 0, 0, 34, 31, 44, 35, 19, 14, 35, 33, 45, 34, 35, 73, 
    57, 0, 0, 28, 29, 46, 66, 80, 0, 2, 21, 3, 0, 57, 58, 33, 29, 67, 0, 0, 28, 40, 40, 33, 24, 13, 20, 30, 38, 32, 46, 83, 
    56, 0, 0, 45, 23, 23, 56, 87, 5, 4, 5, 24, 0, 29, 46, 41, 34, 47, 0, 0, 33, 35, 44, 37, 23, 21, 13, 24, 37, 31, 38, 100, 
    49, 0, 0, 47, 49, 4, 43, 82, 26, 10, 0, 24, 42, 8, 23, 30, 39, 45, 0, 0, 31, 39, 36, 38, 19, 23, 20, 20, 41, 34, 37, 111, 
    36, 0, 0, 35, 70, 0, 30, 66, 52, 0, 0, 0, 50, 33, 16, 20, 27, 44, 0, 1, 15, 42, 39, 37, 15, 8, 19, 21, 34, 34, 44, 112, 
    28, 7, 0, 17, 75, 6, 2, 53, 69, 0, 0, 0, 14, 39, 13, 28, 17, 27, 20, 14, 0, 30, 54, 37, 23, 6, 11, 28, 28, 36, 45, 117, 
    15, 14, 0, 3, 64, 36, 0, 24, 62, 37, 12, 0, 27, 30, 20, 47, 14, 6, 48, 42, 9, 18, 38, 38, 19, 20, 7, 34, 41, 47, 53, 128, 
    0, 18, 0, 0, 44, 57, 0, 0, 31, 51, 54, 0, 35, 17, 17, 64, 32, 0, 34, 50, 51, 29, 23, 39, 13, 33, 14, 30, 42, 45, 51, 122, 
    0, 21, 3, 0, 29, 58, 0, 0, 32, 20, 60, 5, 11, 3, 10, 53, 58, 2, 6, 26, 36, 41, 32, 20, 10, 13, 17, 32, 44, 42, 50, 121, 
    0, 23, 9, 0, 25, 49, 0, 0, 57, 47, 25, 25, 4, 2, 6, 33, 59, 36, 24, 17, 16, 25, 32, 17, 9, 0, 4, 16, 34, 29, 30, 110, 
    0, 14, 14, 3, 28, 45, 0, 0, 22, 74, 54, 13, 0, 0, 0, 12, 35, 28, 40, 33, 25, 15, 16, 17, 11, 0, 0, 12, 29, 27, 25, 95, 
    0, 0, 10, 5, 26, 40, 0, 0, 0, 41, 43, 4, 0, 0, 0, 0, 7, 8, 16, 22, 18, 12, 3, 1, 1, 1, 0, 0, 9, 8, 8, 70, 
    0, 0, 0, 0, 24, 5, 0, 0, 14, 29, 15, 8, 0, 0, 0, 0, 0, 5, 6, 4, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 
    0, 0, 0, 0, 17, 0, 0, 2, 40, 20, 23, 9, 5, 6, 4, 4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 80, 
    1, 0, 0, 0, 0, 0, 0, 31, 41, 16, 8, 2, 2, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 82, 
    0, 0, 0, 0, 0, 0, 0, 54, 36, 21, 0, 0, 4, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 70, 
    0, 0, 0, 0, 0, 0, 0, 63, 26, 15, 3, 0, 4, 5, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 65, 
    0, 0, 0, 0, 0, 0, 0, 29, 23, 3, 0, 0, 0, 3, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 58, 
    0, 0, 0, 0, 0, 0, 0, 0, 21, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 2, 3, 0, 45, 
    0, 4, 0, 0, 0, 0, 0, 0, 11, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 6, 0, 0, 0, 0, 0, 0, 6, 4, 0, 6, 43, 
    0, 5, 2, 0, 0, 1, 6, 8, 12, 13, 6, 8, 7, 9, 6, 0, 0, 0, 0, 0, 5, 5, 5, 0, 0, 0, 0, 6, 12, 3, 9, 36, 
    
    -- channel=7
    109, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    142, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    138, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    135, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 23, 13, 12, 5, 6, 12, 12, 10, 0, 0, 0, 0, 0, 
    134, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 40, 57, 29, 22, 5, 9, 14, 9, 0, 22, 18, 0, 0, 0, 
    141, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 19, 71, 81, 30, 7, 11, 17, 18, 1, 0, 21, 45, 17, 0, 0, 
    153, 0, 0, 52, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 23, 58, 93, 35, 0, 0, 23, 22, 0, 1, 19, 48, 46, 0, 0, 
    177, 0, 0, 75, 21, 0, 0, 0, 0, 0, 0, 0, 23, 2, 0, 0, 35, 24, 32, 79, 62, 0, 0, 15, 22, 12, 6, 13, 32, 65, 18, 0, 
    217, 0, 0, 86, 0, 0, 0, 0, 11, 0, 0, 0, 28, 0, 0, 0, 28, 21, 26, 70, 88, 4, 0, 0, 16, 26, 14, 10, 7, 51, 56, 0, 
    233, 0, 25, 67, 0, 0, 0, 0, 77, 0, 0, 0, 26, 0, 0, 0, 10, 20, 18, 89, 103, 4, 0, 0, 12, 35, 12, 7, 0, 26, 66, 0, 
    247, 0, 72, 52, 0, 0, 0, 0, 107, 61, 0, 0, 27, 0, 0, 0, 0, 7, 16, 131, 98, 0, 0, 0, 12, 46, 17, 8, 1, 12, 50, 8, 
    247, 0, 102, 54, 0, 0, 0, 0, 61, 110, 0, 0, 51, 0, 0, 0, 5, 0, 4, 159, 80, 0, 0, 0, 21, 44, 28, 11, 16, 11, 30, 0, 
    250, 0, 114, 44, 0, 0, 0, 0, 0, 115, 0, 4, 62, 12, 0, 0, 4, 0, 0, 165, 53, 0, 0, 0, 23, 37, 45, 32, 24, 12, 18, 0, 
    252, 0, 117, 26, 0, 0, 0, 0, 0, 90, 24, 41, 27, 5, 0, 0, 0, 0, 12, 153, 34, 0, 0, 0, 18, 36, 44, 47, 25, 1, 9, 0, 
    259, 0, 104, 13, 0, 0, 25, 0, 0, 64, 56, 93, 0, 0, 0, 0, 0, 0, 23, 129, 37, 0, 0, 0, 13, 47, 45, 44, 18, 0, 5, 0, 
    268, 0, 80, 19, 0, 0, 53, 0, 0, 29, 77, 77, 0, 0, 0, 12, 6, 1, 29, 95, 22, 0, 0, 0, 8, 52, 49, 30, 13, 0, 2, 0, 
    284, 0, 54, 30, 0, 0, 72, 21, 0, 0, 83, 51, 0, 0, 0, 22, 12, 29, 12, 20, 10, 41, 0, 0, 8, 50, 61, 36, 7, 0, 0, 0, 
    297, 0, 35, 39, 0, 0, 42, 71, 0, 0, 30, 25, 38, 3, 10, 25, 0, 44, 39, 0, 0, 42, 0, 0, 19, 58, 61, 50, 5, 0, 0, 0, 
    297, 0, 20, 37, 0, 0, 2, 87, 9, 0, 0, 0, 70, 4, 44, 31, 0, 32, 63, 0, 0, 2, 0, 11, 37, 71, 37, 37, 0, 0, 0, 0, 
    283, 18, 6, 27, 8, 0, 0, 99, 28, 0, 0, 0, 84, 36, 72, 22, 0, 0, 45, 1, 1, 0, 0, 39, 57, 76, 34, 20, 0, 0, 0, 0, 
    261, 65, 0, 16, 9, 0, 0, 124, 81, 0, 0, 12, 66, 55, 67, 8, 0, 0, 3, 2, 20, 31, 46, 54, 74, 65, 47, 26, 0, 0, 0, 0, 
    246, 118, 0, 10, 10, 0, 8, 146, 78, 0, 0, 0, 39, 58, 45, 12, 0, 0, 4, 6, 36, 56, 65, 66, 71, 65, 78, 62, 41, 29, 46, 5, 
    227, 149, 35, 25, 17, 0, 23, 144, 46, 0, 0, 0, 50, 69, 54, 50, 41, 28, 40, 38, 61, 71, 77, 80, 79, 81, 87, 86, 77, 66, 76, 26, 
    213, 132, 95, 78, 27, 0, 63, 109, 0, 0, 0, 9, 66, 75, 71, 73, 72, 64, 70, 75, 84, 84, 84, 89, 92, 95, 86, 86, 81, 75, 84, 32, 
    211, 102, 111, 121, 71, 21, 108, 63, 0, 0, 0, 50, 72, 72, 69, 73, 78, 77, 81, 85, 91, 93, 89, 95, 97, 93, 81, 80, 84, 88, 98, 31, 
    214, 74, 95, 117, 103, 78, 131, 19, 0, 0, 52, 76, 75, 73, 75, 78, 76, 77, 81, 86, 90, 95, 95, 91, 90, 83, 81, 88, 104, 100, 96, 20, 
    220, 70, 84, 100, 102, 135, 159, 0, 0, 0, 69, 82, 80, 66, 76, 81, 79, 79, 82, 87, 89, 89, 98, 97, 87, 80, 91, 109, 117, 93, 84, 21, 
    221, 76, 86, 93, 97, 129, 178, 22, 0, 34, 72, 82, 85, 67, 72, 76, 80, 85, 89, 87, 91, 90, 97, 97, 89, 89, 102, 115, 105, 82, 76, 46, 
    223, 68, 89, 97, 93, 106, 139, 79, 0, 56, 77, 90, 93, 76, 72, 71, 83, 86, 87, 86, 87, 86, 88, 95, 101, 107, 107, 109, 84, 64, 66, 69, 
    228, 63, 84, 102, 90, 93, 100, 93, 30, 64, 84, 97, 91, 87, 84, 77, 85, 87, 89, 85, 75, 74, 82, 92, 110, 120, 110, 75, 51, 55, 71, 62, 
    228, 68, 74, 98, 90, 87, 79, 79, 69, 64, 84, 97, 89, 91, 84, 87, 98, 97, 94, 87, 66, 63, 76, 88, 116, 118, 99, 53, 39, 57, 86, 40, 
    170, 76, 74, 89, 87, 85, 77, 75, 77, 70, 80, 87, 79, 85, 80, 84, 92, 92, 91, 87, 68, 64, 76, 79, 101, 101, 90, 64, 52, 68, 89, 45, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 46, 64, 55, 31, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 38, 60, 68, 62, 50, 33, 17, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 10, 24, 40, 42, 38, 34, 26, 29, 31, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 29, 27, 16, 26, 23, 13, 6, 7, 16, 24, 25, 0, 0, 0, 0, 0, 
    37, 53, 47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 18, 30, 29, 9, 6, 13, 13, 5, 6, 11, 23, 25, 7, 0, 0, 0, 0, 
    66, 96, 83, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 18, 14, 27, 22, 14, 3, 13, 30, 19, 14, 16, 22, 30, 20, 0, 0, 0, 0, 
    79, 124, 114, 52, 0, 0, 0, 0, 0, 28, 36, 5, 15, 14, 16, 12, 23, 20, 19, 19, 32, 43, 30, 23, 21, 27, 32, 35, 14, 0, 0, 0, 
    89, 125, 133, 69, 0, 0, 0, 0, 0, 18, 28, 0, 10, 13, 9, 15, 22, 25, 28, 34, 57, 49, 40, 28, 25, 32, 34, 42, 37, 11, 0, 0, 
    94, 125, 131, 79, 0, 0, 0, 0, 0, 0, 2, 0, 10, 25, 16, 14, 27, 31, 33, 50, 73, 54, 43, 30, 28, 29, 38, 44, 47, 23, 0, 0, 
    93, 119, 122, 96, 0, 0, 0, 0, 0, 0, 0, 0, 22, 49, 37, 25, 28, 40, 39, 64, 76, 63, 46, 38, 40, 34, 42, 48, 43, 9, 0, 0, 
    93, 110, 117, 118, 34, 0, 0, 0, 0, 0, 1, 28, 50, 77, 50, 35, 26, 27, 29, 55, 68, 56, 47, 38, 42, 39, 40, 40, 16, 0, 0, 0, 
    99, 115, 122, 132, 77, 13, 0, 0, 0, 0, 0, 52, 64, 55, 35, 27, 22, 4, 0, 0, 29, 32, 41, 38, 39, 44, 36, 13, 0, 0, 0, 0, 
    109, 136, 140, 144, 113, 66, 25, 0, 0, 0, 0, 37, 48, 17, 12, 14, 21, 0, 0, 0, 0, 7, 21, 23, 20, 30, 23, 0, 0, 0, 0, 0, 
    118, 152, 161, 159, 141, 97, 82, 34, 0, 0, 0, 8, 0, 0, 0, 20, 38, 12, 0, 0, 0, 0, 10, 8, 11, 2, 0, 0, 0, 0, 0, 0, 
    109, 145, 163, 164, 152, 110, 92, 76, 49, 14, 0, 0, 0, 0, 9, 42, 52, 30, 0, 0, 0, 0, 10, 5, 18, 0, 0, 0, 0, 0, 0, 0, 
    88, 119, 141, 145, 141, 118, 106, 111, 92, 67, 25, 0, 11, 21, 37, 76, 64, 30, 7, 0, 1, 18, 18, 34, 43, 0, 0, 0, 0, 0, 0, 0, 
    77, 106, 120, 121, 122, 115, 114, 133, 132, 108, 88, 50, 72, 81, 92, 118, 98, 54, 26, 19, 41, 64, 76, 95, 108, 84, 22, 0, 0, 0, 0, 0, 
    97, 145, 134, 120, 119, 115, 117, 132, 168, 150, 129, 128, 132, 144, 150, 157, 144, 116, 86, 85, 107, 140, 161, 175, 195, 188, 168, 151, 138, 140, 149, 105, 
    141, 221, 179, 150, 138, 125, 115, 125, 165, 179, 171, 178, 182, 193, 189, 198, 201, 191, 184, 182, 200, 224, 238, 256, 273, 284, 292, 288, 281, 284, 291, 188, 
    192, 291, 239, 193, 157, 134, 109, 133, 157, 191, 213, 218, 221, 228, 222, 232, 245, 245, 246, 257, 272, 285, 289, 302, 316, 321, 326, 322, 321, 324, 332, 207, 
    236, 332, 285, 234, 179, 143, 117, 142, 167, 218, 232, 251, 254, 256, 251, 253, 261, 269, 274, 288, 301, 311, 318, 325, 332, 330, 328, 327, 335, 344, 353, 217, 
    264, 363, 311, 263, 214, 157, 145, 160, 197, 228, 255, 275, 276, 277, 269, 266, 266, 274, 283, 295, 312, 325, 335, 339, 340, 337, 335, 346, 363, 371, 372, 232, 
    274, 384, 343, 293, 250, 204, 189, 195, 215, 232, 266, 284, 282, 281, 275, 271, 272, 281, 291, 305, 323, 338, 351, 351, 352, 350, 357, 374, 389, 384, 374, 232, 
    274, 394, 371, 335, 287, 248, 237, 225, 226, 245, 272, 288, 288, 285, 279, 278, 279, 289, 301, 315, 332, 344, 356, 358, 357, 361, 377, 394, 403, 381, 361, 212, 
    271, 395, 384, 363, 328, 274, 264, 251, 237, 257, 277, 286, 293, 293, 286, 285, 285, 295, 307, 318, 333, 341, 346, 349, 352, 365, 384, 406, 410, 377, 343, 199, 
    265, 384, 377, 367, 348, 305, 271, 273, 251, 265, 278, 284, 290, 292, 288, 284, 284, 294, 307, 319, 326, 330, 330, 332, 338, 358, 381, 404, 398, 370, 327, 201, 
    260, 368, 356, 354, 345, 322, 288, 276, 268, 272, 276, 279, 283, 284, 279, 273, 272, 286, 302, 313, 316, 315, 310, 313, 321, 340, 364, 377, 377, 362, 329, 201, 
    177, 237, 224, 225, 223, 214, 197, 183, 182, 181, 181, 183, 183, 182, 177, 172, 172, 181, 193, 204, 205, 199, 196, 195, 202, 213, 230, 239, 240, 231, 221, 136, 
    
    -- channel=10
    89, 61, 67, 61, 56, 61, 61, 59, 55, 55, 60, 60, 62, 64, 59, 56, 51, 50, 55, 56, 54, 52, 52, 55, 52, 48, 43, 41, 37, 32, 28, 0, 
    148, 94, 102, 92, 88, 96, 98, 94, 92, 91, 95, 96, 97, 97, 91, 90, 86, 84, 81, 77, 70, 68, 74, 77, 81, 82, 78, 73, 68, 60, 53, 0, 
    145, 87, 99, 93, 90, 100, 101, 96, 92, 98, 124, 122, 100, 96, 92, 90, 90, 70, 72, 79, 81, 71, 63, 67, 62, 72, 80, 78, 73, 66, 59, 0, 
    147, 89, 97, 94, 90, 99, 99, 93, 92, 106, 184, 171, 111, 94, 96, 78, 55, 54, 78, 102, 109, 100, 91, 73, 73, 70, 76, 81, 81, 70, 62, 0, 
    145, 83, 96, 99, 96, 98, 98, 90, 91, 103, 171, 167, 93, 68, 57, 51, 43, 52, 103, 140, 146, 134, 105, 96, 85, 62, 57, 77, 93, 82, 68, 0, 
    145, 46, 59, 100, 105, 98, 96, 92, 90, 100, 155, 139, 90, 74, 55, 52, 44, 67, 146, 184, 168, 142, 126, 117, 100, 68, 38, 58, 96, 91, 71, 0, 
    148, 40, 41, 105, 118, 99, 92, 95, 92, 88, 95, 105, 116, 96, 58, 69, 81, 85, 150, 206, 182, 134, 117, 120, 103, 54, 29, 40, 86, 101, 80, 0, 
    171, 33, 69, 139, 133, 103, 97, 104, 115, 86, 83, 123, 157, 132, 78, 82, 93, 86, 117, 187, 184, 126, 100, 104, 90, 64, 37, 21, 58, 103, 93, 0, 
    221, 82, 129, 187, 143, 104, 100, 154, 205, 183, 132, 167, 187, 149, 93, 88, 90, 68, 86, 170, 191, 144, 110, 92, 87, 75, 59, 29, 24, 77, 100, 0, 
    235, 138, 207, 228, 144, 105, 90, 185, 282, 246, 176, 204, 207, 148, 110, 83, 86, 54, 68, 183, 220, 182, 119, 85, 100, 95, 74, 38, 12, 47, 86, 0, 
    248, 169, 251, 252, 155, 110, 89, 149, 295, 289, 206, 210, 227, 160, 119, 102, 84, 35, 88, 239, 244, 193, 128, 81, 99, 115, 95, 63, 21, 35, 64, 0, 
    232, 177, 276, 253, 158, 115, 90, 110, 243, 264, 184, 211, 261, 196, 139, 118, 113, 44, 123, 282, 257, 182, 120, 79, 101, 114, 99, 82, 53, 48, 49, 0, 
    227, 180, 291, 231, 138, 120, 102, 56, 167, 225, 193, 226, 300, 240, 156, 138, 132, 60, 156, 306, 249, 162, 104, 78, 88, 103, 112, 107, 86, 75, 55, 0, 
    231, 190, 302, 215, 111, 121, 121, 47, 113, 183, 206, 253, 289, 236, 172, 165, 144, 71, 174, 296, 229, 161, 121, 93, 97, 107, 125, 136, 111, 87, 70, 0, 
    252, 214, 305, 208, 97, 129, 141, 71, 109, 170, 262, 329, 276, 216, 170, 156, 136, 87, 173, 269, 223, 149, 109, 82, 90, 113, 137, 147, 110, 91, 86, 0, 
    280, 230, 303, 236, 113, 135, 163, 107, 86, 167, 257, 292, 222, 157, 156, 147, 120, 90, 177, 235, 201, 165, 131, 87, 89, 118, 129, 125, 102, 92, 95, 0, 
    316, 245, 296, 269, 142, 125, 190, 152, 106, 148, 221, 235, 166, 122, 136, 123, 119, 129, 146, 139, 160, 161, 98, 57, 63, 95, 117, 113, 102, 105, 103, 0, 
    346, 261, 297, 292, 180, 125, 191, 200, 132, 130, 142, 157, 150, 129, 150, 126, 112, 152, 163, 128, 126, 128, 80, 33, 48, 76, 113, 117, 111, 113, 100, 0, 
    358, 270, 291, 296, 213, 123, 178, 205, 163, 155, 96, 119, 137, 142, 200, 160, 100, 158, 160, 112, 112, 93, 42, 22, 61, 87, 127, 136, 122, 111, 94, 0, 
    351, 280, 281, 291, 237, 139, 175, 245, 185, 130, 76, 107, 156, 193, 254, 202, 117, 127, 131, 96, 72, 34, 15, 30, 68, 100, 134, 141, 111, 98, 90, 0, 
    333, 291, 273, 283, 238, 132, 178, 304, 296, 200, 137, 168, 216, 260, 304, 249, 152, 134, 110, 77, 52, 43, 56, 74, 109, 129, 143, 144, 119, 106, 102, 0, 
    315, 314, 275, 281, 239, 150, 234, 375, 359, 268, 186, 181, 219, 258, 265, 225, 150, 109, 91, 70, 70, 85, 93, 113, 126, 141, 158, 157, 134, 126, 124, 0, 
    265, 308, 282, 289, 253, 192, 300, 432, 411, 265, 167, 162, 186, 197, 188, 177, 144, 121, 100, 88, 104, 123, 134, 140, 144, 153, 161, 164, 155, 147, 145, 2, 
    212, 247, 267, 293, 243, 236, 363, 436, 353, 236, 139, 130, 151, 151, 146, 145, 128, 120, 118, 123, 132, 136, 143, 151, 160, 165, 169, 172, 162, 157, 162, 10, 
    180, 198, 229, 273, 246, 285, 406, 398, 256, 142, 106, 123, 131, 128, 122, 124, 126, 125, 125, 132, 143, 147, 151, 164, 176, 178, 176, 175, 172, 183, 199, 22, 
    167, 157, 185, 223, 229, 322, 426, 338, 174, 104, 127, 142, 138, 132, 130, 130, 128, 129, 131, 138, 150, 160, 170, 175, 177, 174, 166, 178, 198, 212, 218, 28, 
    176, 151, 157, 180, 202, 341, 425, 279, 126, 116, 139, 151, 143, 129, 128, 131, 132, 134, 139, 150, 154, 160, 174, 181, 174, 161, 168, 198, 216, 210, 207, 19, 
    177, 156, 151, 155, 180, 291, 381, 220, 110, 130, 147, 158, 152, 141, 135, 131, 130, 139, 147, 153, 159, 164, 171, 169, 161, 162, 184, 203, 205, 173, 172, 10, 
    183, 157, 158, 154, 160, 220, 277, 179, 102, 120, 132, 152, 158, 151, 144, 142, 148, 154, 156, 160, 157, 153, 154, 159, 171, 190, 212, 222, 194, 134, 139, 12, 
    186, 155, 158, 159, 153, 167, 199, 151, 102, 112, 123, 135, 139, 141, 139, 142, 152, 165, 177, 176, 161, 151, 146, 159, 192, 233, 249, 215, 160, 122, 124, 9, 
    189, 155, 153, 155, 153, 143, 142, 131, 106, 97, 112, 121, 126, 123, 115, 125, 146, 166, 183, 182, 162, 149, 141, 164, 210, 252, 249, 197, 146, 125, 121, 1, 
    89, 51, 50, 54, 54, 50, 40, 37, 29, 21, 29, 31, 30, 32, 32, 39, 51, 63, 76, 74, 55, 46, 47, 61, 89, 112, 106, 72, 39, 39, 34, 0, 
    
    -- channel=11
    37, 42, 41, 44, 42, 38, 41, 40, 42, 41, 42, 45, 40, 38, 42, 43, 44, 43, 42, 44, 45, 46, 46, 44, 45, 43, 45, 45, 46, 48, 49, 83, 
    2, 19, 20, 29, 25, 20, 22, 22, 24, 20, 18, 24, 24, 20, 24, 22, 23, 23, 27, 35, 42, 44, 41, 37, 36, 31, 31, 28, 29, 31, 34, 87, 
    4, 20, 17, 25, 20, 18, 19, 21, 23, 20, 7, 9, 16, 18, 23, 22, 24, 36, 39, 34, 31, 32, 35, 39, 42, 42, 39, 30, 28, 30, 32, 86, 
    1, 20, 16, 24, 23, 20, 23, 25, 23, 17, 0, 5, 17, 15, 24, 36, 49, 59, 34, 24, 19, 25, 19, 20, 26, 24, 31, 34, 31, 32, 34, 89, 
    1, 31, 26, 26, 25, 20, 23, 25, 22, 17, 0, 55, 57, 40, 49, 61, 54, 34, 17, 17, 17, 26, 31, 29, 22, 35, 33, 33, 29, 30, 28, 88, 
    5, 53, 47, 37, 27, 19, 20, 23, 20, 16, 0, 33, 50, 39, 33, 28, 38, 22, 2, 4, 14, 29, 36, 27, 33, 45, 39, 29, 25, 33, 31, 89, 
    2, 60, 23, 11, 21, 22, 22, 22, 22, 23, 24, 28, 22, 32, 38, 22, 28, 22, 0, 5, 21, 28, 29, 31, 44, 53, 56, 34, 16, 30, 32, 88, 
    2, 62, 15, 0, 2, 17, 18, 17, 17, 27, 26, 9, 2, 26, 43, 34, 38, 37, 14, 9, 35, 38, 28, 34, 43, 48, 48, 48, 22, 21, 30, 89, 
    13, 45, 0, 0, 6, 12, 18, 0, 0, 0, 0, 0, 4, 30, 44, 31, 33, 48, 35, 0, 13, 36, 30, 24, 29, 41, 43, 47, 32, 20, 34, 94, 
    21, 43, 0, 0, 27, 15, 24, 0, 0, 16, 28, 0, 10, 28, 37, 33, 33, 49, 31, 0, 0, 9, 36, 36, 24, 31, 39, 54, 49, 18, 26, 100, 
    22, 15, 0, 5, 30, 12, 27, 0, 0, 31, 41, 0, 8, 24, 26, 40, 28, 58, 11, 0, 0, 8, 48, 45, 29, 33, 32, 43, 53, 28, 19, 87, 
    39, 5, 0, 14, 38, 17, 30, 5, 0, 24, 43, 8, 0, 26, 17, 27, 26, 53, 0, 0, 15, 22, 52, 43, 27, 30, 41, 39, 48, 34, 31, 71, 
    46, 0, 0, 24, 46, 28, 28, 41, 0, 18, 19, 0, 0, 22, 25, 17, 25, 64, 0, 0, 16, 34, 48, 43, 35, 30, 33, 29, 38, 31, 40, 67, 
    44, 0, 0, 37, 34, 21, 23, 49, 0, 23, 0, 0, 0, 38, 45, 20, 20, 60, 0, 0, 23, 33, 34, 29, 26, 20, 12, 19, 33, 33, 40, 76, 
    35, 0, 0, 41, 39, 5, 12, 43, 1, 4, 0, 0, 0, 15, 33, 35, 41, 47, 0, 0, 24, 31, 47, 53, 37, 30, 15, 19, 41, 34, 25, 82, 
    22, 0, 0, 23, 51, 0, 7, 32, 23, 8, 0, 12, 63, 36, 32, 29, 38, 49, 0, 0, 20, 33, 26, 34, 26, 26, 29, 32, 45, 27, 20, 86, 
    6, 0, 0, 8, 62, 12, 7, 19, 26, 0, 5, 17, 52, 54, 26, 31, 30, 27, 0, 35, 38, 45, 56, 61, 46, 35, 34, 31, 24, 17, 22, 91, 
    0, 0, 0, 0, 52, 23, 0, 22, 34, 0, 26, 23, 23, 25, 2, 24, 23, 15, 14, 9, 0, 36, 70, 61, 44, 31, 17, 20, 9, 12, 21, 92, 
    0, 6, 0, 0, 36, 42, 0, 18, 37, 20, 30, 3, 34, 20, 0, 26, 25, 5, 31, 31, 23, 36, 55, 60, 27, 25, 0, 8, 16, 19, 26, 97, 
    0, 8, 0, 0, 22, 48, 0, 0, 11, 38, 72, 8, 24, 0, 0, 27, 35, 3, 33, 55, 75, 72, 57, 51, 30, 40, 10, 15, 29, 31, 34, 100, 
    0, 9, 0, 0, 20, 58, 4, 0, 0, 0, 1, 0, 0, 0, 0, 9, 39, 16, 14, 37, 52, 51, 35, 14, 12, 13, 11, 26, 39, 35, 41, 109, 
    0, 5, 1, 0, 19, 43, 0, 0, 0, 14, 0, 7, 10, 11, 24, 43, 70, 65, 54, 35, 29, 24, 29, 26, 24, 21, 16, 16, 28, 25, 26, 97, 
    0, 15, 12, 0, 13, 21, 0, 0, 0, 45, 80, 47, 34, 40, 43, 47, 60, 48, 45, 43, 38, 28, 24, 28, 31, 25, 22, 23, 29, 26, 28, 102, 
    1, 13, 24, 7, 26, 17, 0, 0, 0, 57, 67, 41, 21, 21, 23, 20, 34, 37, 32, 31, 32, 31, 29, 26, 23, 24, 20, 20, 26, 29, 30, 105, 
    22, 2, 0, 7, 32, 0, 0, 0, 48, 71, 60, 36, 29, 31, 33, 31, 34, 35, 32, 28, 27, 27, 24, 21, 16, 21, 22, 22, 24, 18, 7, 101, 
    43, 27, 6, 2, 28, 0, 0, 10, 70, 53, 42, 28, 30, 34, 33, 30, 31, 31, 29, 27, 25, 23, 19, 17, 24, 29, 32, 28, 20, 7, 9, 120, 
    43, 37, 24, 10, 7, 0, 0, 42, 61, 41, 30, 29, 32, 31, 33, 33, 31, 29, 29, 25, 25, 27, 28, 27, 28, 30, 27, 11, 10, 23, 31, 129, 
    41, 35, 30, 24, 9, 0, 0, 77, 60, 42, 31, 21, 30, 27, 26, 30, 34, 32, 30, 26, 29, 25, 23, 30, 34, 28, 11, 9, 26, 47, 33, 117, 
    35, 31, 30, 29, 24, 0, 0, 89, 60, 45, 42, 32, 32, 32, 31, 24, 21, 18, 22, 24, 27, 31, 30, 29, 23, 12, 2, 12, 22, 43, 21, 110, 
    44, 34, 26, 30, 28, 19, 0, 43, 53, 37, 31, 32, 38, 41, 43, 33, 27, 23, 17, 17, 22, 29, 31, 21, 8, 0, 1, 18, 40, 50, 24, 102, 
    40, 37, 25, 31, 30, 34, 29, 30, 45, 42, 32, 33, 30, 33, 42, 41, 36, 29, 23, 28, 34, 30, 31, 19, 6, 0, 17, 38, 49, 42, 39, 93, 
    82, 93, 82, 81, 81, 82, 82, 79, 83, 79, 72, 76, 75, 76, 70, 63, 66, 72, 77, 89, 95, 89, 86, 73, 73, 79, 97, 110, 102, 82, 85, 110, 
    
    -- channel=12
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 1, 0, 1, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 0, 0, 
    13, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 8, 0, 0, 0, 
    1, 0, 6, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 21, 0, 0, 0, 
    0, 0, 0, 20, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 27, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 24, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=13
    3, 105, 109, 113, 110, 105, 103, 108, 100, 98, 98, 106, 112, 108, 106, 103, 95, 92, 93, 95, 97, 94, 90, 91, 86, 86, 78, 75, 65, 58, 50, 0, 
    83, 204, 209, 214, 215, 208, 211, 213, 208, 203, 206, 217, 219, 211, 205, 201, 193, 192, 188, 188, 176, 171, 167, 167, 174, 178, 175, 169, 154, 143, 132, 17, 
    77, 190, 198, 206, 215, 213, 218, 218, 212, 211, 239, 253, 250, 223, 200, 199, 199, 184, 189, 179, 184, 174, 158, 149, 139, 155, 157, 163, 156, 149, 140, 22, 
    75, 188, 196, 202, 208, 213, 216, 217, 212, 221, 306, 324, 333, 252, 208, 196, 179, 164, 171, 193, 228, 226, 209, 170, 159, 143, 148, 153, 159, 156, 149, 24, 
    75, 191, 201, 201, 206, 211, 214, 212, 209, 215, 297, 348, 342, 238, 175, 160, 136, 134, 172, 241, 302, 307, 273, 235, 191, 156, 137, 131, 153, 166, 165, 31, 
    82, 166, 173, 162, 186, 208, 211, 208, 205, 210, 275, 315, 308, 230, 178, 149, 111, 130, 208, 303, 365, 358, 322, 283, 243, 201, 134, 111, 135, 160, 171, 36, 
    95, 178, 150, 134, 175, 206, 205, 206, 206, 203, 208, 230, 250, 234, 200, 168, 150, 172, 240, 332, 389, 371, 314, 276, 256, 199, 131, 89, 115, 149, 172, 43, 
    132, 220, 178, 157, 219, 223, 208, 215, 237, 217, 222, 229, 279, 304, 267, 220, 196, 198, 224, 310, 365, 358, 295, 251, 227, 190, 137, 84, 87, 125, 159, 49, 
    205, 328, 284, 272, 299, 252, 210, 267, 339, 380, 358, 347, 359, 379, 310, 249, 208, 188, 192, 262, 331, 368, 313, 250, 214, 185, 158, 104, 70, 92, 132, 41, 
    243, 436, 393, 415, 379, 286, 205, 314, 435, 545, 510, 471, 435, 421, 341, 249, 218, 160, 165, 239, 337, 423, 347, 276, 227, 202, 193, 134, 76, 66, 99, 20, 
    266, 496, 466, 506, 436, 321, 214, 292, 475, 611, 608, 541, 491, 449, 373, 280, 230, 150, 175, 277, 407, 488, 379, 298, 231, 228, 224, 185, 112, 79, 77, 2, 
    257, 510, 482, 534, 464, 334, 223, 248, 409, 517, 548, 515, 508, 495, 431, 322, 274, 181, 232, 335, 491, 516, 384, 288, 228, 232, 230, 212, 160, 127, 91, 0, 
    258, 515, 485, 525, 464, 316, 231, 192, 300, 382, 478, 474, 549, 558, 496, 375, 316, 229, 288, 396, 529, 503, 358, 262, 208, 215, 227, 233, 215, 191, 133, 11, 
    263, 526, 500, 527, 437, 291, 232, 180, 242, 300, 420, 466, 569, 576, 518, 418, 357, 273, 322, 415, 522, 485, 355, 273, 230, 218, 238, 263, 260, 232, 173, 26, 
    283, 554, 534, 538, 415, 300, 240, 206, 237, 278, 449, 556, 629, 601, 486, 412, 357, 282, 322, 414, 504, 454, 347, 260, 221, 218, 255, 289, 277, 247, 188, 44, 
    314, 589, 568, 572, 439, 354, 274, 264, 227, 289, 415, 559, 595, 504, 413, 363, 323, 265, 314, 379, 467, 440, 367, 278, 231, 228, 259, 277, 257, 223, 189, 58, 
    353, 631, 603, 609, 486, 393, 335, 329, 294, 298, 371, 497, 480, 396, 336, 290, 291, 275, 279, 296, 359, 349, 319, 243, 175, 182, 224, 241, 232, 210, 204, 67, 
    386, 665, 637, 643, 539, 427, 375, 380, 354, 312, 299, 354, 329, 328, 318, 283, 298, 288, 298, 301, 289, 284, 273, 184, 137, 133, 189, 213, 229, 227, 223, 73, 
    397, 671, 655, 653, 575, 444, 392, 380, 403, 364, 278, 289, 246, 317, 351, 349, 335, 314, 298, 298, 263, 242, 186, 109, 111, 126, 197, 220, 251, 245, 224, 71, 
    381, 641, 654, 646, 593, 473, 420, 423, 433, 397, 270, 246, 256, 359, 434, 464, 401, 319, 276, 264, 232, 170, 98, 70, 97, 153, 211, 234, 250, 234, 207, 64, 
    350, 593, 647, 630, 583, 472, 431, 477, 562, 541, 409, 342, 365, 463, 559, 579, 483, 374, 270, 226, 171, 133, 112, 121, 167, 220, 250, 263, 256, 237, 216, 76, 
    322, 571, 651, 626, 579, 485, 483, 571, 714, 697, 540, 449, 434, 502, 569, 560, 472, 368, 256, 189, 154, 156, 169, 199, 231, 266, 292, 309, 299, 288, 270, 128, 
    273, 539, 626, 630, 595, 526, 561, 687, 852, 778, 624, 472, 422, 444, 458, 445, 400, 346, 269, 223, 212, 231, 256, 282, 300, 314, 329, 342, 339, 331, 319, 173, 
    222, 461, 545, 588, 577, 575, 636, 775, 848, 746, 555, 397, 339, 334, 333, 324, 307, 291, 267, 263, 273, 285, 298, 310, 330, 343, 357, 364, 358, 351, 348, 190, 
    188, 396, 440, 513, 539, 604, 691, 805, 771, 598, 394, 309, 283, 278, 272, 266, 267, 270, 269, 273, 289, 303, 313, 330, 350, 369, 375, 374, 371, 381, 392, 226, 
    182, 359, 359, 407, 461, 577, 715, 786, 677, 459, 330, 309, 303, 298, 287, 280, 275, 275, 275, 283, 300, 321, 341, 357, 370, 377, 369, 377, 396, 424, 444, 270, 
    199, 369, 335, 343, 384, 552, 710, 743, 586, 379, 312, 321, 312, 303, 286, 279, 280, 284, 291, 306, 317, 337, 356, 373, 379, 368, 364, 386, 420, 449, 460, 262, 
    201, 376, 338, 323, 345, 477, 643, 624, 514, 337, 318, 329, 326, 319, 298, 288, 284, 293, 306, 322, 335, 348, 359, 364, 361, 354, 367, 394, 433, 420, 405, 202, 
    206, 387, 350, 331, 335, 392, 495, 481, 408, 299, 292, 308, 325, 331, 318, 310, 306, 316, 329, 339, 341, 339, 337, 339, 351, 372, 410, 450, 449, 376, 331, 151, 
    212, 388, 354, 338, 337, 339, 374, 358, 315, 263, 260, 273, 294, 306, 307, 308, 313, 334, 358, 369, 362, 347, 328, 330, 360, 424, 483, 495, 436, 345, 281, 139, 
    218, 386, 352, 334, 335, 316, 305, 285, 258, 234, 228, 237, 259, 261, 263, 269, 289, 328, 367, 385, 379, 352, 319, 332, 378, 464, 518, 503, 426, 338, 275, 138, 
    103, 205, 182, 171, 173, 167, 150, 135, 119, 106, 100, 101, 106, 106, 109, 114, 130, 161, 196, 216, 207, 182, 162, 172, 208, 267, 299, 283, 223, 172, 136, 55, 
    
    -- channel=14
    0, 18, 17, 16, 21, 26, 23, 25, 25, 25, 21, 18, 21, 24, 27, 27, 29, 30, 27, 21, 16, 14, 11, 14, 15, 19, 18, 18, 18, 19, 21, 0, 
    107, 174, 174, 166, 167, 173, 175, 175, 175, 182, 174, 165, 166, 176, 188, 192, 190, 184, 168, 152, 137, 129, 129, 133, 135, 140, 143, 149, 152, 151, 144, 64, 
    110, 178, 180, 173, 175, 176, 181, 179, 179, 177, 179, 176, 172, 179, 188, 184, 175, 155, 143, 144, 134, 126, 113, 110, 112, 115, 128, 146, 152, 151, 147, 68, 
    111, 179, 181, 170, 170, 176, 179, 178, 180, 179, 190, 164, 160, 172, 167, 150, 127, 115, 132, 110, 93, 81, 89, 97, 99, 120, 119, 130, 142, 146, 142, 65, 
    101, 156, 160, 167, 172, 183, 182, 183, 183, 182, 169, 106, 132, 139, 122, 109, 119, 125, 94, 67, 60, 52, 43, 47, 67, 63, 90, 114, 131, 141, 148, 67, 
    84, 124, 127, 150, 171, 183, 187, 186, 187, 189, 202, 198, 164, 141, 138, 133, 91, 71, 70, 75, 69, 56, 51, 60, 42, 51, 77, 96, 110, 121, 134, 61, 
    79, 103, 143, 154, 158, 175, 185, 183, 181, 180, 170, 170, 152, 109, 81, 69, 51, 56, 73, 72, 73, 79, 77, 59, 49, 50, 41, 69, 99, 113, 131, 63, 
    57, 67, 89, 129, 150, 175, 190, 187, 182, 166, 158, 155, 126, 86, 63, 51, 46, 51, 70, 78, 74, 81, 78, 66, 67, 55, 51, 42, 76, 108, 126, 61, 
    33, 70, 75, 73, 130, 169, 180, 192, 197, 168, 163, 125, 93, 81, 71, 70, 61, 46, 59, 113, 101, 81, 80, 84, 72, 52, 44, 44, 63, 92, 108, 54, 
    35, 55, 69, 82, 113, 161, 165, 175, 128, 81, 56, 96, 91, 90, 73, 60, 54, 51, 66, 97, 99, 98, 67, 56, 64, 58, 44, 30, 41, 85, 104, 38, 
    45, 90, 56, 99, 127, 165, 159, 161, 111, 105, 88, 108, 96, 89, 76, 52, 68, 37, 72, 92, 74, 89, 59, 63, 60, 52, 60, 49, 35, 53, 89, 36, 
    31, 89, 85, 98, 114, 152, 148, 150, 186, 125, 93, 104, 111, 87, 94, 79, 64, 47, 83, 77, 69, 96, 76, 74, 65, 62, 48, 48, 33, 37, 59, 36, 
    30, 98, 94, 83, 109, 145, 152, 124, 147, 110, 122, 148, 131, 100, 97, 89, 64, 31, 83, 87, 103, 98, 81, 62, 53, 62, 65, 62, 44, 43, 56, 31, 
    35, 94, 74, 77, 129, 141, 151, 126, 130, 110, 124, 116, 122, 88, 88, 90, 80, 48, 80, 92, 94, 95, 85, 70, 64, 74, 76, 61, 53, 55, 69, 29, 
    37, 94, 79, 74, 94, 128, 142, 130, 143, 130, 136, 127, 134, 134, 109, 71, 65, 73, 92, 91, 98, 92, 50, 36, 46, 45, 57, 63, 58, 80, 107, 37, 
    45, 89, 88, 82, 61, 106, 114, 121, 108, 102, 114, 67, 56, 104, 88, 92, 88, 66, 93, 113, 106, 91, 98, 81, 67, 56, 54, 65, 79, 109, 117, 50, 
    52, 90, 88, 77, 45, 77, 85, 107, 107, 140, 99, 128, 127, 89, 100, 87, 84, 90, 97, 72, 100, 88, 51, 34, 41, 50, 63, 88, 113, 119, 126, 62, 
    52, 89, 88, 87, 60, 68, 86, 72, 93, 107, 99, 122, 123, 111, 113, 80, 82, 84, 91, 153, 168, 86, 59, 70, 59, 67, 83, 95, 116, 127, 146, 69, 
    67, 93, 90, 95, 72, 50, 77, 68, 70, 83, 97, 104, 59, 81, 89, 64, 74, 83, 75, 81, 66, 81, 83, 48, 57, 59, 91, 106, 123, 146, 157, 69, 
    82, 106, 100, 99, 84, 55, 78, 94, 89, 50, 25, 79, 70, 112, 100, 62, 68, 91, 69, 54, 38, 51, 46, 29, 26, 33, 80, 118, 142, 154, 153, 69, 
    98, 104, 105, 106, 85, 50, 64, 84, 87, 135, 112, 98, 116, 99, 87, 85, 61, 73, 94, 91, 88, 59, 43, 47, 33, 61, 73, 96, 111, 117, 108, 44, 
    98, 89, 106, 105, 89, 81, 114, 102, 53, 43, 60, 24, 15, 20, 45, 44, 23, 17, 22, 54, 47, 24, 0, 0, 0, 19, 47, 81, 80, 77, 77, 25, 
    58, 54, 83, 95, 90, 86, 110, 103, 124, 58, 4, 40, 48, 55, 70, 62, 54, 53, 29, 2, 0, 0, 0, 0, 0, 0, 7, 9, 8, 10, 2, 0, 
    39, 50, 55, 72, 63, 67, 102, 120, 123, 95, 105, 72, 62, 62, 59, 55, 35, 14, 5, 1, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 
    16, 43, 65, 58, 65, 125, 128, 125, 96, 93, 52, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 18, 47, 55, 105, 117, 107, 97, 76, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 21, 46, 71, 98, 94, 91, 35, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 61, 71, 61, 57, 13, 2, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 34, 76, 33, 48, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 0, 0, 0, 0, 0, 56, 56, 23, 14, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 5, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    44, 68, 69, 67, 68, 72, 70, 70, 70, 70, 72, 70, 69, 73, 77, 78, 79, 77, 72, 66, 61, 60, 60, 63, 64, 67, 68, 69, 71, 70, 67, 50, 
    109, 84, 91, 88, 86, 88, 89, 87, 86, 89, 88, 83, 84, 92, 98, 99, 97, 91, 80, 70, 63, 61, 64, 68, 71, 72, 76, 82, 85, 82, 77, 50, 
    110, 87, 97, 96, 93, 90, 90, 86, 90, 85, 84, 76, 74, 87, 95, 94, 89, 76, 62, 55, 38, 34, 38, 47, 60, 60, 68, 74, 81, 79, 76, 52, 
    111, 87, 95, 96, 94, 95, 91, 89, 90, 89, 79, 53, 46, 73, 81, 77, 72, 58, 55, 25, 10, 0, 6, 23, 27, 47, 51, 61, 71, 75, 74, 51, 
    107, 77, 77, 86, 87, 95, 93, 92, 92, 92, 89, 51, 37, 52, 65, 57, 52, 50, 21, 8, 0, 0, 0, 0, 14, 11, 41, 55, 63, 66, 72, 50, 
    95, 58, 58, 73, 80, 88, 97, 93, 94, 91, 79, 86, 22, 26, 37, 39, 19, 15, 18, 2, 0, 0, 0, 0, 0, 0, 16, 41, 58, 64, 69, 51, 
    80, 18, 39, 62, 68, 84, 98, 97, 91, 87, 73, 69, 40, 18, 8, 10, 11, 3, 14, 0, 0, 0, 0, 0, 0, 0, 0, 28, 57, 64, 63, 49, 
    52, 0, 0, 52, 63, 77, 92, 92, 83, 70, 60, 48, 23, 3, 0, 0, 4, 0, 6, 14, 0, 0, 0, 0, 4, 0, 1, 9, 49, 69, 60, 41, 
    30, 0, 0, 8, 43, 67, 84, 78, 60, 16, 18, 11, 6, 0, 0, 0, 1, 0, 0, 29, 8, 0, 0, 2, 2, 0, 0, 8, 31, 66, 62, 35, 
    38, 0, 0, 0, 3, 51, 79, 74, 26, 0, 0, 3, 0, 0, 0, 0, 0, 2, 10, 15, 10, 0, 0, 0, 2, 1, 0, 0, 11, 54, 70, 30, 
    29, 0, 0, 0, 0, 35, 70, 72, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 63, 41, 
    27, 0, 0, 0, 0, 28, 73, 48, 75, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 0, 0, 0, 0, 0, 2, 0, 0, 0, 5, 33, 45, 
    28, 0, 0, 0, 0, 25, 72, 53, 54, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 21, 32, 
    31, 0, 0, 0, 0, 19, 61, 58, 40, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 23, 
    32, 0, 0, 0, 0, 12, 46, 42, 31, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 40, 25, 
    34, 0, 0, 0, 0, 0, 23, 18, 11, 33, 13, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 8, 30, 50, 43, 
    31, 0, 0, 0, 0, 0, 7, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 1, 17, 14, 0, 0, 0, 1, 12, 5, 5, 26, 38, 59, 44, 
    29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 2, 0, 0, 0, 0, 0, 0, 0, 26, 17, 0, 0, 0, 1, 17, 27, 32, 48, 63, 75, 42, 
    38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 0, 3, 0, 0, 0, 0, 6, 0, 0, 18, 10, 0, 15, 13, 30, 53, 55, 71, 72, 43, 
    47, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 17, 0, 0, 0, 0, 0, 12, 0, 0, 0, 1, 9, 7, 13, 25, 54, 54, 57, 56, 34, 
    53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 2, 0, 0, 
    44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end inmem_package;
