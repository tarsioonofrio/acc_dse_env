library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    31766, -20771, 6499, 19371, -20879, -5812, 8847, 13261, 3788, -3044, -15547, 16289, 9585, -36823, -800, 12902,

    -- weights
    -- filter=0 channel=0
    22, 22, -39, 0, 60, -49, -8, 27, 20,
    -- filter=0 channel=1
    43, 31, -78, 8, 25, -38, -43, 47, -23,
    -- filter=0 channel=2
    44, -40, -88, -31, -8, -85, 5, -12, 14,
    -- filter=1 channel=0
    36, -14, 14, -55, -17, 38, 36, 14, 30,
    -- filter=1 channel=1
    46, 38, 17, 75, 75, 55, 84, 20, 22,
    -- filter=1 channel=2
    27, -24, -16, -35, -14, -32, 47, 27, 22,
    -- filter=2 channel=0
    37, 19, 6, 35, -11, 35, 5, -12, 2,
    -- filter=2 channel=1
    -73, -35, 56, -27, -32, 52, -47, -55, 25,
    -- filter=2 channel=2
    -46, -18, 39, -49, -34, 3, -67, 46, 58,
    -- filter=3 channel=0
    35, 52, 38, -84, 9, -47, -43, -41, -21,
    -- filter=3 channel=1
    52, 123, 69, 4, 70, 33, 54, -11, 55,
    -- filter=3 channel=2
    45, -35, -38, -75, -78, -18, -29, -95, -49,
    -- filter=4 channel=0
    49, -29, 44, 32, 15, -18, 6, -7, 67,
    -- filter=4 channel=1
    -2, -23, -76, -21, -41, -50, 19, -48, -79,
    -- filter=4 channel=2
    85, 72, 0, 80, 78, 29, 97, 86, 29,
    -- filter=5 channel=0
    -59, 8, 17, 46, -28, 32, -36, -3, -17,
    -- filter=5 channel=1
    73, 74, 71, 47, 79, 19, -1, 78, 95,
    -- filter=5 channel=2
    -55, -44, 47, 54, -47, 6, -43, -26, -39,
    -- filter=6 channel=0
    41, 0, -20, -19, 19, -46, -20, 58, 18,
    -- filter=6 channel=1
    8, 12, -9, 11, 61, -35, 41, 4, -35,
    -- filter=6 channel=2
    -27, -55, -11, 32, -16, -12, -45, 43, -37,
    -- filter=7 channel=0
    -35, 34, -4, -68, -18, -25, -66, -21, 44,
    -- filter=7 channel=1
    -60, -21, 31, -45, 55, -17, -47, 33, 30,
    -- filter=7 channel=2
    21, 44, 17, -46, 57, 48, -24, 34, -1,
    -- filter=8 channel=0
    3, 19, -31, -3, -17, -31, 30, -10, -9,
    -- filter=8 channel=1
    -3, 31, -22, -36, 34, -24, -33, -36, 31,
    -- filter=8 channel=2
    -6, 0, -32, 21, -32, 3, -17, 33, -45,
    -- filter=9 channel=0
    -58, -60, -79, -103, -97, -92, -87, -32, -93,
    -- filter=9 channel=1
    18, 23, -54, -5, 30, 5, 20, -14, 10,
    -- filter=9 channel=2
    44, 98, 119, 120, 95, 109, 100, 50, 124,
    -- filter=10 channel=0
    -36, -6, 56, -12, -6, -20, -52, 20, 55,
    -- filter=10 channel=1
    -12, 7, 22, -7, 63, 65, 2, 61, 57,
    -- filter=10 channel=2
    8, 46, 52, -10, 6, 30, 45, -10, 68,
    -- filter=11 channel=0
    26, -29, -41, 29, 48, 12, -14, -36, -17,
    -- filter=11 channel=1
    -2, -1, 29, 20, 28, -57, -7, -29, -32,
    -- filter=11 channel=2
    7, 30, -54, -28, 54, -1, -11, 16, -37,
    -- filter=12 channel=0
    -30, -6, 15, -30, -14, 37, -24, -40, 27,
    -- filter=12 channel=1
    -1, 29, -8, -13, -22, 30, 30, -26, 3,
    -- filter=12 channel=2
    -31, -37, -15, 42, -34, -45, -25, 14, -33,
    -- filter=13 channel=0
    -7, 3, 39, -4, -12, 11, 39, 24, 50,
    -- filter=13 channel=1
    37, 35, 27, 43, 31, 34, 70, 11, 60,
    -- filter=13 channel=2
    66, 90, 68, 86, 104, 38, 63, 43, 64,
    -- filter=14 channel=0
    5, 43, 34, -4, -96, -8, 18, -4, 25,
    -- filter=14 channel=1
    80, 114, 80, 46, -13, 25, 51, 70, 87,
    -- filter=14 channel=2
    -65, -14, -43, -31, -101, -50, -53, -11, -28,
    -- filter=15 channel=0
    -31, 65, 53, 58, -7, 27, 52, 37, 48,
    -- filter=15 channel=1
    -54, 39, -29, -21, -52, -29, -55, -18, -36,
    -- filter=15 channel=2
    -36, -17, -52, -31, -21, 32, -39, -44, -17,

    others => 0);
end iwght_package;
