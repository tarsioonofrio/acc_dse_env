library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    -- layer=1
    13182, 857, -1403, -1481, -1386, -1702, 4814, -1112, 3134, -893, -2244, -724, -558, -1042, -665, 4886, -1365, 8574, 9081, -1237, -1695, -4022, 757, 3610, -5065, -546, -1208, -2026, -1548, -5710, -1071, 8699, -2752, -4685, -7459, 1773, 3211, -8344, -867, 9416, -3190, -1046, 2971, 6404, -3892, -503, 2180, -678, -410, -4684, -3199, -3910, -725, -3588, 2659, -334, 5800, 2773, -146, -693, 7196, 2632, 3027, -1515, 12255, -11980, -2840, -2502, 4627, -9782, -360, -726, 18523, -500, -1343, -7138, -203, -869, 4635, -569, -1520, -541, -864, -1825, 2788, -1557, 9287, -403, -2095, -2302, -1554, 4356, -661, -783, -2877, -473, -6341, 9769, 483, -1998, -339, -2337, 9329, -1420, -753, -1441, -1228, -417, -2382, -2463, 9076, -1695, 4187, 13102, 4611, 3616, -1121, -2645, -673, -1274, 2520, 10064, 1994, 15266, -1207, -2008, -437, -3671, -203, 8744, -547, -482, 2470, -1091, -3380, -367, 2901, -4067, -6458, -4651, -1863, 8362, -681, 10452, -6145, -599, -1251, -2348, -2519, -3098, -470, -496, -637, -457, 1125, -902, -5344, -1561, -602, -941, -487, -8230, 4670, -430, -763, 7877, 327, -5405, -3225, -565, -4628, -560, -3130, 4619, -620, -778, 1638, -503, -4925, -2685, -697, -2200, -1647, 11771, -1297, -437, -666, 5216, -769, -1611, 3895, -769, 301, -1081, -1927, 222, -542, 909, -2699, 6271, -1585, -494, -2279, -686, 11000, -679, -1461, -2017, -575, -2877, -1590, -681, -676, -1104, -1120, -4385, -1406, -781, 2038, -695, -751, -1413, -2590, -1495, -542, -882, 16086, -618, -706, -1347, -2728, -104, -979, -695, -538, -526, -3338, -53, -1191, -1360, -2752, -746, 7852, -4932, -606, -922, -558, -493, -1283, -1136, -1324, -438, 964, -4596, -2359, -1293,

    -- weights
    -- layer=1 filter=0 channel=0
    3, -2, -4, -1, -11, 3, -14, 2, 4,
    -- layer=1 filter=0 channel=1
    5, 6, -17, 28, 4, -4, -15, -5, 1,
    -- layer=1 filter=0 channel=2
    -27, 16, 16, 3, -1, -1, -15, 9, 14,
    -- layer=1 filter=0 channel=3
    0, -4, 1, 1, -3, 2, 0, 7, 10,
    -- layer=1 filter=0 channel=4
    0, 5, 7, -6, -14, -2, -3, -7, -8,
    -- layer=1 filter=0 channel=5
    8, 10, -2, 9, 5, 8, 18, -4, 11,
    -- layer=1 filter=0 channel=6
    -28, -15, -1, -59, -58, -30, 1, -10, -29,
    -- layer=1 filter=0 channel=7
    -18, -14, -19, -14, -74, -51, -12, -32, -15,
    -- layer=1 filter=0 channel=8
    13, -12, -20, 17, 14, -2, 12, 1, 21,
    -- layer=1 filter=0 channel=9
    -38, -55, -33, -26, -44, -52, -27, -21, -18,
    -- layer=1 filter=0 channel=10
    16, -7, -12, -10, -43, -43, 4, -6, 0,
    -- layer=1 filter=0 channel=11
    -16, -10, -7, 1, -14, -5, -6, -22, -15,
    -- layer=1 filter=0 channel=12
    -80, -65, -54, -45, -60, -23, 2, -5, -24,
    -- layer=1 filter=0 channel=13
    3, -4, -14, -33, -30, -18, -8, -1, -4,
    -- layer=1 filter=0 channel=14
    -12, -3, -27, -19, 6, -6, -14, 42, -27,
    -- layer=1 filter=0 channel=15
    -19, -26, -6, -40, -50, -48, -43, -41, -57,
    -- layer=1 filter=0 channel=16
    21, -10, -19, 4, 21, 1, 24, 5, 16,
    -- layer=1 filter=0 channel=17
    -4, 0, -14, -19, -34, -21, -17, -9, -8,
    -- layer=1 filter=0 channel=18
    7, -7, -18, 9, 16, 13, -15, -17, -20,
    -- layer=1 filter=0 channel=19
    19, -6, 7, -3, 0, 0, 24, -4, -1,
    -- layer=1 filter=0 channel=20
    14, -3, 0, -19, -23, -24, -12, 8, 9,
    -- layer=1 filter=0 channel=21
    -12, 7, -9, -3, 3, -10, -12, 6, -7,
    -- layer=1 filter=0 channel=22
    -18, 8, -15, -12, -37, -43, -19, -12, 1,
    -- layer=1 filter=0 channel=23
    -13, -45, -17, 16, -36, -33, 1, -30, -30,
    -- layer=1 filter=0 channel=24
    20, -10, 7, 5, 7, 20, 16, 23, 39,
    -- layer=1 filter=0 channel=25
    8, -13, -21, 1, -38, -16, 10, 3, 4,
    -- layer=1 filter=0 channel=26
    20, -29, -6, -13, -37, -14, 3, -5, 1,
    -- layer=1 filter=0 channel=27
    -46, -39, -50, -6, -29, -28, -6, -3, -4,
    -- layer=1 filter=0 channel=28
    -22, 12, -28, -6, -18, -48, 5, 3, -15,
    -- layer=1 filter=0 channel=29
    -22, -17, -25, -28, -28, -10, -18, -28, -17,
    -- layer=1 filter=0 channel=30
    56, 16, -6, 11, 9, 31, 24, -3, -25,
    -- layer=1 filter=0 channel=31
    -21, -14, -38, 6, 7, 3, -12, -15, -18,
    -- layer=1 filter=0 channel=32
    38, -23, 0, 0, -29, 7, 8, -40, 3,
    -- layer=1 filter=0 channel=33
    0, 3, -11, -8, -2, -3, 14, 7, 3,
    -- layer=1 filter=0 channel=34
    -31, 6, -2, 0, -14, -9, 2, 0, -3,
    -- layer=1 filter=0 channel=35
    -12, -12, -10, -5, -8, -19, -8, -4, -16,
    -- layer=1 filter=0 channel=36
    8, 7, 11, 11, 1, 8, 3, 0, 0,
    -- layer=1 filter=0 channel=37
    34, 8, 6, 3, 17, 19, 9, 3, 13,
    -- layer=1 filter=0 channel=38
    9, 5, -9, -19, -8, -9, -4, -8, -5,
    -- layer=1 filter=0 channel=39
    -19, -18, -17, -9, -16, -12, 11, -2, -3,
    -- layer=1 filter=0 channel=40
    -14, -43, -49, -27, -49, -40, 11, 7, -28,
    -- layer=1 filter=0 channel=41
    37, -7, -5, 5, -14, -3, 19, -35, 45,
    -- layer=1 filter=0 channel=42
    -29, -25, 18, -27, -4, 2, -31, -14, -11,
    -- layer=1 filter=0 channel=43
    -4, -13, -33, 17, 2, -11, 20, 0, 14,
    -- layer=1 filter=0 channel=44
    3, -61, 2, -19, -54, -12, -9, -44, -3,
    -- layer=1 filter=0 channel=45
    -26, -18, -6, -7, -30, -4, -28, -28, -23,
    -- layer=1 filter=0 channel=46
    0, -12, -12, -42, -23, -16, 3, -36, -47,
    -- layer=1 filter=0 channel=47
    13, -47, -24, -18, -38, -53, -21, -32, -10,
    -- layer=1 filter=0 channel=48
    12, 3, 9, -2, 20, -4, 7, 5, -5,
    -- layer=1 filter=0 channel=49
    -7, -10, -3, -35, -22, -20, -23, -25, -15,
    -- layer=1 filter=0 channel=50
    -7, -13, -13, -14, -18, -29, -15, -30, -20,
    -- layer=1 filter=0 channel=51
    5, 22, -2, 3, 14, -16, 8, 8, -6,
    -- layer=1 filter=0 channel=52
    0, 6, 5, 19, 1, 9, -14, -21, -2,
    -- layer=1 filter=0 channel=53
    0, 1, -2, -20, -13, -3, -14, -17, -6,
    -- layer=1 filter=0 channel=54
    -5, -1, -19, -13, -19, -5, 8, 0, 16,
    -- layer=1 filter=0 channel=55
    10, -6, -2, 29, 15, 4, 16, 6, 23,
    -- layer=1 filter=0 channel=56
    -4, 4, -5, -4, 9, 2, -11, -10, 7,
    -- layer=1 filter=0 channel=57
    -12, -43, -27, -26, -70, -48, -27, -39, -18,
    -- layer=1 filter=0 channel=58
    -17, -85, -33, -4, -81, -16, 6, -28, -12,
    -- layer=1 filter=0 channel=59
    -3, 2, -1, -4, -1, -11, -3, -14, -6,
    -- layer=1 filter=0 channel=60
    6, 9, 4, 2, 5, -2, 3, 12, 5,
    -- layer=1 filter=0 channel=61
    6, 8, -8, 2, -1, -6, 10, 5, 8,
    -- layer=1 filter=0 channel=62
    1, -24, -10, 16, 15, 0, 18, 0, 14,
    -- layer=1 filter=0 channel=63
    10, -11, 2, 6, 8, 25, -9, -9, 10,
    -- layer=1 filter=0 channel=64
    8, 5, 10, 8, 7, 0, -2, 7, 13,
    -- layer=1 filter=0 channel=65
    -5, 15, -9, 1, 6, -2, -14, -3, -10,
    -- layer=1 filter=0 channel=66
    2, 6, 5, 0, 9, 9, -12, 8, 4,
    -- layer=1 filter=0 channel=67
    -12, -25, -29, -21, -31, -41, -60, -58, -54,
    -- layer=1 filter=0 channel=68
    -7, -54, -4, -26, -48, -19, -2, -55, -23,
    -- layer=1 filter=0 channel=69
    -2, -24, -8, -3, -2, -9, 10, 1, -13,
    -- layer=1 filter=0 channel=70
    20, 0, -28, 28, 14, -3, -65, -38, -53,
    -- layer=1 filter=0 channel=71
    -11, 6, 6, 15, 21, 21, 27, 36, 24,
    -- layer=1 filter=0 channel=72
    23, -21, -29, 2, -8, -26, 4, -28, -26,
    -- layer=1 filter=0 channel=73
    1, -2, 6, -1, 3, -6, -3, -9, 3,
    -- layer=1 filter=0 channel=74
    7, -1, -32, -18, -16, -7, 16, -13, -47,
    -- layer=1 filter=0 channel=75
    -7, -19, -31, -6, -25, -4, 14, 14, -30,
    -- layer=1 filter=0 channel=76
    14, 6, 7, 3, -3, -4, 6, -18, -4,
    -- layer=1 filter=0 channel=77
    2, 11, -8, 8, 8, -5, -6, 3, 5,
    -- layer=1 filter=0 channel=78
    3, -4, 3, -11, -5, -3, 6, -9, -7,
    -- layer=1 filter=0 channel=79
    10, -16, -8, 12, 20, 10, 2, 0, 8,
    -- layer=1 filter=0 channel=80
    -1, -1, -5, 0, -6, -9, -8, -5, -1,
    -- layer=1 filter=0 channel=81
    -5, 2, 3, 19, 29, 16, 13, 17, 33,
    -- layer=1 filter=0 channel=82
    -14, -4, -13, 10, 19, -2, 8, 9, 5,
    -- layer=1 filter=0 channel=83
    -8, 1, 0, 3, -5, -14, -13, -25, -12,
    -- layer=1 filter=0 channel=84
    23, -11, -8, 6, 19, 18, 21, -22, 30,
    -- layer=1 filter=0 channel=85
    -23, -48, 2, -27, -48, -31, -16, -39, -5,
    -- layer=1 filter=0 channel=86
    0, 5, -5, 5, 2, -4, -5, -2, -17,
    -- layer=1 filter=0 channel=87
    20, -21, 31, -27, -20, -45, -9, -27, -7,
    -- layer=1 filter=0 channel=88
    -14, -8, -16, -9, -18, -2, -17, -24, -21,
    -- layer=1 filter=0 channel=89
    -12, 0, 2, -11, 2, 7, -3, 9, -3,
    -- layer=1 filter=0 channel=90
    -12, -80, -23, -14, -61, -18, -29, -43, -29,
    -- layer=1 filter=0 channel=91
    23, 9, 0, -17, -20, -14, -19, -14, -16,
    -- layer=1 filter=0 channel=92
    23, -8, -13, -3, -12, -47, 25, -6, 4,
    -- layer=1 filter=0 channel=93
    20, 25, 22, 25, 30, 18, 13, 17, 17,
    -- layer=1 filter=0 channel=94
    -1, -9, 6, -13, -8, -10, -6, -23, -16,
    -- layer=1 filter=0 channel=95
    37, 0, -2, 0, 21, 40, 17, 0, 16,
    -- layer=1 filter=0 channel=96
    3, 9, 7, 2, 0, -11, 9, 6, 11,
    -- layer=1 filter=0 channel=97
    6, 10, 5, 18, 6, 15, 10, 14, 18,
    -- layer=1 filter=0 channel=98
    19, 6, -16, 39, 11, -18, -9, -9, 4,
    -- layer=1 filter=0 channel=99
    -32, 12, 3, -49, -16, -81, 1, -3, -65,
    -- layer=1 filter=0 channel=100
    -9, -21, -32, 6, -12, -19, -11, -31, -18,
    -- layer=1 filter=0 channel=101
    16, 7, 9, -14, 1, -1, -10, 2, -12,
    -- layer=1 filter=0 channel=102
    -5, 12, 0, -3, -14, -11, -10, -22, -18,
    -- layer=1 filter=0 channel=103
    -12, -19, -17, 1, -9, -3, -25, -27, -2,
    -- layer=1 filter=0 channel=104
    -7, -1, 7, -17, -22, -20, -10, -16, -8,
    -- layer=1 filter=0 channel=105
    -1, 14, 14, 16, 14, 0, 13, 4, 5,
    -- layer=1 filter=0 channel=106
    -2, -2, 0, -38, -27, -14, -29, -14, 3,
    -- layer=1 filter=0 channel=107
    2, 19, 10, 13, 1, 17, 6, 5, 10,
    -- layer=1 filter=0 channel=108
    1, -86, -19, -18, -53, -25, -5, -31, 0,
    -- layer=1 filter=0 channel=109
    -2, 1, 7, 10, 1, -6, -5, 8, 2,
    -- layer=1 filter=0 channel=110
    2, 3, 6, -10, 10, 0, 0, -6, -1,
    -- layer=1 filter=0 channel=111
    41, -3, 5, 11, 34, 30, 16, -10, -3,
    -- layer=1 filter=0 channel=112
    22, -9, -13, 14, 18, 20, -29, -49, 18,
    -- layer=1 filter=0 channel=113
    -75, -61, -45, -34, -40, -37, -56, -53, -9,
    -- layer=1 filter=0 channel=114
    -3, -37, -42, 0, 10, 0, 38, 26, 10,
    -- layer=1 filter=0 channel=115
    15, 8, -2, -2, 1, -10, 8, -19, 13,
    -- layer=1 filter=0 channel=116
    -4, 5, -8, -8, -7, -2, -7, 5, 0,
    -- layer=1 filter=0 channel=117
    34, -34, -10, 6, -5, -1, -9, -42, 8,
    -- layer=1 filter=0 channel=118
    41, 6, -8, 12, 11, 23, 38, 2, -9,
    -- layer=1 filter=0 channel=119
    14, -49, 14, -19, -46, 2, -10, -36, 1,
    -- layer=1 filter=0 channel=120
    1, 11, -18, 6, -11, -22, -1, 9, 4,
    -- layer=1 filter=0 channel=121
    17, 4, -14, 21, -4, 16, 38, 13, -25,
    -- layer=1 filter=0 channel=122
    -8, 6, -5, -10, -9, 6, -2, 0, -9,
    -- layer=1 filter=0 channel=123
    10, -6, -22, 25, 0, 22, 24, 16, 5,
    -- layer=1 filter=0 channel=124
    -18, -2, 0, -18, -4, -21, -12, -20, -5,
    -- layer=1 filter=0 channel=125
    5, 1, -1, -43, -19, -13, -66, -70, -41,
    -- layer=1 filter=0 channel=126
    7, -5, 0, 37, -11, -44, -20, -23, 9,
    -- layer=1 filter=0 channel=127
    39, 6, -5, 6, 42, 28, 25, 5, -6,
    -- layer=1 filter=1 channel=0
    -1, 2, 8, 12, 0, 5, 5, 2, -6,
    -- layer=1 filter=1 channel=1
    -15, -12, -12, 22, 6, 20, 11, -20, 5,
    -- layer=1 filter=1 channel=2
    5, 11, 37, 37, 31, 13, 46, 66, 59,
    -- layer=1 filter=1 channel=3
    -6, 1, 9, -7, -1, 7, 0, -5, -10,
    -- layer=1 filter=1 channel=4
    6, -8, -5, -4, 2, -8, 7, 3, -6,
    -- layer=1 filter=1 channel=5
    -8, 20, 8, -20, -4, 11, -9, -31, -8,
    -- layer=1 filter=1 channel=6
    -62, -53, -67, -1, -5, -16, 37, 41, 38,
    -- layer=1 filter=1 channel=7
    -30, -51, -8, -50, -83, -54, -34, -54, -37,
    -- layer=1 filter=1 channel=8
    -2, 22, 5, 33, 24, 20, 8, -16, 18,
    -- layer=1 filter=1 channel=9
    24, 16, 45, -13, 0, 18, 38, 28, 31,
    -- layer=1 filter=1 channel=10
    -21, -64, 20, -57, -91, -48, -20, -41, -15,
    -- layer=1 filter=1 channel=11
    14, -8, -5, 2, 17, 12, -7, -11, -3,
    -- layer=1 filter=1 channel=12
    58, 33, 27, 18, 26, 43, 16, 32, 80,
    -- layer=1 filter=1 channel=13
    -39, -42, -49, 0, 15, 6, 32, 32, 14,
    -- layer=1 filter=1 channel=14
    24, 7, 58, -29, -22, -12, -41, -23, 19,
    -- layer=1 filter=1 channel=15
    -49, -14, -23, -18, 20, 31, -8, -17, -12,
    -- layer=1 filter=1 channel=16
    0, 8, 0, 11, 19, 21, -6, -4, 17,
    -- layer=1 filter=1 channel=17
    0, -1, -6, 12, 0, -6, 7, 15, 6,
    -- layer=1 filter=1 channel=18
    -1, 2, 21, 5, -12, 3, -9, -6, 13,
    -- layer=1 filter=1 channel=19
    48, 47, 24, -31, 16, -9, -18, -42, -23,
    -- layer=1 filter=1 channel=20
    -26, -10, -29, 2, 1, 14, 49, 42, 26,
    -- layer=1 filter=1 channel=21
    -33, -28, -31, -5, -11, 3, 4, -13, -8,
    -- layer=1 filter=1 channel=22
    -27, -38, -32, 37, 20, 2, 31, 35, 26,
    -- layer=1 filter=1 channel=23
    -29, -13, -21, -57, -36, -46, -36, -59, -35,
    -- layer=1 filter=1 channel=24
    9, 1, -3, -15, -1, -15, -31, -39, 12,
    -- layer=1 filter=1 channel=25
    -36, -38, -25, -7, -39, -43, -14, -63, -23,
    -- layer=1 filter=1 channel=26
    -13, -18, -22, 0, 37, 13, 37, 6, 34,
    -- layer=1 filter=1 channel=27
    -27, -6, -6, -21, -19, -8, -37, -25, -31,
    -- layer=1 filter=1 channel=28
    -15, -39, 6, -8, -39, -26, -27, -35, -8,
    -- layer=1 filter=1 channel=29
    -39, -21, -28, -37, -20, -12, -25, -22, -27,
    -- layer=1 filter=1 channel=30
    38, 12, 27, -29, -19, -18, -28, -7, -5,
    -- layer=1 filter=1 channel=31
    -9, 0, -21, -2, -11, 17, 1, 29, 39,
    -- layer=1 filter=1 channel=32
    -43, -59, -46, -62, -41, -33, -1, -44, -5,
    -- layer=1 filter=1 channel=33
    -27, -1, -14, -19, -8, -6, 1, -3, -4,
    -- layer=1 filter=1 channel=34
    -25, -29, -23, 13, 4, 24, 0, 15, -23,
    -- layer=1 filter=1 channel=35
    -2, -2, 5, 0, -9, 5, 3, -3, -2,
    -- layer=1 filter=1 channel=36
    24, 12, 26, 9, 19, 18, -11, -4, -17,
    -- layer=1 filter=1 channel=37
    10, 18, 6, -21, -10, -4, -34, -42, -1,
    -- layer=1 filter=1 channel=38
    -34, -43, -23, -2, 2, 0, 33, 34, 28,
    -- layer=1 filter=1 channel=39
    13, 10, 9, 3, 5, -2, -4, -11, -10,
    -- layer=1 filter=1 channel=40
    -52, -55, -36, 15, 1, 3, 44, 67, 43,
    -- layer=1 filter=1 channel=41
    12, -20, 26, -58, -53, -19, 0, -18, 6,
    -- layer=1 filter=1 channel=42
    23, 14, 32, 36, 56, 35, 58, 66, 58,
    -- layer=1 filter=1 channel=43
    -14, -5, -10, 14, 24, 13, -9, -14, -4,
    -- layer=1 filter=1 channel=44
    -47, -29, -32, -21, -2, 21, -8, -29, 5,
    -- layer=1 filter=1 channel=45
    -11, -32, -28, -26, 15, 1, 1, -4, 11,
    -- layer=1 filter=1 channel=46
    76, 73, 50, -5, -3, 0, 21, -14, 26,
    -- layer=1 filter=1 channel=47
    -42, -22, -41, -78, -52, -52, -9, -22, -25,
    -- layer=1 filter=1 channel=48
    -1, -9, 3, -5, 1, 0, 21, 20, 12,
    -- layer=1 filter=1 channel=49
    -10, -5, -8, -7, -18, -6, 21, 28, 8,
    -- layer=1 filter=1 channel=50
    -6, -21, -1, -5, -8, 0, -6, 7, -4,
    -- layer=1 filter=1 channel=51
    -16, -39, -15, -9, -46, -29, 30, 23, 24,
    -- layer=1 filter=1 channel=52
    4, 20, 10, 15, -3, 2, 10, 5, -2,
    -- layer=1 filter=1 channel=53
    6, 14, 7, 13, 12, 10, 9, 14, 21,
    -- layer=1 filter=1 channel=54
    -5, -7, -7, -28, -33, -38, -66, -68, 0,
    -- layer=1 filter=1 channel=55
    15, 10, 14, 3, 12, 21, -27, -6, -13,
    -- layer=1 filter=1 channel=56
    7, 10, -8, -3, 2, -5, -9, -9, 6,
    -- layer=1 filter=1 channel=57
    -36, -69, -19, -18, -43, -8, 11, 28, 36,
    -- layer=1 filter=1 channel=58
    -66, -86, -26, -120, -123, -103, -81, -93, -56,
    -- layer=1 filter=1 channel=59
    -12, -10, -4, -10, -3, -3, 2, -4, -3,
    -- layer=1 filter=1 channel=60
    12, 4, -6, 0, 16, 12, 18, 0, 0,
    -- layer=1 filter=1 channel=61
    8, 11, 4, 11, -1, 1, 5, 3, 0,
    -- layer=1 filter=1 channel=62
    13, 2, -3, -7, 33, 23, -25, -28, 26,
    -- layer=1 filter=1 channel=63
    16, 9, 5, 14, 11, 1, -17, -18, 0,
    -- layer=1 filter=1 channel=64
    -14, -19, -16, 9, -7, -13, 23, 24, 14,
    -- layer=1 filter=1 channel=65
    -10, -5, -8, -2, -7, -4, 14, 16, 14,
    -- layer=1 filter=1 channel=66
    1, 16, 17, -9, -3, 3, -10, -8, -8,
    -- layer=1 filter=1 channel=67
    -4, -4, -28, -14, -45, -24, 51, 27, 31,
    -- layer=1 filter=1 channel=68
    -60, -41, -41, -66, -27, -7, -50, -37, 18,
    -- layer=1 filter=1 channel=69
    2, 4, 3, -8, 29, 24, -9, -19, -9,
    -- layer=1 filter=1 channel=70
    -16, 9, -41, -44, -51, -18, 49, 29, 20,
    -- layer=1 filter=1 channel=71
    -1, -9, 0, -31, -9, 9, -28, -37, -35,
    -- layer=1 filter=1 channel=72
    52, 24, 8, 0, 0, -6, -8, -22, 39,
    -- layer=1 filter=1 channel=73
    10, 9, -5, -1, 0, 6, -7, -6, 2,
    -- layer=1 filter=1 channel=74
    -35, -3, -20, -2, -22, -12, 3, -1, 27,
    -- layer=1 filter=1 channel=75
    46, 45, 3, -2, -9, 0, -32, 10, 40,
    -- layer=1 filter=1 channel=76
    -2, -1, 4, 11, -4, 5, 2, 5, 9,
    -- layer=1 filter=1 channel=77
    -13, -23, -19, 2, -19, -7, -9, -16, -4,
    -- layer=1 filter=1 channel=78
    5, -11, -4, 11, -11, -9, -5, -7, -7,
    -- layer=1 filter=1 channel=79
    -6, 11, -9, 1, 28, 21, 0, -1, 30,
    -- layer=1 filter=1 channel=80
    -8, 9, -2, -4, 4, -2, 4, 5, 9,
    -- layer=1 filter=1 channel=81
    -7, -10, -23, 4, 13, -13, -37, -25, 0,
    -- layer=1 filter=1 channel=82
    -19, -15, -21, 2, -15, -9, 21, 19, 17,
    -- layer=1 filter=1 channel=83
    0, -14, 7, 5, 38, 1, 7, -17, 27,
    -- layer=1 filter=1 channel=84
    -33, -2, 13, -1, -28, -9, -11, 10, -2,
    -- layer=1 filter=1 channel=85
    -34, -77, -31, -90, -48, -60, -66, -106, -16,
    -- layer=1 filter=1 channel=86
    14, 18, 21, 12, 16, 12, -21, -19, -16,
    -- layer=1 filter=1 channel=87
    73, 60, 72, -23, -18, -43, 49, 2, 47,
    -- layer=1 filter=1 channel=88
    -9, -18, 14, 6, -10, 10, 17, 16, 21,
    -- layer=1 filter=1 channel=89
    -12, 1, -2, -6, -16, -1, 11, 16, 23,
    -- layer=1 filter=1 channel=90
    -31, -25, -32, -36, 0, -9, -38, -61, 9,
    -- layer=1 filter=1 channel=91
    -28, -24, -17, 16, 3, -8, 48, 33, 26,
    -- layer=1 filter=1 channel=92
    -2, 28, -3, -27, 5, 48, 62, 11, 1,
    -- layer=1 filter=1 channel=93
    7, -5, 0, -5, 4, 5, -2, 1, 3,
    -- layer=1 filter=1 channel=94
    13, 4, 3, 7, 3, 11, -14, 3, -7,
    -- layer=1 filter=1 channel=95
    -10, 12, 28, -14, -36, -14, -31, -9, 10,
    -- layer=1 filter=1 channel=96
    -6, -8, 6, 9, 2, 0, 2, 11, 15,
    -- layer=1 filter=1 channel=97
    1, -3, 1, 12, 5, -4, 4, 3, -5,
    -- layer=1 filter=1 channel=98
    11, -1, -8, 34, 30, 18, 7, 6, 24,
    -- layer=1 filter=1 channel=99
    -68, -77, 15, -67, -89, -107, -29, -26, -40,
    -- layer=1 filter=1 channel=100
    14, 13, 0, -2, -10, 11, -23, -15, -4,
    -- layer=1 filter=1 channel=101
    -16, -17, -11, 5, 2, -1, 21, 41, 15,
    -- layer=1 filter=1 channel=102
    -7, -10, -6, 12, 6, 0, 15, 19, -3,
    -- layer=1 filter=1 channel=103
    -8, -8, 0, 2, 4, -12, -3, -26, -4,
    -- layer=1 filter=1 channel=104
    -26, -14, -10, -45, -8, -15, -24, -26, -10,
    -- layer=1 filter=1 channel=105
    -1, 11, 21, 9, 8, -1, -4, 2, -1,
    -- layer=1 filter=1 channel=106
    -39, -30, -27, -3, -8, 1, 37, 29, 40,
    -- layer=1 filter=1 channel=107
    -2, 4, 9, -1, 5, 14, 1, 4, 2,
    -- layer=1 filter=1 channel=108
    -28, -40, -44, -47, -3, -7, -35, -72, -30,
    -- layer=1 filter=1 channel=109
    -3, 7, 2, 4, 0, 0, -5, -7, 2,
    -- layer=1 filter=1 channel=110
    -6, -6, 2, -3, 7, -6, -11, -8, -11,
    -- layer=1 filter=1 channel=111
    4, 14, 43, -13, -11, -9, -11, -1, -4,
    -- layer=1 filter=1 channel=112
    -12, 11, 50, -3, -17, 3, -4, 7, 2,
    -- layer=1 filter=1 channel=113
    -19, -45, -34, 10, -4, 2, 13, 8, 16,
    -- layer=1 filter=1 channel=114
    3, 27, 16, -9, 0, 5, -23, -31, -35,
    -- layer=1 filter=1 channel=115
    0, 0, 12, 5, -5, 9, -8, -3, -2,
    -- layer=1 filter=1 channel=116
    -2, -7, -7, -3, -10, 9, 9, 2, -3,
    -- layer=1 filter=1 channel=117
    12, 2, 86, 16, 2, 0, 9, 2, -9,
    -- layer=1 filter=1 channel=118
    -16, 10, 14, 2, -15, -11, 12, 10, 27,
    -- layer=1 filter=1 channel=119
    -25, -62, -55, -81, -42, -30, -45, -60, -1,
    -- layer=1 filter=1 channel=120
    -19, -35, -32, -16, -4, -13, 22, 13, 16,
    -- layer=1 filter=1 channel=121
    54, 67, 44, -10, 13, 18, -19, -22, -12,
    -- layer=1 filter=1 channel=122
    1, 3, -9, -4, -9, -5, 0, 6, 3,
    -- layer=1 filter=1 channel=123
    26, 28, 9, -8, 13, 7, -18, -11, -7,
    -- layer=1 filter=1 channel=124
    5, -6, -2, -4, 3, 13, 2, 1, 3,
    -- layer=1 filter=1 channel=125
    -40, -38, -51, -38, -52, -24, 45, 36, 36,
    -- layer=1 filter=1 channel=126
    16, 18, 16, 52, 55, 4, -4, 10, 33,
    -- layer=1 filter=1 channel=127
    13, 18, 32, -18, -21, -19, 4, 13, 15,
    -- layer=1 filter=2 channel=0
    0, -15, -3, -7, -4, -5, -19, -4, -9,
    -- layer=1 filter=2 channel=1
    -11, -10, -9, 3, 0, -7, -15, -19, -15,
    -- layer=1 filter=2 channel=2
    9, 1, 16, -12, 0, 1, -9, -10, 0,
    -- layer=1 filter=2 channel=3
    -10, -11, -7, -4, 4, -8, -10, -2, 6,
    -- layer=1 filter=2 channel=4
    5, 6, 3, -7, 5, 3, 1, -2, 5,
    -- layer=1 filter=2 channel=5
    13, -13, -16, 8, 0, -1, 0, 13, -8,
    -- layer=1 filter=2 channel=6
    -11, 0, 8, 9, -5, 3, 9, 0, -4,
    -- layer=1 filter=2 channel=7
    -5, -2, -21, -24, -15, -20, -10, -2, -7,
    -- layer=1 filter=2 channel=8
    -5, -14, -25, -10, -15, 0, -8, -6, 2,
    -- layer=1 filter=2 channel=9
    -17, -28, -21, -1, -10, -16, -11, -27, -13,
    -- layer=1 filter=2 channel=10
    -12, -11, -20, -12, -12, -24, -25, 2, -7,
    -- layer=1 filter=2 channel=11
    -21, -22, -18, -7, -18, -21, -21, -24, -19,
    -- layer=1 filter=2 channel=12
    6, -7, -14, -8, -8, -3, -1, -12, -4,
    -- layer=1 filter=2 channel=13
    17, 7, -4, 2, 13, -1, 4, -5, 15,
    -- layer=1 filter=2 channel=14
    0, -17, -3, -26, -16, -18, -18, -16, -15,
    -- layer=1 filter=2 channel=15
    16, -6, -11, -8, -2, 10, -9, 3, -5,
    -- layer=1 filter=2 channel=16
    -2, -7, -7, -5, 2, -8, 11, 11, 7,
    -- layer=1 filter=2 channel=17
    -20, -5, -10, -3, -8, -20, -4, -16, -14,
    -- layer=1 filter=2 channel=18
    -19, -31, -21, -6, -14, -17, -22, -11, 4,
    -- layer=1 filter=2 channel=19
    -22, -14, -14, -6, -17, -1, -18, -3, -4,
    -- layer=1 filter=2 channel=20
    0, 7, 2, 1, -4, 0, 4, 4, 6,
    -- layer=1 filter=2 channel=21
    1, -16, -11, 2, -1, 1, -17, -10, -9,
    -- layer=1 filter=2 channel=22
    16, 0, 5, 11, 8, 16, 11, 12, 15,
    -- layer=1 filter=2 channel=23
    -14, -12, -16, -20, -12, -19, -7, -10, -18,
    -- layer=1 filter=2 channel=24
    6, -7, -15, -3, -8, -14, -2, -5, 0,
    -- layer=1 filter=2 channel=25
    10, -2, -17, -23, -19, -7, -10, -6, -3,
    -- layer=1 filter=2 channel=26
    8, -21, -18, 2, -4, -15, -2, -13, -11,
    -- layer=1 filter=2 channel=27
    -1, -13, 5, 0, -18, -4, 4, -17, -8,
    -- layer=1 filter=2 channel=28
    -1, -14, -18, -22, -26, -18, -24, -2, -10,
    -- layer=1 filter=2 channel=29
    0, 7, 0, 5, 1, 6, -3, -4, -5,
    -- layer=1 filter=2 channel=30
    -10, -29, -13, -6, -5, -5, -9, -23, -16,
    -- layer=1 filter=2 channel=31
    2, 0, 10, 1, -7, -7, 17, -3, -4,
    -- layer=1 filter=2 channel=32
    8, -8, -11, 4, -26, -20, 0, -21, -7,
    -- layer=1 filter=2 channel=33
    2, -9, 9, 15, 10, 18, 6, 4, 9,
    -- layer=1 filter=2 channel=34
    13, 8, 7, 18, 3, 3, 3, 11, 11,
    -- layer=1 filter=2 channel=35
    -5, -8, -3, 3, -8, 8, -3, -6, -3,
    -- layer=1 filter=2 channel=36
    -26, -30, -26, -18, -24, -23, -5, -14, -29,
    -- layer=1 filter=2 channel=37
    0, -4, -10, -17, 0, 8, 8, 10, -5,
    -- layer=1 filter=2 channel=38
    -1, -2, 7, -2, 11, -5, 0, -1, 12,
    -- layer=1 filter=2 channel=39
    -10, 3, -10, 3, -9, -9, -15, -16, -15,
    -- layer=1 filter=2 channel=40
    5, -11, 5, 9, 0, -2, 8, 2, -4,
    -- layer=1 filter=2 channel=41
    -5, -21, -18, 0, -14, -2, -14, -23, -14,
    -- layer=1 filter=2 channel=42
    0, 6, 17, -4, 0, 8, 4, -17, -1,
    -- layer=1 filter=2 channel=43
    0, -17, -22, -17, -14, 0, -17, -12, -4,
    -- layer=1 filter=2 channel=44
    -2, -16, -21, -5, -8, -19, -11, -6, -1,
    -- layer=1 filter=2 channel=45
    18, -3, -12, 2, -11, -9, -5, -9, -10,
    -- layer=1 filter=2 channel=46
    -8, -16, -6, 8, 17, -2, 6, 11, 9,
    -- layer=1 filter=2 channel=47
    -5, -16, -28, 1, -23, 0, -20, -11, 9,
    -- layer=1 filter=2 channel=48
    -2, -7, -5, -6, -3, -2, 0, -5, -4,
    -- layer=1 filter=2 channel=49
    8, -5, 10, -3, -6, -21, -1, -5, -6,
    -- layer=1 filter=2 channel=50
    -5, 5, 5, -10, -3, -6, 6, -11, -1,
    -- layer=1 filter=2 channel=51
    -12, 4, -12, 1, -13, -17, 1, -2, -5,
    -- layer=1 filter=2 channel=52
    2, -8, 2, -9, -7, -10, -8, 10, 6,
    -- layer=1 filter=2 channel=53
    -6, -10, -13, -2, -1, 6, 7, -6, 6,
    -- layer=1 filter=2 channel=54
    -14, -20, -20, -23, -16, -3, -11, 6, -14,
    -- layer=1 filter=2 channel=55
    1, 0, -6, -14, -7, -3, -10, -6, 5,
    -- layer=1 filter=2 channel=56
    -6, 2, -6, -6, 0, 0, -10, -3, -6,
    -- layer=1 filter=2 channel=57
    -7, -11, -24, 0, -10, -6, 2, 3, -19,
    -- layer=1 filter=2 channel=58
    -18, -36, -24, 6, -17, -24, 0, 0, -19,
    -- layer=1 filter=2 channel=59
    2, -5, 2, -1, 2, 7, -3, 6, -9,
    -- layer=1 filter=2 channel=60
    -5, -6, -2, 9, 11, -3, -1, -11, -8,
    -- layer=1 filter=2 channel=61
    -5, 1, -2, -5, -11, 9, 5, -7, 0,
    -- layer=1 filter=2 channel=62
    7, -13, -18, 4, -2, 5, 6, 6, -8,
    -- layer=1 filter=2 channel=63
    -9, -25, -29, -18, -16, -14, -18, -20, -26,
    -- layer=1 filter=2 channel=64
    -10, -5, -9, -5, -15, -12, -11, -15, 0,
    -- layer=1 filter=2 channel=65
    -13, -13, -16, 0, -8, -4, -14, -13, -15,
    -- layer=1 filter=2 channel=66
    -18, -19, -8, -5, -13, -12, -22, -28, -9,
    -- layer=1 filter=2 channel=67
    -15, -10, -16, -2, -13, -22, -3, -21, -3,
    -- layer=1 filter=2 channel=68
    10, -25, 2, -7, -11, -13, -8, -15, -1,
    -- layer=1 filter=2 channel=69
    18, -26, -12, 6, -2, 18, -1, 2, 10,
    -- layer=1 filter=2 channel=70
    9, 0, 10, 12, -1, 8, 4, 7, 3,
    -- layer=1 filter=2 channel=71
    -16, -8, -1, -20, 0, 0, -4, -1, -3,
    -- layer=1 filter=2 channel=72
    -15, -29, -13, -5, -14, -10, -14, -1, -1,
    -- layer=1 filter=2 channel=73
    3, -2, 3, -7, 4, 5, -10, 0, 0,
    -- layer=1 filter=2 channel=74
    6, -1, -11, -4, -12, -4, -2, -4, -9,
    -- layer=1 filter=2 channel=75
    -16, -25, -7, -11, -16, -6, -16, -10, 10,
    -- layer=1 filter=2 channel=76
    -10, -14, -15, 0, -15, -20, -6, 0, -12,
    -- layer=1 filter=2 channel=77
    -5, -4, -8, -6, -10, -2, -10, -22, -10,
    -- layer=1 filter=2 channel=78
    -7, 3, 4, -6, -1, -8, -6, 5, 0,
    -- layer=1 filter=2 channel=79
    7, -8, -4, -9, -5, 10, -1, 2, -11,
    -- layer=1 filter=2 channel=80
    -5, -13, -4, -5, -8, -4, -4, -3, -5,
    -- layer=1 filter=2 channel=81
    -17, -9, -17, -7, -20, -14, -7, -8, -1,
    -- layer=1 filter=2 channel=82
    -15, 0, 2, -15, -16, -12, -4, -13, -8,
    -- layer=1 filter=2 channel=83
    0, -2, -8, -9, -4, -1, 0, -3, -10,
    -- layer=1 filter=2 channel=84
    3, -21, -14, -4, -15, -16, -6, -12, -17,
    -- layer=1 filter=2 channel=85
    -11, -21, -16, -1, -23, -14, -20, -6, -25,
    -- layer=1 filter=2 channel=86
    -24, -17, -19, -19, -17, -6, -16, -6, -2,
    -- layer=1 filter=2 channel=87
    -3, -8, -10, -1, -3, -16, -11, 11, -10,
    -- layer=1 filter=2 channel=88
    -9, -2, -12, -17, -6, -18, -20, -8, -9,
    -- layer=1 filter=2 channel=89
    2, -17, 0, -5, -13, -17, -17, -11, -14,
    -- layer=1 filter=2 channel=90
    -13, -30, -11, -3, -8, -3, -7, -12, -18,
    -- layer=1 filter=2 channel=91
    -6, 0, 6, 0, 1, -5, -3, 5, 8,
    -- layer=1 filter=2 channel=92
    0, -25, -13, -15, -14, -8, -23, -18, -15,
    -- layer=1 filter=2 channel=93
    -16, -10, -1, -13, -5, 1, -13, -14, -11,
    -- layer=1 filter=2 channel=94
    -24, -14, -21, -14, -7, -9, -19, -3, -23,
    -- layer=1 filter=2 channel=95
    -20, -12, -25, -14, -6, -1, -12, -15, -12,
    -- layer=1 filter=2 channel=96
    -7, 4, 7, -2, -13, -12, 0, -10, 0,
    -- layer=1 filter=2 channel=97
    -12, -12, -24, -20, -8, -8, -11, -14, -24,
    -- layer=1 filter=2 channel=98
    -6, -5, -15, -18, -7, -5, 3, 2, 1,
    -- layer=1 filter=2 channel=99
    -11, -15, -23, -23, -13, -17, -15, -12, -14,
    -- layer=1 filter=2 channel=100
    -7, -4, -7, -21, -9, -13, -1, -1, -4,
    -- layer=1 filter=2 channel=101
    5, 7, -8, 6, -6, 0, -4, -10, -6,
    -- layer=1 filter=2 channel=102
    -16, -14, -6, -18, -2, -15, -8, -8, -5,
    -- layer=1 filter=2 channel=103
    -8, -11, -5, -9, -19, 2, -3, -11, -7,
    -- layer=1 filter=2 channel=104
    -14, 3, -3, -10, -15, 3, -1, -12, 1,
    -- layer=1 filter=2 channel=105
    -11, -10, -28, -17, -10, -23, -17, -15, -19,
    -- layer=1 filter=2 channel=106
    -1, 5, -3, -5, -7, -12, -9, -5, 3,
    -- layer=1 filter=2 channel=107
    -2, 4, 0, -2, -10, -4, -1, -11, 5,
    -- layer=1 filter=2 channel=108
    7, -4, -7, 1, -8, -14, -9, -9, 1,
    -- layer=1 filter=2 channel=109
    4, -1, -1, -4, 7, -8, 7, -2, -1,
    -- layer=1 filter=2 channel=110
    4, 3, 5, -12, 4, -11, 3, 2, -10,
    -- layer=1 filter=2 channel=111
    -7, -6, -18, -8, -16, -13, -25, -26, -8,
    -- layer=1 filter=2 channel=112
    -3, -19, -20, -17, -2, 1, -5, -9, -5,
    -- layer=1 filter=2 channel=113
    15, 13, 16, 0, -1, 13, 4, 5, -7,
    -- layer=1 filter=2 channel=114
    8, -16, -3, 6, 15, -10, 5, 12, -1,
    -- layer=1 filter=2 channel=115
    -17, -20, -16, -25, -17, -25, -14, -2, -17,
    -- layer=1 filter=2 channel=116
    -4, 8, -10, -5, 5, -7, -11, 7, -5,
    -- layer=1 filter=2 channel=117
    0, -6, -12, -18, 0, -16, -12, -4, -13,
    -- layer=1 filter=2 channel=118
    -1, -27, -2, -14, -14, -12, -9, -18, -20,
    -- layer=1 filter=2 channel=119
    4, -20, -2, 0, -20, -18, 6, -23, -17,
    -- layer=1 filter=2 channel=120
    5, -7, -9, -10, -10, -17, -12, -10, -9,
    -- layer=1 filter=2 channel=121
    -18, -20, -23, -7, -4, -4, -16, -5, -3,
    -- layer=1 filter=2 channel=122
    -1, 4, 6, -1, 0, 8, 4, -5, 10,
    -- layer=1 filter=2 channel=123
    -22, -13, -8, -15, -6, -9, 2, -1, -9,
    -- layer=1 filter=2 channel=124
    -10, 0, 0, -7, -6, 6, 6, 2, -2,
    -- layer=1 filter=2 channel=125
    15, -8, 7, -3, 1, -7, 7, 17, 13,
    -- layer=1 filter=2 channel=126
    4, -18, -7, -15, -7, -16, -4, -12, -5,
    -- layer=1 filter=2 channel=127
    -7, -23, -16, -14, -11, -8, -19, -20, -13,
    -- layer=1 filter=3 channel=0
    8, -3, 0, -6, 0, 0, -10, -10, 3,
    -- layer=1 filter=3 channel=1
    3, 0, 5, -8, -9, 2, -10, -4, 4,
    -- layer=1 filter=3 channel=2
    -3, -16, 3, 3, -14, -3, -6, 5, 1,
    -- layer=1 filter=3 channel=3
    -7, -7, -5, -4, 1, 8, -7, 0, -3,
    -- layer=1 filter=3 channel=4
    -9, 4, 7, -6, 3, 1, 0, -4, -4,
    -- layer=1 filter=3 channel=5
    -6, -2, 1, 4, -11, 2, -6, -5, -5,
    -- layer=1 filter=3 channel=6
    6, -6, -2, -8, 4, -4, -7, 5, -2,
    -- layer=1 filter=3 channel=7
    -13, 6, -5, 0, 0, -7, -13, 2, -3,
    -- layer=1 filter=3 channel=8
    0, -9, -5, 8, -7, -3, 5, -2, -9,
    -- layer=1 filter=3 channel=9
    1, -9, 4, 7, -2, -6, -1, 0, -5,
    -- layer=1 filter=3 channel=10
    5, 7, -11, -3, -7, -4, -11, -12, 0,
    -- layer=1 filter=3 channel=11
    -1, 8, 5, -6, 0, -12, 6, 2, -2,
    -- layer=1 filter=3 channel=12
    3, -3, 10, 8, -5, 0, 3, -4, 0,
    -- layer=1 filter=3 channel=13
    -9, -6, -9, -3, 4, 7, -7, -9, 3,
    -- layer=1 filter=3 channel=14
    -8, -5, -8, -1, -8, -5, 1, -8, 0,
    -- layer=1 filter=3 channel=15
    3, -2, -1, -9, 1, 6, -7, -7, 9,
    -- layer=1 filter=3 channel=16
    12, -8, -7, -7, -1, -3, -7, -6, 6,
    -- layer=1 filter=3 channel=17
    -3, 7, 2, 8, -4, -2, -8, -9, 7,
    -- layer=1 filter=3 channel=18
    -6, 2, -9, -9, -7, -10, 7, 8, 0,
    -- layer=1 filter=3 channel=19
    6, 8, -11, -3, -5, 4, 1, -1, 7,
    -- layer=1 filter=3 channel=20
    -8, 6, -5, 1, 0, -9, -4, -10, -2,
    -- layer=1 filter=3 channel=21
    1, -12, 5, -7, 4, 1, 0, 0, -3,
    -- layer=1 filter=3 channel=22
    -3, 6, -12, 2, -11, -2, 5, -6, -3,
    -- layer=1 filter=3 channel=23
    6, -1, -4, 5, 1, -8, 7, 9, -1,
    -- layer=1 filter=3 channel=24
    4, -7, 4, 2, -8, 5, -9, -10, 6,
    -- layer=1 filter=3 channel=25
    4, 4, 5, 3, -13, 0, 0, 2, 8,
    -- layer=1 filter=3 channel=26
    -10, -11, -11, 2, -4, -1, -8, 4, 0,
    -- layer=1 filter=3 channel=27
    -3, -2, 7, -6, 5, -7, 3, 1, -7,
    -- layer=1 filter=3 channel=28
    -8, -11, -13, -7, -9, -5, 7, -12, 6,
    -- layer=1 filter=3 channel=29
    11, 11, 8, -5, 6, 6, -11, 3, 0,
    -- layer=1 filter=3 channel=30
    -8, 6, -3, -11, 9, -10, -8, -4, -9,
    -- layer=1 filter=3 channel=31
    4, 0, 1, -4, -8, 1, -1, -4, 0,
    -- layer=1 filter=3 channel=32
    1, 4, -7, 2, 5, -9, -4, 1, 8,
    -- layer=1 filter=3 channel=33
    2, 5, -2, -8, 7, -3, 0, -5, -2,
    -- layer=1 filter=3 channel=34
    8, 7, -11, 5, -6, -11, 6, 8, -8,
    -- layer=1 filter=3 channel=35
    0, 1, -9, -8, 7, 8, 2, 10, 8,
    -- layer=1 filter=3 channel=36
    2, 9, 3, 0, 9, -2, -10, -4, -2,
    -- layer=1 filter=3 channel=37
    0, -12, -10, -1, -3, -5, -9, 0, -6,
    -- layer=1 filter=3 channel=38
    -9, -1, -11, -3, 6, 6, -11, -6, 3,
    -- layer=1 filter=3 channel=39
    6, 2, -8, 6, -7, -2, 3, 6, 2,
    -- layer=1 filter=3 channel=40
    -12, -9, 7, 0, 5, -2, -1, 2, 5,
    -- layer=1 filter=3 channel=41
    0, 0, -1, 0, 1, 9, -8, 4, 7,
    -- layer=1 filter=3 channel=42
    -3, -7, 0, -10, 5, 0, 7, -4, -10,
    -- layer=1 filter=3 channel=43
    5, 3, -6, 7, 3, 3, 7, 0, -12,
    -- layer=1 filter=3 channel=44
    -11, 0, -2, 7, 5, 7, 4, -7, -3,
    -- layer=1 filter=3 channel=45
    2, -3, -3, 3, -12, 0, 8, -7, -4,
    -- layer=1 filter=3 channel=46
    0, 4, -2, 0, -9, 0, -10, 8, 7,
    -- layer=1 filter=3 channel=47
    -1, -11, -11, 10, -7, -12, -8, -6, -5,
    -- layer=1 filter=3 channel=48
    -11, -9, -9, 0, 4, 3, 0, -6, 5,
    -- layer=1 filter=3 channel=49
    -3, 7, 5, -4, 2, 7, 4, -5, -5,
    -- layer=1 filter=3 channel=50
    -7, 2, 9, -8, -3, 8, 4, 3, -11,
    -- layer=1 filter=3 channel=51
    6, -7, 0, 7, -5, 4, 0, -6, -1,
    -- layer=1 filter=3 channel=52
    0, 9, -7, 1, -4, 7, 3, -11, -13,
    -- layer=1 filter=3 channel=53
    6, 0, 2, 2, 6, -1, -9, -7, -4,
    -- layer=1 filter=3 channel=54
    5, -4, -9, 5, -8, -6, -5, 0, 0,
    -- layer=1 filter=3 channel=55
    -11, -7, 2, 0, 3, -8, 6, 2, -9,
    -- layer=1 filter=3 channel=56
    5, 8, -1, 2, 8, 1, 3, -8, 5,
    -- layer=1 filter=3 channel=57
    0, -1, 0, -10, -3, 2, -5, -2, 1,
    -- layer=1 filter=3 channel=58
    -14, -13, 1, -2, 0, 8, 0, 0, -10,
    -- layer=1 filter=3 channel=59
    9, -8, -10, 5, -8, -8, -9, -2, 1,
    -- layer=1 filter=3 channel=60
    -2, 5, 0, 6, -4, 3, 2, 10, 1,
    -- layer=1 filter=3 channel=61
    -10, 6, 7, 0, -7, -2, 4, 1, 5,
    -- layer=1 filter=3 channel=62
    -7, -2, 0, 0, 5, -8, 0, 7, -8,
    -- layer=1 filter=3 channel=63
    1, -8, -5, -4, -1, 1, -10, 1, -9,
    -- layer=1 filter=3 channel=64
    0, -8, -4, -5, -12, -6, -12, -4, 5,
    -- layer=1 filter=3 channel=65
    -3, -11, 0, -6, 7, -9, 7, 2, 7,
    -- layer=1 filter=3 channel=66
    -10, -2, -10, -9, -9, 0, 5, -10, -13,
    -- layer=1 filter=3 channel=67
    0, -7, 11, -2, -7, 5, 7, 0, -1,
    -- layer=1 filter=3 channel=68
    -3, -4, -3, -7, 2, 1, -11, -5, -2,
    -- layer=1 filter=3 channel=69
    6, 0, 6, 2, -5, 0, -1, -3, 2,
    -- layer=1 filter=3 channel=70
    3, -1, 9, 0, -2, -3, 0, -6, -10,
    -- layer=1 filter=3 channel=71
    7, 1, 7, 9, -11, -3, 0, 0, 8,
    -- layer=1 filter=3 channel=72
    -4, -1, 4, 9, 3, 1, 0, -2, -4,
    -- layer=1 filter=3 channel=73
    -5, 3, -2, 3, -5, 0, 5, -6, 5,
    -- layer=1 filter=3 channel=74
    -10, -5, 6, 5, 1, 8, -5, 5, 7,
    -- layer=1 filter=3 channel=75
    0, -4, -6, 2, -3, 4, -1, 0, 6,
    -- layer=1 filter=3 channel=76
    0, 4, -11, 5, -2, 6, -5, 6, -11,
    -- layer=1 filter=3 channel=77
    -3, 0, 2, -9, 5, -5, -2, 1, -10,
    -- layer=1 filter=3 channel=78
    3, -8, 0, -8, 0, 2, 6, -2, -5,
    -- layer=1 filter=3 channel=79
    -8, -11, 7, 4, -4, 8, 8, 4, 1,
    -- layer=1 filter=3 channel=80
    -4, 7, -1, -5, 0, -6, -5, -5, 1,
    -- layer=1 filter=3 channel=81
    5, -7, 1, -11, 4, 5, -5, -3, -2,
    -- layer=1 filter=3 channel=82
    2, 4, 0, -4, 6, 0, -3, 7, 5,
    -- layer=1 filter=3 channel=83
    -5, 4, -10, -5, -9, 0, -10, 7, -9,
    -- layer=1 filter=3 channel=84
    0, -6, 0, 0, 5, 4, 0, -9, -3,
    -- layer=1 filter=3 channel=85
    2, -8, 4, 0, -1, 4, -9, 4, -12,
    -- layer=1 filter=3 channel=86
    2, 0, -6, -12, 4, -5, -2, -2, -3,
    -- layer=1 filter=3 channel=87
    -3, 5, -7, 8, -7, 6, 7, 0, -5,
    -- layer=1 filter=3 channel=88
    0, 5, -3, -2, -2, -7, -2, -13, -6,
    -- layer=1 filter=3 channel=89
    -7, -1, 0, 0, -10, 7, 8, -12, -8,
    -- layer=1 filter=3 channel=90
    -5, -2, 0, 2, 6, 5, -8, -2, 5,
    -- layer=1 filter=3 channel=91
    1, -5, 3, -12, -9, -2, -7, -6, -11,
    -- layer=1 filter=3 channel=92
    0, 1, 2, 2, 0, -2, 6, 8, 6,
    -- layer=1 filter=3 channel=93
    6, -2, -5, 5, 7, -4, 6, 2, 4,
    -- layer=1 filter=3 channel=94
    3, -8, 4, -4, -8, 2, 0, -4, 0,
    -- layer=1 filter=3 channel=95
    2, -4, -2, 7, -6, -5, 8, 6, -4,
    -- layer=1 filter=3 channel=96
    6, 1, -8, 0, -3, -1, 0, 2, -2,
    -- layer=1 filter=3 channel=97
    -1, 8, -11, -6, -2, -9, 7, -8, -5,
    -- layer=1 filter=3 channel=98
    2, -9, -3, -10, 1, 0, -6, 0, 1,
    -- layer=1 filter=3 channel=99
    4, 4, 7, -6, 2, -10, 1, -3, 3,
    -- layer=1 filter=3 channel=100
    8, 6, -10, 1, 7, 8, -4, -5, -10,
    -- layer=1 filter=3 channel=101
    -11, -10, -4, 0, 1, 5, 8, 4, -7,
    -- layer=1 filter=3 channel=102
    5, 1, -5, 5, 6, 2, -1, 4, 4,
    -- layer=1 filter=3 channel=103
    -11, 1, -1, -9, -9, 4, -7, 5, 0,
    -- layer=1 filter=3 channel=104
    -9, 9, 9, 1, -2, 0, -8, -6, 0,
    -- layer=1 filter=3 channel=105
    -6, 8, -7, -8, 2, 5, -9, -5, 4,
    -- layer=1 filter=3 channel=106
    2, 3, 6, 2, 1, -6, -10, -7, -7,
    -- layer=1 filter=3 channel=107
    -8, -4, 0, -8, 1, 4, 7, -8, 1,
    -- layer=1 filter=3 channel=108
    5, 3, 4, -9, -8, 2, 3, -5, 5,
    -- layer=1 filter=3 channel=109
    -9, -4, 9, 3, 2, -11, 0, -8, 7,
    -- layer=1 filter=3 channel=110
    9, -6, 2, -1, 5, -1, -4, 7, -12,
    -- layer=1 filter=3 channel=111
    -6, -7, 9, 1, -10, -6, -8, 3, 8,
    -- layer=1 filter=3 channel=112
    6, -4, -3, 1, 4, -6, 2, 0, 4,
    -- layer=1 filter=3 channel=113
    2, 2, -4, -5, -4, -8, 5, 0, 7,
    -- layer=1 filter=3 channel=114
    -6, -1, -10, 5, 0, 8, 3, 2, 7,
    -- layer=1 filter=3 channel=115
    -8, -3, 7, -3, -1, -1, -9, -11, 5,
    -- layer=1 filter=3 channel=116
    -2, -4, 8, 10, 6, 0, 2, 0, 7,
    -- layer=1 filter=3 channel=117
    -4, 8, 0, -2, 0, 2, -1, 2, 8,
    -- layer=1 filter=3 channel=118
    5, -6, 7, 1, -12, -10, 4, -4, -5,
    -- layer=1 filter=3 channel=119
    -11, -5, 5, -2, -3, -8, 1, -13, -11,
    -- layer=1 filter=3 channel=120
    -5, -10, -6, 5, -1, -6, -10, -4, -2,
    -- layer=1 filter=3 channel=121
    -3, -3, -8, 0, -2, -8, -2, -6, -6,
    -- layer=1 filter=3 channel=122
    -3, 6, 8, -9, -2, -1, -1, -9, 2,
    -- layer=1 filter=3 channel=123
    0, 2, 0, 2, 5, 0, -4, 7, 0,
    -- layer=1 filter=3 channel=124
    1, -8, -1, 9, -5, -5, -7, 0, -3,
    -- layer=1 filter=3 channel=125
    -8, -1, -8, -1, -1, -10, 4, -3, -9,
    -- layer=1 filter=3 channel=126
    -5, 1, -5, -1, -6, -9, -2, 3, -2,
    -- layer=1 filter=3 channel=127
    -3, 5, -2, -10, -1, 2, 0, 10, 0,
    -- layer=1 filter=4 channel=0
    -6, -7, -2, 3, 0, 2, 2, -1, -4,
    -- layer=1 filter=4 channel=1
    -8, 8, 3, -10, -1, -1, 0, 3, -3,
    -- layer=1 filter=4 channel=2
    3, -3, 4, -7, -5, 3, -1, 8, 0,
    -- layer=1 filter=4 channel=3
    -3, 9, -8, 4, -4, -8, -2, -6, -4,
    -- layer=1 filter=4 channel=4
    3, -6, -3, 5, -8, -7, -4, 0, 8,
    -- layer=1 filter=4 channel=5
    0, -5, -3, -11, 5, -11, 2, 7, 0,
    -- layer=1 filter=4 channel=6
    -3, 7, 3, -1, 5, -4, -13, 9, -1,
    -- layer=1 filter=4 channel=7
    -5, 3, -5, -14, 7, -9, -2, -4, 1,
    -- layer=1 filter=4 channel=8
    -5, -3, -3, -7, -7, 4, 2, -3, -1,
    -- layer=1 filter=4 channel=9
    6, 0, 6, -6, 1, -13, -7, -5, -1,
    -- layer=1 filter=4 channel=10
    -13, -2, -9, -1, 0, 1, 1, -3, 6,
    -- layer=1 filter=4 channel=11
    -11, 0, -11, -6, 0, -15, -3, -2, -5,
    -- layer=1 filter=4 channel=12
    -9, -7, 3, -1, 1, -8, -5, -1, 8,
    -- layer=1 filter=4 channel=13
    -11, -3, 3, -3, 2, -5, -7, 0, 4,
    -- layer=1 filter=4 channel=14
    -9, -4, 0, 5, -12, -9, -9, 10, 5,
    -- layer=1 filter=4 channel=15
    -4, -2, 1, -1, -9, -8, -9, 11, -5,
    -- layer=1 filter=4 channel=16
    2, -11, -9, -12, 2, 8, -1, 10, 0,
    -- layer=1 filter=4 channel=17
    -9, 4, -1, -13, -2, 7, 2, 5, -8,
    -- layer=1 filter=4 channel=18
    0, 2, -11, -1, -5, -7, 0, -2, -13,
    -- layer=1 filter=4 channel=19
    0, -13, -11, -11, -3, 4, 0, -4, -2,
    -- layer=1 filter=4 channel=20
    1, -14, -11, -15, -1, -7, -6, -9, 4,
    -- layer=1 filter=4 channel=21
    -5, 1, -5, -16, 0, 4, -9, 3, 0,
    -- layer=1 filter=4 channel=22
    -1, 0, -9, -5, 4, 1, 2, 0, 9,
    -- layer=1 filter=4 channel=23
    -1, -5, -4, 5, 0, -9, -5, -8, -5,
    -- layer=1 filter=4 channel=24
    -11, 1, -2, -9, -3, 3, -1, 2, 1,
    -- layer=1 filter=4 channel=25
    -5, -12, -7, 5, 8, 1, -5, -7, -4,
    -- layer=1 filter=4 channel=26
    -11, -15, -9, 0, -6, -10, 4, 2, 1,
    -- layer=1 filter=4 channel=27
    0, -10, 4, -4, 0, -5, -6, -4, 6,
    -- layer=1 filter=4 channel=28
    7, -3, 3, -3, -2, 7, 3, 6, 1,
    -- layer=1 filter=4 channel=29
    6, 4, 2, -7, 1, -11, -10, -1, -9,
    -- layer=1 filter=4 channel=30
    2, -9, 0, 5, -8, -11, 4, 1, 3,
    -- layer=1 filter=4 channel=31
    -2, 6, 7, 3, -7, -1, 2, 6, 1,
    -- layer=1 filter=4 channel=32
    -13, 1, -5, 1, -12, 0, 2, 4, -13,
    -- layer=1 filter=4 channel=33
    10, 8, 8, 3, 1, -7, 3, 0, 4,
    -- layer=1 filter=4 channel=34
    0, -3, -1, -11, 2, -11, 0, -11, 3,
    -- layer=1 filter=4 channel=35
    -5, -6, -3, -6, -5, 1, -1, 3, -11,
    -- layer=1 filter=4 channel=36
    -13, 1, -11, 4, 4, 4, -10, -1, -5,
    -- layer=1 filter=4 channel=37
    -14, -17, -12, -2, -7, 0, -9, -3, 0,
    -- layer=1 filter=4 channel=38
    0, -7, -10, 0, 2, -5, -9, 3, -7,
    -- layer=1 filter=4 channel=39
    -10, -4, -12, -6, -5, 0, -2, 0, 1,
    -- layer=1 filter=4 channel=40
    -7, -5, 8, 0, 4, -10, -6, -7, -4,
    -- layer=1 filter=4 channel=41
    -9, 4, -2, -1, 3, -7, 6, 2, -9,
    -- layer=1 filter=4 channel=42
    -10, 3, 5, -5, -5, -12, 6, -9, 1,
    -- layer=1 filter=4 channel=43
    -5, 3, -3, 4, -1, -4, -8, -4, 0,
    -- layer=1 filter=4 channel=44
    -16, -3, -8, -1, -2, -1, -2, -4, 1,
    -- layer=1 filter=4 channel=45
    -12, -3, -13, -2, -3, 0, -7, -2, -11,
    -- layer=1 filter=4 channel=46
    6, -14, -6, 1, -6, -2, -4, -7, 6,
    -- layer=1 filter=4 channel=47
    5, 5, 1, 6, 0, 3, 6, 4, -11,
    -- layer=1 filter=4 channel=48
    -6, -3, 0, 8, 8, -4, -4, 8, 2,
    -- layer=1 filter=4 channel=49
    -6, 7, -9, -3, 10, -4, -11, -11, 0,
    -- layer=1 filter=4 channel=50
    -4, 1, 0, 8, 6, 1, 4, -1, -4,
    -- layer=1 filter=4 channel=51
    -12, 9, 6, -5, 7, -7, -10, 3, -7,
    -- layer=1 filter=4 channel=52
    1, 8, -6, 0, -4, 7, 5, 3, -7,
    -- layer=1 filter=4 channel=53
    7, -4, -10, -7, 4, -5, -11, -10, 10,
    -- layer=1 filter=4 channel=54
    -7, 1, -3, 4, 6, 5, 3, 2, -2,
    -- layer=1 filter=4 channel=55
    -6, -9, -13, 6, -3, -12, 7, 5, -15,
    -- layer=1 filter=4 channel=56
    0, 5, 10, -7, 8, 7, 6, -3, 5,
    -- layer=1 filter=4 channel=57
    -13, 6, 3, -8, 5, -4, -2, 9, 5,
    -- layer=1 filter=4 channel=58
    -13, -14, -3, 3, 10, -4, 5, -6, 0,
    -- layer=1 filter=4 channel=59
    -10, 7, 0, -2, 0, 2, -5, 1, -1,
    -- layer=1 filter=4 channel=60
    -5, 0, -1, 0, -3, 3, -9, 3, 6,
    -- layer=1 filter=4 channel=61
    1, 2, -5, 8, 0, -2, 1, -4, 0,
    -- layer=1 filter=4 channel=62
    -3, -18, -3, -4, -5, 8, 11, -7, -18,
    -- layer=1 filter=4 channel=63
    -11, -1, -3, -2, -9, -9, -4, -1, -3,
    -- layer=1 filter=4 channel=64
    0, 0, -10, 6, -10, -5, -4, -7, 8,
    -- layer=1 filter=4 channel=65
    -4, 5, -10, -3, 7, 0, 2, -1, -9,
    -- layer=1 filter=4 channel=66
    -14, -6, -6, -9, 4, -7, 4, -11, -8,
    -- layer=1 filter=4 channel=67
    -8, 12, -2, 2, -5, 4, -1, -8, 5,
    -- layer=1 filter=4 channel=68
    -1, -10, 0, 2, -11, 0, 0, 3, 5,
    -- layer=1 filter=4 channel=69
    -13, -6, -1, 0, 0, -13, 0, -8, -4,
    -- layer=1 filter=4 channel=70
    0, 9, 6, -5, 11, 0, 0, -4, 5,
    -- layer=1 filter=4 channel=71
    -3, -4, -5, -12, -3, 0, 4, 3, -12,
    -- layer=1 filter=4 channel=72
    7, 5, -4, 9, -4, -6, -2, -10, 5,
    -- layer=1 filter=4 channel=73
    -6, -9, -1, 8, 7, 3, 0, -2, 1,
    -- layer=1 filter=4 channel=74
    -6, -3, -10, -9, 0, -10, 4, 0, 7,
    -- layer=1 filter=4 channel=75
    6, -2, 0, 0, -3, -5, -2, -10, -10,
    -- layer=1 filter=4 channel=76
    -4, -3, 7, 7, -5, 4, -15, -10, -6,
    -- layer=1 filter=4 channel=77
    -6, -8, 1, -11, -5, 9, 8, -3, 2,
    -- layer=1 filter=4 channel=78
    -5, -5, 1, 5, -8, -5, -1, -7, -6,
    -- layer=1 filter=4 channel=79
    -8, -1, -12, 7, -2, 1, 0, 0, 4,
    -- layer=1 filter=4 channel=80
    -6, 10, 0, -5, -7, 4, 2, -7, -1,
    -- layer=1 filter=4 channel=81
    -4, -12, 2, -10, 5, -8, 2, -2, -5,
    -- layer=1 filter=4 channel=82
    -12, -8, 10, -10, -3, -2, 0, -7, -3,
    -- layer=1 filter=4 channel=83
    4, -4, -7, -12, 0, -5, -5, 6, -4,
    -- layer=1 filter=4 channel=84
    1, 1, -5, -14, -10, 2, -4, -14, 4,
    -- layer=1 filter=4 channel=85
    -3, -3, 0, -2, 0, -7, 5, -12, -15,
    -- layer=1 filter=4 channel=86
    1, -13, -1, -1, -1, -13, 3, -12, -9,
    -- layer=1 filter=4 channel=87
    -7, 5, -10, -3, 0, 2, -3, 7, -8,
    -- layer=1 filter=4 channel=88
    -7, -9, -3, 5, 6, -12, -3, 0, 5,
    -- layer=1 filter=4 channel=89
    -8, 0, -10, -10, -15, -6, 0, -5, 5,
    -- layer=1 filter=4 channel=90
    -3, 6, 3, -2, -6, 6, -13, 0, -6,
    -- layer=1 filter=4 channel=91
    -7, -7, 1, -8, -2, 5, -3, 1, -7,
    -- layer=1 filter=4 channel=92
    6, 1, -7, -7, -10, 0, -5, 10, -5,
    -- layer=1 filter=4 channel=93
    3, 1, 2, -1, -5, 0, -2, 2, 5,
    -- layer=1 filter=4 channel=94
    0, -9, -9, -7, -2, 3, -1, -1, -10,
    -- layer=1 filter=4 channel=95
    -11, 1, -4, -10, 5, -8, 0, -8, -1,
    -- layer=1 filter=4 channel=96
    4, 1, -3, -4, 1, -6, -1, 0, -1,
    -- layer=1 filter=4 channel=97
    -1, -8, 5, -2, -6, -9, -9, 7, -3,
    -- layer=1 filter=4 channel=98
    -9, 3, 0, -12, 1, 8, 8, 3, -10,
    -- layer=1 filter=4 channel=99
    4, -9, -4, 8, -6, 0, -10, -2, 2,
    -- layer=1 filter=4 channel=100
    2, 5, 4, 6, -3, 6, -14, 0, 6,
    -- layer=1 filter=4 channel=101
    -6, -3, -9, -9, -1, 2, -8, 0, 7,
    -- layer=1 filter=4 channel=102
    -8, -11, -2, 8, 5, -1, 5, -3, -1,
    -- layer=1 filter=4 channel=103
    -14, 0, -1, -6, -13, -10, 3, -11, 7,
    -- layer=1 filter=4 channel=104
    -12, -1, -9, 5, -4, -5, -11, -8, 2,
    -- layer=1 filter=4 channel=105
    -8, 0, -3, 2, 4, -2, 3, -7, 1,
    -- layer=1 filter=4 channel=106
    -5, 4, -1, 3, -15, -1, -3, 0, -3,
    -- layer=1 filter=4 channel=107
    4, -1, 10, -9, -5, -1, -2, 5, -3,
    -- layer=1 filter=4 channel=108
    -2, -2, -9, 2, -12, -18, 9, -8, -16,
    -- layer=1 filter=4 channel=109
    -9, 9, -2, -11, -2, -4, -3, -7, -10,
    -- layer=1 filter=4 channel=110
    3, 0, -3, -4, -9, 8, -2, 3, -8,
    -- layer=1 filter=4 channel=111
    0, 1, 2, -11, 3, 3, 3, 0, -9,
    -- layer=1 filter=4 channel=112
    -7, -8, -9, 4, 7, 5, 1, -12, -7,
    -- layer=1 filter=4 channel=113
    -4, -3, -8, -4, -1, -7, -4, 11, 9,
    -- layer=1 filter=4 channel=114
    -14, -2, 2, 0, 2, -5, -3, -6, -6,
    -- layer=1 filter=4 channel=115
    1, -9, -9, -13, -6, 8, -12, -2, -3,
    -- layer=1 filter=4 channel=116
    -2, 9, -8, 0, 9, -9, -6, -6, 5,
    -- layer=1 filter=4 channel=117
    4, -8, -10, -4, -2, -9, -6, 2, 1,
    -- layer=1 filter=4 channel=118
    -5, -4, -9, -12, -3, -7, -16, -10, -8,
    -- layer=1 filter=4 channel=119
    -2, -16, -4, -11, -12, -6, -1, 1, 0,
    -- layer=1 filter=4 channel=120
    -2, -4, 2, 1, 6, -7, -7, 3, -11,
    -- layer=1 filter=4 channel=121
    -3, -5, -8, 4, 12, -12, 0, -6, 0,
    -- layer=1 filter=4 channel=122
    -5, 0, -1, 0, 4, -10, 8, -2, -10,
    -- layer=1 filter=4 channel=123
    0, 5, 0, -9, 0, -12, -8, 0, -11,
    -- layer=1 filter=4 channel=124
    8, 4, 6, 1, -2, 5, -8, -11, -10,
    -- layer=1 filter=4 channel=125
    0, -4, -3, -1, 13, -7, 0, -7, -4,
    -- layer=1 filter=4 channel=126
    -3, -9, -1, 2, -4, -3, 7, -5, -7,
    -- layer=1 filter=4 channel=127
    -3, 7, 0, 2, 2, -3, 0, -1, -2,
    -- layer=1 filter=5 channel=0
    -7, -9, -14, -5, 1, -11, -13, -5, -13,
    -- layer=1 filter=5 channel=1
    5, 1, -5, 0, -11, 1, 3, -13, 5,
    -- layer=1 filter=5 channel=2
    -11, -5, 0, 0, 0, -5, -7, -11, 1,
    -- layer=1 filter=5 channel=3
    5, 8, -4, -6, 4, -9, 0, 6, 7,
    -- layer=1 filter=5 channel=4
    -3, 6, -5, -5, 5, 0, -5, 0, 2,
    -- layer=1 filter=5 channel=5
    1, -11, -1, -3, -14, -19, 6, -8, 6,
    -- layer=1 filter=5 channel=6
    7, 0, -6, 2, -15, -13, -6, -9, 0,
    -- layer=1 filter=5 channel=7
    -15, -7, 3, -17, 7, 6, -12, 0, -5,
    -- layer=1 filter=5 channel=8
    -4, 0, -8, -1, -10, -8, -10, 0, -6,
    -- layer=1 filter=5 channel=9
    -15, -7, -12, 0, 10, 3, -1, 3, -5,
    -- layer=1 filter=5 channel=10
    -7, -4, 15, -11, 0, 0, -13, -15, 3,
    -- layer=1 filter=5 channel=11
    0, -13, -6, -10, -15, -14, -2, -12, 0,
    -- layer=1 filter=5 channel=12
    7, -6, 0, 6, -5, 0, -7, 4, 1,
    -- layer=1 filter=5 channel=13
    1, -8, -2, -12, -3, -4, 5, 0, -3,
    -- layer=1 filter=5 channel=14
    -3, 0, -5, -9, -13, 19, -17, 0, -4,
    -- layer=1 filter=5 channel=15
    8, 0, -13, -16, 9, -1, 2, -8, 0,
    -- layer=1 filter=5 channel=16
    -1, -15, 5, -15, -11, -4, 7, 4, -6,
    -- layer=1 filter=5 channel=17
    -7, -14, -8, 1, 0, -8, -1, -13, -7,
    -- layer=1 filter=5 channel=18
    -13, -1, -2, 9, 0, -8, -3, 0, 5,
    -- layer=1 filter=5 channel=19
    4, -3, -4, -11, 7, -8, -1, -5, 1,
    -- layer=1 filter=5 channel=20
    3, -6, -12, -2, -7, 1, -12, -4, -1,
    -- layer=1 filter=5 channel=21
    9, 1, 0, -2, -9, -7, 4, -13, 3,
    -- layer=1 filter=5 channel=22
    -3, -1, -9, -17, 0, -7, -10, -7, -13,
    -- layer=1 filter=5 channel=23
    -10, 5, -16, -11, -6, -2, -9, -4, -12,
    -- layer=1 filter=5 channel=24
    -9, -5, -4, -8, -9, -6, 2, -13, -11,
    -- layer=1 filter=5 channel=25
    -8, -6, 9, -11, 0, 2, -8, -10, -7,
    -- layer=1 filter=5 channel=26
    -4, -7, -1, -2, -4, -13, -13, -12, 4,
    -- layer=1 filter=5 channel=27
    4, -9, -9, -9, 3, -4, -15, 8, -9,
    -- layer=1 filter=5 channel=28
    -8, -15, -14, -12, -5, -9, -13, -10, -12,
    -- layer=1 filter=5 channel=29
    1, 1, 9, 0, 0, 11, -6, -9, -7,
    -- layer=1 filter=5 channel=30
    -8, 1, -7, 12, -4, -14, -11, -10, 12,
    -- layer=1 filter=5 channel=31
    6, 11, -4, -4, -11, -14, -16, -13, -2,
    -- layer=1 filter=5 channel=32
    -12, 1, 1, 1, -11, -15, -2, 6, -2,
    -- layer=1 filter=5 channel=33
    6, 8, 8, -14, -4, -17, -14, 1, -5,
    -- layer=1 filter=5 channel=34
    -11, 2, -8, -10, -3, 3, -3, 7, 3,
    -- layer=1 filter=5 channel=35
    0, -4, -12, -10, 0, -2, -12, -6, 4,
    -- layer=1 filter=5 channel=36
    0, 2, -12, -3, -12, -19, -14, -13, -12,
    -- layer=1 filter=5 channel=37
    -11, -2, 2, -9, -8, -21, 6, 2, 0,
    -- layer=1 filter=5 channel=38
    -11, 0, -13, -2, 3, -2, -9, -6, -9,
    -- layer=1 filter=5 channel=39
    -12, -4, -2, -7, 1, -14, -5, -4, -5,
    -- layer=1 filter=5 channel=40
    1, -8, 3, -5, -17, 0, -6, -15, -4,
    -- layer=1 filter=5 channel=41
    -6, 2, -8, -7, 3, -9, 1, -1, -2,
    -- layer=1 filter=5 channel=42
    -8, 7, 4, 2, 8, 6, 6, 3, 10,
    -- layer=1 filter=5 channel=43
    -16, -12, -10, -1, -10, -9, 4, -10, -1,
    -- layer=1 filter=5 channel=44
    0, -9, -17, -11, -7, -2, -6, -3, 4,
    -- layer=1 filter=5 channel=45
    -1, -11, 3, -5, -5, 2, -3, 1, 1,
    -- layer=1 filter=5 channel=46
    0, 11, 8, -6, -1, 3, 10, -8, 9,
    -- layer=1 filter=5 channel=47
    -9, -9, -8, 1, -10, -14, 0, -13, 6,
    -- layer=1 filter=5 channel=48
    -7, -9, -13, 0, -9, -15, 2, -8, -6,
    -- layer=1 filter=5 channel=49
    -9, -5, -4, -4, -3, -12, -5, -7, 0,
    -- layer=1 filter=5 channel=50
    1, -5, -1, -11, 0, 1, 6, -9, -3,
    -- layer=1 filter=5 channel=51
    -4, 3, 1, -2, -12, -11, 2, 0, -10,
    -- layer=1 filter=5 channel=52
    14, 1, -8, 0, 0, -14, 6, -3, -9,
    -- layer=1 filter=5 channel=53
    2, -2, 2, -5, -5, -9, -4, 6, -7,
    -- layer=1 filter=5 channel=54
    -9, -10, -1, -4, 4, -8, 3, -10, 1,
    -- layer=1 filter=5 channel=55
    -12, -10, -16, -7, -14, -19, 0, 5, -16,
    -- layer=1 filter=5 channel=56
    -6, 6, 0, 6, 4, -9, 6, -8, -3,
    -- layer=1 filter=5 channel=57
    0, -2, 5, -13, -11, 4, -4, -12, -2,
    -- layer=1 filter=5 channel=58
    -11, -12, 9, 1, -1, 2, -14, -7, 4,
    -- layer=1 filter=5 channel=59
    8, 5, 6, 0, -4, -5, 7, 0, 7,
    -- layer=1 filter=5 channel=60
    10, 1, -8, 6, 6, -7, 6, 1, -8,
    -- layer=1 filter=5 channel=61
    5, 11, 6, 8, 3, 6, 3, -1, -8,
    -- layer=1 filter=5 channel=62
    8, -14, 5, -2, -6, -14, 9, -8, -2,
    -- layer=1 filter=5 channel=63
    -7, -4, -4, 6, -13, -18, -11, -4, -4,
    -- layer=1 filter=5 channel=64
    4, -14, -5, -4, 0, -4, 1, -14, -6,
    -- layer=1 filter=5 channel=65
    2, -8, -11, -13, -6, 0, -16, -12, -5,
    -- layer=1 filter=5 channel=66
    -2, -15, -2, -7, -13, -15, -6, -10, -10,
    -- layer=1 filter=5 channel=67
    11, 1, 6, -4, 1, -1, -3, 8, -1,
    -- layer=1 filter=5 channel=68
    -2, 7, -18, -8, -14, -10, -11, 1, -5,
    -- layer=1 filter=5 channel=69
    0, 3, 2, -4, -9, -4, 6, 0, -10,
    -- layer=1 filter=5 channel=70
    1, 3, -17, -4, -7, 7, -16, -11, -2,
    -- layer=1 filter=5 channel=71
    -14, -12, -12, 3, -1, -8, -1, -3, -15,
    -- layer=1 filter=5 channel=72
    -10, -1, -10, -10, -10, -16, -3, -12, -7,
    -- layer=1 filter=5 channel=73
    -2, 8, 2, 5, 6, -6, -9, 6, -5,
    -- layer=1 filter=5 channel=74
    -2, -4, -8, -6, -12, -3, -13, -5, -2,
    -- layer=1 filter=5 channel=75
    4, -2, 4, -5, -5, 2, -6, -10, 8,
    -- layer=1 filter=5 channel=76
    1, 5, -16, 0, -1, -17, 2, -2, -8,
    -- layer=1 filter=5 channel=77
    -3, -3, -3, -4, -13, -2, 3, -6, -10,
    -- layer=1 filter=5 channel=78
    -16, -7, -16, -16, -3, -3, -3, -12, -16,
    -- layer=1 filter=5 channel=79
    -3, -4, -1, -11, -12, -4, 6, -1, -1,
    -- layer=1 filter=5 channel=80
    -7, 2, -11, -4, -13, 3, 8, 0, -4,
    -- layer=1 filter=5 channel=81
    0, -6, 3, 2, -5, -5, 0, -7, -17,
    -- layer=1 filter=5 channel=82
    -3, -2, 3, -7, -1, 1, -5, -5, -2,
    -- layer=1 filter=5 channel=83
    -9, -8, -9, -11, 3, -13, 3, 0, -10,
    -- layer=1 filter=5 channel=84
    -10, 8, -2, 7, 0, -6, -12, 1, 3,
    -- layer=1 filter=5 channel=85
    -8, -7, -4, 0, -6, 6, -2, 3, 5,
    -- layer=1 filter=5 channel=86
    0, -2, -7, -17, -7, -5, -4, -17, -20,
    -- layer=1 filter=5 channel=87
    -11, 6, -10, 2, 6, 6, 4, 2, -6,
    -- layer=1 filter=5 channel=88
    -6, 9, -5, -7, 7, -9, -1, 6, 0,
    -- layer=1 filter=5 channel=89
    1, 0, -15, -9, -11, 0, -9, -8, -6,
    -- layer=1 filter=5 channel=90
    4, 1, -9, -5, -13, -16, 1, 1, -9,
    -- layer=1 filter=5 channel=91
    -10, -11, -14, 4, -8, 3, 1, -5, -14,
    -- layer=1 filter=5 channel=92
    -3, 5, 5, 0, -6, -2, 5, 0, -6,
    -- layer=1 filter=5 channel=93
    -2, -3, 0, -16, -9, -10, -12, -10, -9,
    -- layer=1 filter=5 channel=94
    -3, -5, -16, -16, -13, 2, -9, -8, -11,
    -- layer=1 filter=5 channel=95
    6, 5, -5, -2, 0, -16, 2, 0, 3,
    -- layer=1 filter=5 channel=96
    9, -4, -10, -12, -5, -4, 0, -5, 1,
    -- layer=1 filter=5 channel=97
    -2, -2, 2, -14, 3, -12, -10, -9, -6,
    -- layer=1 filter=5 channel=98
    -9, -11, 19, 0, -9, -8, -3, 0, -17,
    -- layer=1 filter=5 channel=99
    0, 2, -4, -6, -13, -4, -7, 1, -12,
    -- layer=1 filter=5 channel=100
    -3, -7, -7, -13, -1, -4, -17, -15, -8,
    -- layer=1 filter=5 channel=101
    1, 0, -6, -10, -14, 0, -13, -9, -3,
    -- layer=1 filter=5 channel=102
    0, -2, -7, -11, -2, -9, -7, 2, -10,
    -- layer=1 filter=5 channel=103
    -5, 3, 1, 2, -13, -13, -15, -11, 0,
    -- layer=1 filter=5 channel=104
    -4, -7, -11, -2, -8, -16, -7, -10, -9,
    -- layer=1 filter=5 channel=105
    -12, 1, 2, -5, -13, -7, -13, -5, 0,
    -- layer=1 filter=5 channel=106
    3, 1, -3, -1, -9, -7, 0, -13, -3,
    -- layer=1 filter=5 channel=107
    0, -4, 0, 6, -5, -7, -10, -3, -6,
    -- layer=1 filter=5 channel=108
    -1, 13, -3, 10, 6, 0, 0, 7, 9,
    -- layer=1 filter=5 channel=109
    -10, -4, 0, -11, -6, -8, 9, -7, 9,
    -- layer=1 filter=5 channel=110
    -4, -9, 0, -12, -1, -14, -16, -15, -7,
    -- layer=1 filter=5 channel=111
    0, -7, 4, 7, -16, -7, -3, -5, 4,
    -- layer=1 filter=5 channel=112
    5, 0, 0, -8, -14, -4, -10, -9, 5,
    -- layer=1 filter=5 channel=113
    -18, -5, -5, -14, 6, -3, -1, -9, 0,
    -- layer=1 filter=5 channel=114
    6, -19, -9, -11, -16, -19, 6, -6, -8,
    -- layer=1 filter=5 channel=115
    -9, -4, -15, -10, -17, 1, 2, -7, -1,
    -- layer=1 filter=5 channel=116
    0, 2, 2, -8, -2, 1, 4, 10, -8,
    -- layer=1 filter=5 channel=117
    -6, -4, -2, 0, -9, 4, -4, 7, -2,
    -- layer=1 filter=5 channel=118
    3, -3, -7, 0, 0, -1, -5, 0, 3,
    -- layer=1 filter=5 channel=119
    -8, 5, -7, 0, 8, -11, -12, -6, 9,
    -- layer=1 filter=5 channel=120
    -10, -9, -7, -7, -2, -9, 4, -6, -8,
    -- layer=1 filter=5 channel=121
    1, -2, -10, -8, -1, 8, 2, -1, -8,
    -- layer=1 filter=5 channel=122
    0, 7, -6, -5, -1, 0, 0, 10, -8,
    -- layer=1 filter=5 channel=123
    0, -1, -1, -12, -3, -6, -13, -6, -16,
    -- layer=1 filter=5 channel=124
    4, -7, -7, -1, -1, -7, 4, 2, 3,
    -- layer=1 filter=5 channel=125
    1, -5, 0, -17, -5, -4, -21, -16, 6,
    -- layer=1 filter=5 channel=126
    0, -8, 3, -3, -7, -18, -9, -6, -15,
    -- layer=1 filter=5 channel=127
    10, -6, -2, -2, -12, 0, 8, 0, 9,
    -- layer=1 filter=6 channel=0
    -25, -8, -6, -25, -10, -9, -15, -27, -14,
    -- layer=1 filter=6 channel=1
    -24, -9, 6, -10, -20, -12, 0, -17, 3,
    -- layer=1 filter=6 channel=2
    -2, 0, 6, 2, 6, 0, 43, -12, -24,
    -- layer=1 filter=6 channel=3
    -1, 15, 1, 9, -8, 2, 0, 8, -1,
    -- layer=1 filter=6 channel=4
    -11, -5, 0, 1, 2, -8, -8, -14, -6,
    -- layer=1 filter=6 channel=5
    -8, -2, 13, 9, -4, -10, 9, 9, 53,
    -- layer=1 filter=6 channel=6
    -11, -14, -58, 3, -1, 1, -35, -1, -24,
    -- layer=1 filter=6 channel=7
    20, -18, 11, 19, 24, 12, 22, 54, 29,
    -- layer=1 filter=6 channel=8
    -4, 13, 1, 16, 17, 6, 7, -15, 13,
    -- layer=1 filter=6 channel=9
    18, 4, 28, -7, -17, 11, -38, -25, -43,
    -- layer=1 filter=6 channel=10
    9, -3, 8, 9, 15, 6, 13, 52, 25,
    -- layer=1 filter=6 channel=11
    0, -25, -18, -1, 5, -16, 15, 23, 17,
    -- layer=1 filter=6 channel=12
    -20, 21, -19, 10, 11, 11, -58, -29, -58,
    -- layer=1 filter=6 channel=13
    4, 20, 37, -2, 19, 17, -22, 3, -17,
    -- layer=1 filter=6 channel=14
    -10, -29, -10, -12, -5, -11, -7, -5, -21,
    -- layer=1 filter=6 channel=15
    -22, 23, 30, -37, -38, -30, 17, 13, 16,
    -- layer=1 filter=6 channel=16
    -21, -5, 12, 28, 0, 4, 0, -3, 20,
    -- layer=1 filter=6 channel=17
    8, 19, 33, -10, 2, 15, -8, -7, 1,
    -- layer=1 filter=6 channel=18
    22, 23, -13, 16, 31, 10, 13, 19, -5,
    -- layer=1 filter=6 channel=19
    -7, -3, -3, 39, -13, -38, -21, 5, 26,
    -- layer=1 filter=6 channel=20
    32, 40, 29, 18, 27, 35, 2, 11, 8,
    -- layer=1 filter=6 channel=21
    -36, -12, -8, -24, -12, -25, -12, -38, -13,
    -- layer=1 filter=6 channel=22
    36, 53, 35, 19, 32, 15, 10, 5, 0,
    -- layer=1 filter=6 channel=23
    -63, -58, -44, -77, -98, -44, -15, -43, -21,
    -- layer=1 filter=6 channel=24
    -36, -1, 15, -49, -31, -33, -18, -14, -28,
    -- layer=1 filter=6 channel=25
    0, -24, 20, 10, -10, -13, -1, 21, 28,
    -- layer=1 filter=6 channel=26
    17, 28, 53, -21, -13, 11, 18, 16, 8,
    -- layer=1 filter=6 channel=27
    -10, -23, 24, 17, -32, 5, 75, 54, 27,
    -- layer=1 filter=6 channel=28
    -17, -1, 12, 1, 12, -6, -19, 16, 6,
    -- layer=1 filter=6 channel=29
    11, 3, -18, 31, 11, 10, 29, 1, -20,
    -- layer=1 filter=6 channel=30
    13, 8, 13, 39, 18, 23, 10, 22, -12,
    -- layer=1 filter=6 channel=31
    6, 9, -45, 34, 36, 15, -8, 6, -11,
    -- layer=1 filter=6 channel=32
    -25, 16, 9, 6, -20, 0, 26, 2, 12,
    -- layer=1 filter=6 channel=33
    -2, -21, -10, -6, -12, -17, -15, -16, -32,
    -- layer=1 filter=6 channel=34
    -58, -36, -37, -52, -42, -33, -26, -24, -24,
    -- layer=1 filter=6 channel=35
    -27, -16, 2, -5, -10, -4, -4, -2, -9,
    -- layer=1 filter=6 channel=36
    -20, -42, -13, -30, -17, -18, 1, 7, 10,
    -- layer=1 filter=6 channel=37
    -18, -10, 1, 14, -7, -15, 6, 36, 58,
    -- layer=1 filter=6 channel=38
    19, 26, -2, 18, 39, 17, -2, 8, 0,
    -- layer=1 filter=6 channel=39
    -11, -28, -10, -14, -19, -33, -28, -13, -6,
    -- layer=1 filter=6 channel=40
    69, 30, -17, 42, 68, 44, 47, 60, 7,
    -- layer=1 filter=6 channel=41
    0, -43, 19, -5, -73, -24, -4, -10, -77,
    -- layer=1 filter=6 channel=42
    8, -6, 8, 30, 10, 16, 14, 0, -32,
    -- layer=1 filter=6 channel=43
    -39, -19, -10, -4, -43, -30, 0, -24, 8,
    -- layer=1 filter=6 channel=44
    5, 20, 36, -34, -4, 1, 45, -4, 25,
    -- layer=1 filter=6 channel=45
    -22, 13, 14, -15, -14, -11, -6, -16, -1,
    -- layer=1 filter=6 channel=46
    -8, -19, 24, 72, -1, -29, 27, 24, 51,
    -- layer=1 filter=6 channel=47
    -60, -45, -12, -20, -63, -26, 6, 17, -3,
    -- layer=1 filter=6 channel=48
    13, 0, 5, -19, -14, -3, -23, -1, -11,
    -- layer=1 filter=6 channel=49
    -23, -24, -18, -10, -23, -21, -4, -15, -15,
    -- layer=1 filter=6 channel=50
    4, 0, -18, -5, -3, 24, 8, -1, -4,
    -- layer=1 filter=6 channel=51
    9, -10, -20, -16, 12, -16, -10, 9, -1,
    -- layer=1 filter=6 channel=52
    2, -3, -4, -17, -11, 1, -11, -17, -9,
    -- layer=1 filter=6 channel=53
    10, 12, -5, 10, 6, 0, 17, 1, 11,
    -- layer=1 filter=6 channel=54
    0, -53, -16, 9, -22, -38, -6, 30, 23,
    -- layer=1 filter=6 channel=55
    -38, -65, -34, -29, -35, -25, 21, 3, 1,
    -- layer=1 filter=6 channel=56
    -2, -8, 0, -2, 0, 9, 11, -6, 11,
    -- layer=1 filter=6 channel=57
    54, 13, 6, 39, 56, 16, 40, 74, 37,
    -- layer=1 filter=6 channel=58
    -35, -90, -45, -29, -71, -61, 20, 22, 4,
    -- layer=1 filter=6 channel=59
    -11, -19, -5, -2, 1, 13, -13, 2, -1,
    -- layer=1 filter=6 channel=60
    12, -2, 20, 8, 11, 13, 16, 6, 14,
    -- layer=1 filter=6 channel=61
    1, -10, 13, 7, -16, 1, 7, 0, 1,
    -- layer=1 filter=6 channel=62
    -4, 12, 8, 4, 2, 1, -16, -11, 17,
    -- layer=1 filter=6 channel=63
    -22, -29, -22, -29, -32, -28, -20, -14, -19,
    -- layer=1 filter=6 channel=64
    -5, 0, -4, -6, 10, -11, -12, -18, -10,
    -- layer=1 filter=6 channel=65
    -15, -8, -3, -7, -16, -5, -36, -32, -14,
    -- layer=1 filter=6 channel=66
    -14, -22, -26, -25, -24, -16, 6, 4, 0,
    -- layer=1 filter=6 channel=67
    -61, -54, -50, -45, -41, -59, -70, -63, -50,
    -- layer=1 filter=6 channel=68
    -4, 5, 20, -41, -31, -28, 27, 8, 17,
    -- layer=1 filter=6 channel=69
    -2, 30, 15, -21, 12, 1, 11, -2, 27,
    -- layer=1 filter=6 channel=70
    -40, -58, -52, -18, -30, -38, -62, -14, -24,
    -- layer=1 filter=6 channel=71
    -46, -41, -14, -19, -44, -25, -40, -36, -2,
    -- layer=1 filter=6 channel=72
    10, 16, 20, 40, 7, -5, 9, -11, -17,
    -- layer=1 filter=6 channel=73
    -5, -1, -4, -14, -12, -13, -7, -13, -7,
    -- layer=1 filter=6 channel=74
    -2, 0, -17, -4, 3, -18, -6, 17, 19,
    -- layer=1 filter=6 channel=75
    -4, 20, -28, 9, -12, -9, -47, -23, -58,
    -- layer=1 filter=6 channel=76
    21, -19, 10, 3, -32, -1, -11, -37, -15,
    -- layer=1 filter=6 channel=77
    -36, -16, -17, -41, -34, -27, -29, -37, -11,
    -- layer=1 filter=6 channel=78
    -1, 0, -15, -30, 9, 6, -21, -5, 25,
    -- layer=1 filter=6 channel=79
    -12, 26, 2, 19, 21, 21, -10, -13, 0,
    -- layer=1 filter=6 channel=80
    -7, -19, -8, 3, 2, 1, -12, -8, -1,
    -- layer=1 filter=6 channel=81
    -26, -19, -3, -66, -73, -5, -41, -49, -27,
    -- layer=1 filter=6 channel=82
    -11, -2, -11, -25, -5, -5, -11, -14, -7,
    -- layer=1 filter=6 channel=83
    -20, 1, 6, -20, -19, 9, 7, -5, 1,
    -- layer=1 filter=6 channel=84
    36, 12, 1, 0, -10, -3, 0, 25, -19,
    -- layer=1 filter=6 channel=85
    -16, -44, -37, -41, -68, -44, 3, 9, -3,
    -- layer=1 filter=6 channel=86
    9, 4, 0, 40, 15, 18, 12, 24, 29,
    -- layer=1 filter=6 channel=87
    12, 15, 7, 40, 9, -25, 15, -27, -25,
    -- layer=1 filter=6 channel=88
    -11, 0, 3, -1, -10, -1, -8, -2, -2,
    -- layer=1 filter=6 channel=89
    -24, 3, -10, -27, -36, -22, -10, -20, -18,
    -- layer=1 filter=6 channel=90
    -10, 21, 51, -44, -34, 0, 11, -22, 13,
    -- layer=1 filter=6 channel=91
    32, 20, 8, 22, 40, 25, 12, 24, 15,
    -- layer=1 filter=6 channel=92
    16, -25, 34, -48, -52, -26, -10, 16, -18,
    -- layer=1 filter=6 channel=93
    -8, -12, -11, -23, -23, -5, -29, -28, -23,
    -- layer=1 filter=6 channel=94
    -10, 14, 4, -3, 17, -2, -15, -2, -3,
    -- layer=1 filter=6 channel=95
    19, 5, -20, 21, 1, 0, 0, -11, -11,
    -- layer=1 filter=6 channel=96
    -22, -18, -5, -19, -13, -23, -7, 0, -13,
    -- layer=1 filter=6 channel=97
    3, 8, 7, -24, -11, 1, -17, -17, -7,
    -- layer=1 filter=6 channel=98
    -9, 25, 2, 19, 17, 23, 0, -19, -9,
    -- layer=1 filter=6 channel=99
    -5, -23, -26, -51, -23, -38, 18, 6, 10,
    -- layer=1 filter=6 channel=100
    -38, -30, -28, -35, -14, -26, -1, -3, 14,
    -- layer=1 filter=6 channel=101
    27, 21, 10, 17, 33, 16, 2, 0, 1,
    -- layer=1 filter=6 channel=102
    3, 4, -12, -6, 11, 16, -29, -8, 0,
    -- layer=1 filter=6 channel=103
    -26, -40, -13, -15, -9, 8, 25, 19, 9,
    -- layer=1 filter=6 channel=104
    -4, -12, 6, 11, -20, 7, 4, -15, 2,
    -- layer=1 filter=6 channel=105
    6, -8, 4, -26, -6, -10, -19, -17, -1,
    -- layer=1 filter=6 channel=106
    11, 9, 17, 11, 12, 1, 5, 3, -11,
    -- layer=1 filter=6 channel=107
    -16, -16, -16, -4, -11, -12, -9, -8, -8,
    -- layer=1 filter=6 channel=108
    3, -14, 30, -23, -56, -24, 23, 2, -12,
    -- layer=1 filter=6 channel=109
    8, 3, -4, 0, -8, -5, 8, 2, 5,
    -- layer=1 filter=6 channel=110
    10, 0, 4, 5, 3, 0, -17, -1, -8,
    -- layer=1 filter=6 channel=111
    46, 10, 25, 1, 16, 0, 5, 11, -11,
    -- layer=1 filter=6 channel=112
    -3, 7, -29, 5, -30, -18, -16, -29, -32,
    -- layer=1 filter=6 channel=113
    -30, -54, -29, -8, -33, -56, -42, -12, -49,
    -- layer=1 filter=6 channel=114
    -17, -23, -6, 0, -45, -33, 2, -15, 35,
    -- layer=1 filter=6 channel=115
    36, 15, 1, 42, 27, 8, 4, 27, 17,
    -- layer=1 filter=6 channel=116
    -8, 6, 0, 0, 5, 7, 0, 7, 6,
    -- layer=1 filter=6 channel=117
    36, 0, -2, -1, -5, -6, -5, -27, -29,
    -- layer=1 filter=6 channel=118
    22, 6, 7, 18, 6, 12, 22, 8, 17,
    -- layer=1 filter=6 channel=119
    -8, -10, 30, -39, -41, -11, 7, -2, -24,
    -- layer=1 filter=6 channel=120
    -5, -7, -6, -4, 6, 6, -28, -7, 16,
    -- layer=1 filter=6 channel=121
    0, -8, 26, 40, 15, -8, -15, -17, -24,
    -- layer=1 filter=6 channel=122
    10, -10, -10, 5, 0, 4, 0, -3, -5,
    -- layer=1 filter=6 channel=123
    -32, -43, -36, 1, -44, -38, 14, -5, -25,
    -- layer=1 filter=6 channel=124
    -1, 4, 16, -6, 0, 1, -1, 9, 0,
    -- layer=1 filter=6 channel=125
    -5, -42, -40, -29, -30, -56, -37, -1, -25,
    -- layer=1 filter=6 channel=126
    -33, -4, -3, -59, 3, 2, 16, -17, -32,
    -- layer=1 filter=6 channel=127
    36, 17, 17, 45, 35, 25, 32, 17, 18,
    -- layer=1 filter=7 channel=0
    -4, -3, 3, -8, 6, 6, 0, -9, -4,
    -- layer=1 filter=7 channel=1
    -7, -7, -6, 0, 4, -4, -4, -6, -7,
    -- layer=1 filter=7 channel=2
    -1, 0, -2, -15, 3, -15, -9, 0, -3,
    -- layer=1 filter=7 channel=3
    6, -10, -10, -6, -8, 2, -8, 2, 2,
    -- layer=1 filter=7 channel=4
    -1, 2, 6, 0, 6, 0, 5, 0, 0,
    -- layer=1 filter=7 channel=5
    -2, -7, 3, -4, -2, 2, -14, -4, -10,
    -- layer=1 filter=7 channel=6
    -10, 4, 5, -4, -5, -2, -6, 6, 3,
    -- layer=1 filter=7 channel=7
    0, -10, -3, -5, -8, -1, 0, -6, -9,
    -- layer=1 filter=7 channel=8
    5, -7, 0, -7, -12, 5, -1, -7, 7,
    -- layer=1 filter=7 channel=9
    8, 8, 4, -14, -1, -8, -10, -10, -7,
    -- layer=1 filter=7 channel=10
    -15, 0, 2, -6, -2, 7, -1, -14, -2,
    -- layer=1 filter=7 channel=11
    -4, -4, 4, 3, -1, 0, 1, -1, -11,
    -- layer=1 filter=7 channel=12
    -5, 9, -2, -6, -2, -9, -12, -15, -12,
    -- layer=1 filter=7 channel=13
    -12, -13, -3, -3, 2, -8, -12, -1, 0,
    -- layer=1 filter=7 channel=14
    1, -10, -12, -7, -12, -10, -9, 4, -5,
    -- layer=1 filter=7 channel=15
    -10, -6, -11, -1, -6, 0, 0, -5, -15,
    -- layer=1 filter=7 channel=16
    -3, 8, -8, -3, 1, 3, -12, 4, 3,
    -- layer=1 filter=7 channel=17
    -2, 2, -9, 0, 2, -3, 5, 0, -5,
    -- layer=1 filter=7 channel=18
    -5, -6, -10, -12, 4, -5, 6, -10, -4,
    -- layer=1 filter=7 channel=19
    5, -6, 4, -1, 6, -3, 0, -6, 1,
    -- layer=1 filter=7 channel=20
    7, -7, -7, 2, -10, -11, -2, -11, -10,
    -- layer=1 filter=7 channel=21
    1, -11, -4, -6, 6, -7, 6, -5, -8,
    -- layer=1 filter=7 channel=22
    -1, 5, -1, 1, -8, 4, -12, 0, -5,
    -- layer=1 filter=7 channel=23
    5, -4, -12, 6, 6, 0, 1, -12, 7,
    -- layer=1 filter=7 channel=24
    -7, -7, -6, 0, -6, -9, -16, -10, 1,
    -- layer=1 filter=7 channel=25
    -4, 1, -5, 3, 2, 0, -7, -6, -15,
    -- layer=1 filter=7 channel=26
    -2, -5, 1, -13, -3, -15, -9, -10, -13,
    -- layer=1 filter=7 channel=27
    1, -7, 3, -14, -14, -4, 0, -2, -3,
    -- layer=1 filter=7 channel=28
    3, 0, 2, 4, -7, -10, -12, -11, -5,
    -- layer=1 filter=7 channel=29
    4, 10, -7, 4, 3, -9, -3, -2, -6,
    -- layer=1 filter=7 channel=30
    -6, -11, -4, 4, -18, -10, -9, -9, 4,
    -- layer=1 filter=7 channel=31
    3, -7, -8, 1, -13, -4, -3, -2, -17,
    -- layer=1 filter=7 channel=32
    -7, -2, -1, -1, 0, -4, 6, 2, -7,
    -- layer=1 filter=7 channel=33
    -3, -6, -5, 9, 3, -2, 5, -2, -2,
    -- layer=1 filter=7 channel=34
    -6, 7, 8, 1, 2, -5, -13, -7, -2,
    -- layer=1 filter=7 channel=35
    -11, -6, 5, 1, 1, -9, -6, -8, 6,
    -- layer=1 filter=7 channel=36
    -6, -5, 2, -3, 8, -11, -9, 1, -7,
    -- layer=1 filter=7 channel=37
    -12, 4, 2, 4, 6, 1, -4, 1, -4,
    -- layer=1 filter=7 channel=38
    0, -8, 4, 0, 2, 6, -9, 3, 0,
    -- layer=1 filter=7 channel=39
    -3, -11, 4, 1, -1, -10, 0, -7, 2,
    -- layer=1 filter=7 channel=40
    0, 6, 2, 3, -1, -13, 0, 2, -7,
    -- layer=1 filter=7 channel=41
    -7, -2, -10, -9, 5, -8, -7, -5, 0,
    -- layer=1 filter=7 channel=42
    -15, -9, -2, -1, 0, -14, -11, 3, -6,
    -- layer=1 filter=7 channel=43
    5, 2, 6, 2, -10, 1, 2, 6, 0,
    -- layer=1 filter=7 channel=44
    -6, -5, 4, -5, -13, -8, -9, -1, -9,
    -- layer=1 filter=7 channel=45
    -6, 5, 8, -1, -11, -3, -7, -9, -11,
    -- layer=1 filter=7 channel=46
    -12, -3, -3, -2, -4, -9, 0, -6, 3,
    -- layer=1 filter=7 channel=47
    -12, -12, -5, 2, -12, -7, 0, -9, -12,
    -- layer=1 filter=7 channel=48
    0, 6, 8, 3, -3, 7, -13, 5, -6,
    -- layer=1 filter=7 channel=49
    -4, 2, 7, -2, 0, 7, 6, 0, -1,
    -- layer=1 filter=7 channel=50
    5, 5, -6, 7, -12, 3, -7, -1, -8,
    -- layer=1 filter=7 channel=51
    0, -4, 0, 7, 6, -4, 3, -6, 5,
    -- layer=1 filter=7 channel=52
    2, 3, -8, 2, 7, -7, 2, -10, 1,
    -- layer=1 filter=7 channel=53
    7, 8, -7, -11, -6, -10, -3, -5, -9,
    -- layer=1 filter=7 channel=54
    4, 2, -12, 1, -15, 1, -3, -11, 1,
    -- layer=1 filter=7 channel=55
    0, 3, 2, -8, 0, -16, -15, -4, 2,
    -- layer=1 filter=7 channel=56
    5, -10, -7, 8, -7, 1, -7, 8, 4,
    -- layer=1 filter=7 channel=57
    -6, -11, 4, 1, -5, -7, -8, -10, 4,
    -- layer=1 filter=7 channel=58
    -9, 1, -6, -8, 5, -7, -9, 6, -2,
    -- layer=1 filter=7 channel=59
    2, -11, -10, -3, -8, 5, -7, -3, -11,
    -- layer=1 filter=7 channel=60
    1, 5, 0, 0, 6, 1, 5, 10, 4,
    -- layer=1 filter=7 channel=61
    1, -2, 9, -6, -2, -5, -5, -8, 8,
    -- layer=1 filter=7 channel=62
    -14, 1, 7, -2, 2, -2, -5, 8, 4,
    -- layer=1 filter=7 channel=63
    0, -6, -7, -3, -5, -2, -2, 7, -12,
    -- layer=1 filter=7 channel=64
    -9, -11, -12, -8, -12, -10, 5, -5, 0,
    -- layer=1 filter=7 channel=65
    7, 1, 8, -11, 7, 6, 1, 3, 0,
    -- layer=1 filter=7 channel=66
    -8, -10, -2, -1, 7, -7, 7, -10, 6,
    -- layer=1 filter=7 channel=67
    2, 8, -10, 6, 10, 5, 6, 6, 8,
    -- layer=1 filter=7 channel=68
    4, -14, 4, 5, 0, -12, -1, -10, 7,
    -- layer=1 filter=7 channel=69
    -5, -9, -10, -3, 6, 6, -11, -2, -2,
    -- layer=1 filter=7 channel=70
    3, -4, -2, -5, -5, -8, -3, 4, -6,
    -- layer=1 filter=7 channel=71
    4, 0, -3, -6, -6, 3, -6, -10, 0,
    -- layer=1 filter=7 channel=72
    8, 4, 4, -9, 4, -9, 2, 6, 3,
    -- layer=1 filter=7 channel=73
    -7, -9, -8, -2, -8, -11, -7, -4, 6,
    -- layer=1 filter=7 channel=74
    -9, 6, -6, 4, -9, -11, 7, 1, -9,
    -- layer=1 filter=7 channel=75
    -4, -14, -9, -3, -10, -8, 2, 3, -13,
    -- layer=1 filter=7 channel=76
    -3, 5, -11, -7, -7, -5, 3, -4, 0,
    -- layer=1 filter=7 channel=77
    -6, -10, 1, -6, -3, -7, -4, 3, 6,
    -- layer=1 filter=7 channel=78
    -7, 7, -5, 6, 2, 7, 3, -1, -1,
    -- layer=1 filter=7 channel=79
    -12, -7, -7, -3, 7, -10, 4, 2, -8,
    -- layer=1 filter=7 channel=80
    -5, 1, 0, 5, 7, 0, -1, -10, -9,
    -- layer=1 filter=7 channel=81
    0, -10, 2, 2, 7, -4, -7, 7, 4,
    -- layer=1 filter=7 channel=82
    2, -9, 6, -7, 6, -4, 0, 2, -3,
    -- layer=1 filter=7 channel=83
    -6, 7, 3, 8, -9, -7, -7, 5, -12,
    -- layer=1 filter=7 channel=84
    -3, 4, 0, 2, -18, 2, -1, -6, -8,
    -- layer=1 filter=7 channel=85
    0, -12, -8, -5, 4, -11, -4, -3, -11,
    -- layer=1 filter=7 channel=86
    0, -8, 0, 0, -3, 5, 4, -1, 0,
    -- layer=1 filter=7 channel=87
    5, -9, 5, -1, 1, -11, -12, 4, -10,
    -- layer=1 filter=7 channel=88
    -6, 2, -3, 10, -5, 11, 4, -2, -1,
    -- layer=1 filter=7 channel=89
    -7, -8, -11, -5, 1, -8, -1, -7, 1,
    -- layer=1 filter=7 channel=90
    5, 4, 7, -10, 1, -4, 0, -6, -10,
    -- layer=1 filter=7 channel=91
    0, 4, -4, -3, -4, 3, 3, -10, -7,
    -- layer=1 filter=7 channel=92
    -11, -8, 7, 0, 0, 0, 4, -13, 6,
    -- layer=1 filter=7 channel=93
    4, 5, -10, -5, -4, -5, -1, 0, 6,
    -- layer=1 filter=7 channel=94
    -9, -5, 4, 3, -8, 1, -13, -3, -4,
    -- layer=1 filter=7 channel=95
    7, 5, -6, -2, 0, -12, 2, -6, 4,
    -- layer=1 filter=7 channel=96
    -5, -4, 1, -8, -2, 0, -2, 2, -4,
    -- layer=1 filter=7 channel=97
    0, -9, -3, 3, -2, 5, -10, -11, 5,
    -- layer=1 filter=7 channel=98
    -5, -5, 1, 5, 4, -10, -9, 4, -14,
    -- layer=1 filter=7 channel=99
    9, -8, -6, 6, 5, -2, -1, 1, -6,
    -- layer=1 filter=7 channel=100
    -1, -2, -10, -4, -5, 8, 4, 5, -2,
    -- layer=1 filter=7 channel=101
    8, 2, 9, 0, -9, -3, -12, 0, 1,
    -- layer=1 filter=7 channel=102
    -8, 3, 6, 0, -8, 6, -2, 1, 4,
    -- layer=1 filter=7 channel=103
    5, -8, -11, 5, -6, 6, -9, 8, 3,
    -- layer=1 filter=7 channel=104
    4, -1, -6, -2, -5, 4, -12, 0, 7,
    -- layer=1 filter=7 channel=105
    -1, 0, -2, -1, 7, 0, -7, -9, -6,
    -- layer=1 filter=7 channel=106
    -9, -10, -10, 5, -12, -3, -3, -7, -3,
    -- layer=1 filter=7 channel=107
    -3, -1, -4, -6, 5, -4, 9, -6, -10,
    -- layer=1 filter=7 channel=108
    0, -19, -11, -8, -13, -2, -13, 3, 7,
    -- layer=1 filter=7 channel=109
    -8, 10, 9, 3, -2, -4, 11, 5, -1,
    -- layer=1 filter=7 channel=110
    0, 4, 1, -2, -5, 4, -6, -7, 7,
    -- layer=1 filter=7 channel=111
    -10, -3, -11, -16, 1, 4, -6, 8, -4,
    -- layer=1 filter=7 channel=112
    -7, 6, 1, -7, -9, -5, 1, 3, -8,
    -- layer=1 filter=7 channel=113
    -11, 0, -10, 2, -8, 3, 5, -12, 3,
    -- layer=1 filter=7 channel=114
    -4, 1, 0, 3, -7, 0, -5, -10, -10,
    -- layer=1 filter=7 channel=115
    -7, -7, 2, -7, -8, 5, 7, -5, 0,
    -- layer=1 filter=7 channel=116
    -1, 6, 0, 5, 5, 8, -9, 0, -3,
    -- layer=1 filter=7 channel=117
    3, -9, -8, 7, -7, -1, 1, 4, 0,
    -- layer=1 filter=7 channel=118
    7, -2, -11, 0, 3, 6, -8, 1, -8,
    -- layer=1 filter=7 channel=119
    3, -9, -2, -3, 0, -9, -7, -7, -5,
    -- layer=1 filter=7 channel=120
    -7, -3, -11, -5, -6, -7, 4, -8, 8,
    -- layer=1 filter=7 channel=121
    -2, -10, -8, -11, -14, -14, -2, -16, -13,
    -- layer=1 filter=7 channel=122
    9, -8, 8, -6, 3, -3, -1, -9, 1,
    -- layer=1 filter=7 channel=123
    -9, -2, -6, 4, -5, 3, -13, -3, -13,
    -- layer=1 filter=7 channel=124
    -9, 0, 5, 7, 9, 3, -7, 7, 6,
    -- layer=1 filter=7 channel=125
    -2, 0, 9, -8, -8, -9, -4, 0, 6,
    -- layer=1 filter=7 channel=126
    3, 3, -4, 8, -6, -9, -5, 7, 0,
    -- layer=1 filter=7 channel=127
    -3, 8, -3, 3, -18, -12, 1, -10, -7,
    -- layer=1 filter=8 channel=0
    5, 7, 10, 10, 4, -3, 3, 7, -7,
    -- layer=1 filter=8 channel=1
    -12, 2, -19, -18, -26, -7, -6, -41, -40,
    -- layer=1 filter=8 channel=2
    63, 14, 1, 43, 13, -14, 47, 20, -6,
    -- layer=1 filter=8 channel=3
    1, 5, -3, -2, -6, -2, -13, 0, 2,
    -- layer=1 filter=8 channel=4
    4, -5, 5, -8, -6, -6, 6, 3, -10,
    -- layer=1 filter=8 channel=5
    -21, 3, -34, -51, -73, -38, -41, -85, -106,
    -- layer=1 filter=8 channel=6
    -12, 4, 4, 7, -12, 0, -18, -22, -21,
    -- layer=1 filter=8 channel=7
    36, 57, 43, 22, 47, 8, 28, 62, 5,
    -- layer=1 filter=8 channel=8
    -16, -22, -32, -45, -61, -37, -23, -78, -93,
    -- layer=1 filter=8 channel=9
    -37, -57, -3, -22, -17, -59, -14, -27, -21,
    -- layer=1 filter=8 channel=10
    32, 46, 36, 6, 36, 12, 16, 41, 17,
    -- layer=1 filter=8 channel=11
    0, 6, 2, 2, -10, -11, 3, 9, 3,
    -- layer=1 filter=8 channel=12
    -28, -77, -61, -11, -104, -80, -18, -63, 13,
    -- layer=1 filter=8 channel=13
    5, 5, 1, -2, 1, 0, -9, -17, 1,
    -- layer=1 filter=8 channel=14
    -1, 31, 26, -8, -13, -40, -19, 3, -19,
    -- layer=1 filter=8 channel=15
    14, 31, -25, -7, -36, -8, 34, -15, -42,
    -- layer=1 filter=8 channel=16
    -40, -35, -37, -51, -57, -22, -27, -77, -51,
    -- layer=1 filter=8 channel=17
    9, -2, -5, -5, 12, -15, 0, -1, -11,
    -- layer=1 filter=8 channel=18
    -6, -16, -3, -28, -29, -24, -16, -31, -6,
    -- layer=1 filter=8 channel=19
    -65, -55, -17, -15, -48, -32, -26, -58, 9,
    -- layer=1 filter=8 channel=20
    6, 2, 9, -7, -5, 0, -11, -8, -2,
    -- layer=1 filter=8 channel=21
    -9, -17, 2, -11, -9, 5, -8, -2, -4,
    -- layer=1 filter=8 channel=22
    1, 0, -10, -10, -20, -6, 16, -9, -13,
    -- layer=1 filter=8 channel=23
    0, 25, 10, 65, 28, 36, 59, 59, 42,
    -- layer=1 filter=8 channel=24
    -9, -19, 6, -32, 15, -13, -7, -10, -4,
    -- layer=1 filter=8 channel=25
    11, 20, 16, -13, 12, -15, -11, 27, -4,
    -- layer=1 filter=8 channel=26
    7, 38, -4, -1, 23, -9, 8, 17, 7,
    -- layer=1 filter=8 channel=27
    -19, -17, 11, -34, -24, 14, -53, -29, -26,
    -- layer=1 filter=8 channel=28
    -6, 9, 28, 1, 8, 7, -14, 13, 2,
    -- layer=1 filter=8 channel=29
    -3, -8, -1, -10, -4, 5, -28, 4, 4,
    -- layer=1 filter=8 channel=30
    -18, -41, -6, -31, -47, -52, -13, -38, -17,
    -- layer=1 filter=8 channel=31
    17, 4, 7, 9, -20, -20, -9, 3, 0,
    -- layer=1 filter=8 channel=32
    12, 52, 11, 4, 35, 4, 24, 46, 23,
    -- layer=1 filter=8 channel=33
    7, -14, -1, 4, 8, 11, 14, 26, 23,
    -- layer=1 filter=8 channel=34
    -4, 6, -5, -22, -10, -9, 0, -1, 8,
    -- layer=1 filter=8 channel=35
    0, 1, 3, 11, 8, -7, -4, -6, 7,
    -- layer=1 filter=8 channel=36
    11, 7, -10, 9, 0, -18, 6, 4, -20,
    -- layer=1 filter=8 channel=37
    -40, -34, -42, -56, -72, -43, -49, -110, -67,
    -- layer=1 filter=8 channel=38
    2, 2, 6, -8, 13, 1, -11, 4, 0,
    -- layer=1 filter=8 channel=39
    1, -6, -9, -4, -15, -6, -19, -19, -12,
    -- layer=1 filter=8 channel=40
    19, 19, 7, 7, -6, -6, -30, -9, -12,
    -- layer=1 filter=8 channel=41
    -16, -28, 20, -4, 14, -24, -9, -6, 2,
    -- layer=1 filter=8 channel=42
    57, 56, 10, 58, 27, 14, 34, 27, 6,
    -- layer=1 filter=8 channel=43
    -17, -12, -22, -32, -25, 6, -5, -56, -35,
    -- layer=1 filter=8 channel=44
    24, 64, -9, -7, 17, 0, 6, 39, 8,
    -- layer=1 filter=8 channel=45
    -6, 27, -7, -20, -14, 3, 9, -3, -13,
    -- layer=1 filter=8 channel=46
    -13, -16, -48, 17, -52, -12, 2, -29, 3,
    -- layer=1 filter=8 channel=47
    15, 0, 7, 62, 34, 10, 39, 44, 35,
    -- layer=1 filter=8 channel=48
    -4, -4, 0, -9, -11, 0, 3, -10, -4,
    -- layer=1 filter=8 channel=49
    22, 1, -8, 18, -3, -4, 9, -9, 12,
    -- layer=1 filter=8 channel=50
    -25, 9, 0, -6, -6, -3, -7, 9, 4,
    -- layer=1 filter=8 channel=51
    4, 3, 6, -3, 2, 1, -5, -15, 9,
    -- layer=1 filter=8 channel=52
    -2, 9, -9, 10, 14, 11, 1, -9, -10,
    -- layer=1 filter=8 channel=53
    0, 2, -5, -5, -2, 22, 5, -16, -1,
    -- layer=1 filter=8 channel=54
    2, 8, 7, -10, -24, -36, -10, 0, -4,
    -- layer=1 filter=8 channel=55
    20, -15, -17, 11, -7, -6, -4, -2, -24,
    -- layer=1 filter=8 channel=56
    6, 4, 1, 8, 4, 4, 13, 0, -3,
    -- layer=1 filter=8 channel=57
    24, 49, 16, 7, 37, 1, 8, 27, 8,
    -- layer=1 filter=8 channel=58
    46, 50, 32, 92, 58, 43, 76, 71, 46,
    -- layer=1 filter=8 channel=59
    8, -11, 1, 0, -1, -4, -5, -10, -8,
    -- layer=1 filter=8 channel=60
    -8, 7, -2, -11, -8, -2, -15, 4, -7,
    -- layer=1 filter=8 channel=61
    -1, -10, -11, 5, -5, -10, 3, 3, -7,
    -- layer=1 filter=8 channel=62
    -37, -31, -38, -67, -55, -16, -30, -91, -47,
    -- layer=1 filter=8 channel=63
    -3, -5, -2, -5, -6, -1, 7, -3, 1,
    -- layer=1 filter=8 channel=64
    -6, 5, 13, -14, 6, -6, -13, 3, 0,
    -- layer=1 filter=8 channel=65
    4, 2, 10, -1, -4, 6, -8, 2, 13,
    -- layer=1 filter=8 channel=66
    8, 8, 0, 5, 7, -1, 5, 9, -3,
    -- layer=1 filter=8 channel=67
    -40, -57, -14, -33, -46, 0, -7, -26, 1,
    -- layer=1 filter=8 channel=68
    38, 62, 9, 2, 52, -1, 30, 46, 8,
    -- layer=1 filter=8 channel=69
    -9, 31, -32, -30, -31, -5, 25, -21, -25,
    -- layer=1 filter=8 channel=70
    -20, -45, -15, -21, -41, -15, -16, -47, -12,
    -- layer=1 filter=8 channel=71
    -17, -26, -7, -1, -33, -6, -19, -22, 2,
    -- layer=1 filter=8 channel=72
    -25, -9, 3, -21, -63, -39, -2, -34, 7,
    -- layer=1 filter=8 channel=73
    -11, -1, 0, 5, -13, -12, -3, 6, -6,
    -- layer=1 filter=8 channel=74
    -4, 16, -14, -21, 9, -6, -19, 23, 1,
    -- layer=1 filter=8 channel=75
    -15, -1, -19, 15, -52, -37, -36, -49, -29,
    -- layer=1 filter=8 channel=76
    7, 14, -4, -6, 0, -32, -10, 8, -2,
    -- layer=1 filter=8 channel=77
    -14, -13, 1, -15, 5, 14, -7, -4, 6,
    -- layer=1 filter=8 channel=78
    -17, -7, -10, -13, -15, -30, -6, -8, -10,
    -- layer=1 filter=8 channel=79
    -34, -12, -39, -34, -39, -18, -25, -55, -22,
    -- layer=1 filter=8 channel=80
    4, -5, -8, 9, 1, 6, 0, -2, -11,
    -- layer=1 filter=8 channel=81
    0, -33, -13, -16, -32, 13, 12, -36, -17,
    -- layer=1 filter=8 channel=82
    -1, -7, 0, -18, 3, 21, 0, -1, 17,
    -- layer=1 filter=8 channel=83
    3, 36, -15, -29, -1, 9, -1, -20, -29,
    -- layer=1 filter=8 channel=84
    -17, -14, -8, -28, -17, -32, -18, -12, 0,
    -- layer=1 filter=8 channel=85
    10, 0, 17, 44, 18, 9, 49, 33, 21,
    -- layer=1 filter=8 channel=86
    5, 4, -16, 1, 3, -12, -5, 3, -12,
    -- layer=1 filter=8 channel=87
    10, -18, -3, 7, -20, -43, 17, -31, -11,
    -- layer=1 filter=8 channel=88
    6, -13, -9, -3, -18, 2, -1, -13, 9,
    -- layer=1 filter=8 channel=89
    -27, 0, 2, -23, -23, 1, 4, -8, 8,
    -- layer=1 filter=8 channel=90
    29, 40, 11, 5, 52, -1, 30, 39, 13,
    -- layer=1 filter=8 channel=91
    13, 7, 10, 2, -2, -10, -8, 4, 2,
    -- layer=1 filter=8 channel=92
    31, -17, -30, -21, -21, -73, 9, -12, -30,
    -- layer=1 filter=8 channel=93
    -11, -14, 1, -16, -14, 3, 0, -18, 3,
    -- layer=1 filter=8 channel=94
    12, 13, 12, 10, 6, 1, -3, -11, -1,
    -- layer=1 filter=8 channel=95
    -38, -24, -10, -25, -34, -42, -33, -36, -10,
    -- layer=1 filter=8 channel=96
    -8, -9, -1, -3, -10, -3, -16, -11, -10,
    -- layer=1 filter=8 channel=97
    2, -4, 3, -12, -3, 0, 4, 2, 2,
    -- layer=1 filter=8 channel=98
    -15, -26, -14, -24, -17, -6, -10, -50, -21,
    -- layer=1 filter=8 channel=99
    26, 38, 39, 9, 66, 45, 28, 55, 57,
    -- layer=1 filter=8 channel=100
    3, -5, 0, -7, -10, -20, -8, -11, 1,
    -- layer=1 filter=8 channel=101
    -7, 6, 7, -8, 12, 14, 0, 6, 6,
    -- layer=1 filter=8 channel=102
    22, 19, 2, 1, -6, -3, -8, -10, -24,
    -- layer=1 filter=8 channel=103
    -19, -21, -5, 0, -25, -12, -14, 7, 5,
    -- layer=1 filter=8 channel=104
    14, -26, 10, 59, -6, 12, 50, 14, 17,
    -- layer=1 filter=8 channel=105
    6, -10, -5, -1, 3, 3, 9, 0, 6,
    -- layer=1 filter=8 channel=106
    0, 7, 1, -13, 1, 8, 0, -1, 13,
    -- layer=1 filter=8 channel=107
    0, -4, 6, -3, -22, -5, -19, -7, -14,
    -- layer=1 filter=8 channel=108
    10, 38, 14, 8, 33, -3, 6, 34, 6,
    -- layer=1 filter=8 channel=109
    -5, 3, -7, -9, 0, 1, 1, 8, 6,
    -- layer=1 filter=8 channel=110
    -7, 0, -9, 5, -4, 3, 5, 2, 3,
    -- layer=1 filter=8 channel=111
    -27, -29, -7, -25, -26, -28, -21, -38, -29,
    -- layer=1 filter=8 channel=112
    -43, -9, -28, -10, -19, -4, -21, -34, 4,
    -- layer=1 filter=8 channel=113
    13, 25, 7, 0, 9, -9, 3, 5, 18,
    -- layer=1 filter=8 channel=114
    -19, -11, -57, -37, -68, -34, -26, -93, -88,
    -- layer=1 filter=8 channel=115
    0, 5, 8, 10, -10, -15, -14, -1, -11,
    -- layer=1 filter=8 channel=116
    -6, 0, 6, -9, 6, -8, -2, 0, 6,
    -- layer=1 filter=8 channel=117
    -33, -26, -14, -31, -10, 3, -21, -47, -20,
    -- layer=1 filter=8 channel=118
    -17, -17, 5, -13, 0, -32, -17, -4, -14,
    -- layer=1 filter=8 channel=119
    10, 34, -1, 16, 41, 0, 25, 46, 15,
    -- layer=1 filter=8 channel=120
    -4, -2, 9, 3, -10, -6, 1, -15, -4,
    -- layer=1 filter=8 channel=121
    14, -12, 8, 4, -11, -24, -21, -16, -10,
    -- layer=1 filter=8 channel=122
    -2, 2, 0, 6, 3, 10, -9, 7, 10,
    -- layer=1 filter=8 channel=123
    -6, -19, -19, 1, -7, -39, -17, -3, -12,
    -- layer=1 filter=8 channel=124
    12, 11, -3, 8, -7, 5, 1, 4, -8,
    -- layer=1 filter=8 channel=125
    -9, -9, 4, -6, -10, -18, -12, -7, -8,
    -- layer=1 filter=8 channel=126
    -37, -33, -22, -62, -48, 2, -35, -79, -49,
    -- layer=1 filter=8 channel=127
    -24, -3, 0, -11, -33, -24, -20, -29, -6,
    -- layer=1 filter=9 channel=0
    -4, 5, -10, 0, -2, 0, -7, -1, -7,
    -- layer=1 filter=9 channel=1
    -8, -6, -8, -10, -8, -9, 4, 7, -9,
    -- layer=1 filter=9 channel=2
    -3, -1, 2, -1, 1, -1, 2, 7, -6,
    -- layer=1 filter=9 channel=3
    5, 9, 2, -3, 6, 0, 1, 0, -3,
    -- layer=1 filter=9 channel=4
    -11, 1, 2, 5, -3, -4, -4, -4, -5,
    -- layer=1 filter=9 channel=5
    0, -8, 10, -2, -5, 0, 4, 2, -10,
    -- layer=1 filter=9 channel=6
    0, -7, 10, 5, -10, 3, -4, 8, 2,
    -- layer=1 filter=9 channel=7
    0, 7, 6, 8, -8, -11, 9, -10, -5,
    -- layer=1 filter=9 channel=8
    -11, 3, -12, -1, 9, -7, 0, -5, -8,
    -- layer=1 filter=9 channel=9
    -5, 9, 5, -6, -8, -12, 1, -2, 6,
    -- layer=1 filter=9 channel=10
    2, -1, -8, -10, -10, -3, 8, -12, -1,
    -- layer=1 filter=9 channel=11
    9, -7, -2, 4, 0, -9, 4, -8, 0,
    -- layer=1 filter=9 channel=12
    -3, 5, 0, 1, -5, -7, 1, 2, 3,
    -- layer=1 filter=9 channel=13
    -1, -10, 0, -2, 7, 10, -6, -2, -10,
    -- layer=1 filter=9 channel=14
    3, 0, 11, 8, 0, -2, 3, 5, 6,
    -- layer=1 filter=9 channel=15
    6, 6, 7, -1, -3, -9, 0, -2, -3,
    -- layer=1 filter=9 channel=16
    6, 6, -9, 7, -8, -10, -3, -6, -6,
    -- layer=1 filter=9 channel=17
    3, -10, -2, 1, 2, 8, 4, -7, 1,
    -- layer=1 filter=9 channel=18
    -7, -7, -8, 0, -6, -7, 5, -1, 8,
    -- layer=1 filter=9 channel=19
    0, 3, -3, -11, -4, 5, -8, 2, -6,
    -- layer=1 filter=9 channel=20
    -5, -5, -3, 7, -4, 0, -6, 0, 2,
    -- layer=1 filter=9 channel=21
    2, 6, 6, 0, -3, -9, 0, 2, 8,
    -- layer=1 filter=9 channel=22
    -9, 2, 5, 4, 2, -11, 4, -4, -8,
    -- layer=1 filter=9 channel=23
    9, -10, 3, 6, 0, -11, 1, 5, -2,
    -- layer=1 filter=9 channel=24
    7, -6, 4, -11, 0, 7, -2, -10, 2,
    -- layer=1 filter=9 channel=25
    1, 9, -2, -6, 10, -12, 5, -7, -1,
    -- layer=1 filter=9 channel=26
    -1, 0, 7, 2, 1, 9, 9, -4, 8,
    -- layer=1 filter=9 channel=27
    0, 1, -1, 0, -6, 2, 3, -2, 3,
    -- layer=1 filter=9 channel=28
    0, -7, -6, -5, 2, 7, -8, 6, -6,
    -- layer=1 filter=9 channel=29
    -11, 9, 7, 8, 6, 3, 0, 3, -1,
    -- layer=1 filter=9 channel=30
    -10, -6, 5, 7, 5, 2, 2, 2, -1,
    -- layer=1 filter=9 channel=31
    0, 4, -2, -3, -6, 1, 6, -11, -11,
    -- layer=1 filter=9 channel=32
    0, -1, 0, -1, 2, 6, -6, 0, 0,
    -- layer=1 filter=9 channel=33
    3, 1, 9, 4, -9, -7, 3, 1, 5,
    -- layer=1 filter=9 channel=34
    0, 0, -4, 6, -4, -9, 4, -6, -2,
    -- layer=1 filter=9 channel=35
    1, 0, -6, 0, -2, -7, -3, 0, -1,
    -- layer=1 filter=9 channel=36
    8, 9, 9, 1, -10, 4, -3, 0, -7,
    -- layer=1 filter=9 channel=37
    2, -3, 4, 2, -4, -11, -4, -1, -11,
    -- layer=1 filter=9 channel=38
    3, -6, 2, -1, -8, -7, -9, -11, -11,
    -- layer=1 filter=9 channel=39
    -12, -7, -4, 2, -3, 0, -8, 3, 8,
    -- layer=1 filter=9 channel=40
    9, 4, -8, -3, 4, 6, 5, 0, -4,
    -- layer=1 filter=9 channel=41
    -1, 4, 4, 8, -3, 6, -7, -5, 0,
    -- layer=1 filter=9 channel=42
    -11, -10, -8, -10, -9, 5, -5, -9, 3,
    -- layer=1 filter=9 channel=43
    -2, -6, 7, -3, 5, -2, -9, 4, -1,
    -- layer=1 filter=9 channel=44
    7, -1, -11, -5, -6, -12, 6, 0, -3,
    -- layer=1 filter=9 channel=45
    7, 2, 0, -4, 8, -2, 5, 1, 0,
    -- layer=1 filter=9 channel=46
    -8, 0, 7, 8, 0, -3, 7, 6, -3,
    -- layer=1 filter=9 channel=47
    2, -4, -8, 1, 2, -2, -7, 2, -3,
    -- layer=1 filter=9 channel=48
    3, 0, 0, -10, 2, -1, 1, -2, 0,
    -- layer=1 filter=9 channel=49
    0, -10, -4, 0, -8, 3, 5, 1, -9,
    -- layer=1 filter=9 channel=50
    5, -3, -2, -5, -11, -8, -3, -3, -3,
    -- layer=1 filter=9 channel=51
    6, 0, -4, 3, 6, 4, -2, 1, 7,
    -- layer=1 filter=9 channel=52
    10, -10, -3, -2, 3, -7, 9, -3, -8,
    -- layer=1 filter=9 channel=53
    -9, -2, -4, 0, -1, 0, 1, 0, 0,
    -- layer=1 filter=9 channel=54
    3, 7, 5, 8, -3, -5, -3, -3, -2,
    -- layer=1 filter=9 channel=55
    3, 0, 8, -4, 0, 0, -2, -4, 1,
    -- layer=1 filter=9 channel=56
    6, -2, 2, 4, 8, 0, 0, 7, -11,
    -- layer=1 filter=9 channel=57
    -9, -2, 6, 7, 2, -2, -8, -7, -7,
    -- layer=1 filter=9 channel=58
    -5, -4, 0, -7, -4, -1, -6, 6, -4,
    -- layer=1 filter=9 channel=59
    1, -8, 2, 0, 0, -3, 8, 8, -3,
    -- layer=1 filter=9 channel=60
    -5, -8, 8, 8, -6, 8, 4, -8, -4,
    -- layer=1 filter=9 channel=61
    -3, 6, 8, -2, 3, 5, 1, 0, -6,
    -- layer=1 filter=9 channel=62
    -1, 0, 8, -5, 2, 6, -6, 0, 1,
    -- layer=1 filter=9 channel=63
    -6, -8, 0, 3, 5, 4, 3, -1, -2,
    -- layer=1 filter=9 channel=64
    5, -6, -11, -11, -9, 6, 3, -7, -5,
    -- layer=1 filter=9 channel=65
    3, -3, 3, -7, -3, 5, -8, 1, -6,
    -- layer=1 filter=9 channel=66
    -11, -2, -1, -12, -5, 2, 3, -2, 6,
    -- layer=1 filter=9 channel=67
    4, -4, -9, 2, 5, -1, 7, -5, -7,
    -- layer=1 filter=9 channel=68
    -1, -9, -9, -9, 6, 0, 1, -4, 1,
    -- layer=1 filter=9 channel=69
    -4, 9, -5, 1, 3, 8, -12, -1, 0,
    -- layer=1 filter=9 channel=70
    0, -4, 6, 2, 0, -7, -1, 4, 7,
    -- layer=1 filter=9 channel=71
    -5, 4, 4, -2, -4, 3, 0, -2, 3,
    -- layer=1 filter=9 channel=72
    5, -4, -10, 8, -8, -9, -2, 7, -6,
    -- layer=1 filter=9 channel=73
    -6, -5, -9, -11, -4, -8, 5, -4, 5,
    -- layer=1 filter=9 channel=74
    1, 8, 1, 2, -6, -7, -4, -8, 7,
    -- layer=1 filter=9 channel=75
    -7, 2, 7, -6, 2, 1, -4, 7, -5,
    -- layer=1 filter=9 channel=76
    8, -12, 0, 3, 2, -1, -8, 9, 8,
    -- layer=1 filter=9 channel=77
    1, -2, -7, 2, -6, -3, -11, 0, 0,
    -- layer=1 filter=9 channel=78
    0, 0, 6, 7, 0, -6, -7, 9, 2,
    -- layer=1 filter=9 channel=79
    -1, -10, -8, -7, 1, 7, 6, -5, -2,
    -- layer=1 filter=9 channel=80
    8, -2, 7, 8, 10, 8, 7, -3, -10,
    -- layer=1 filter=9 channel=81
    -7, 2, -9, -2, 7, 4, -1, -11, -10,
    -- layer=1 filter=9 channel=82
    4, 2, -6, -6, -1, -5, -6, 7, 3,
    -- layer=1 filter=9 channel=83
    -8, 0, 3, 0, 6, -6, -11, 0, 0,
    -- layer=1 filter=9 channel=84
    -9, -7, -4, -8, 3, 1, 10, 0, 7,
    -- layer=1 filter=9 channel=85
    5, 6, -11, 3, 8, -11, 2, 1, 1,
    -- layer=1 filter=9 channel=86
    8, -3, 9, 7, -4, 0, -5, 2, 7,
    -- layer=1 filter=9 channel=87
    3, -9, 5, 8, 8, 2, 6, -3, -3,
    -- layer=1 filter=9 channel=88
    1, 3, 7, -7, -2, 4, 3, -7, -7,
    -- layer=1 filter=9 channel=89
    -4, -5, -9, 6, 3, -6, -6, 9, 2,
    -- layer=1 filter=9 channel=90
    -11, -11, -4, 3, 2, -5, -5, 5, 0,
    -- layer=1 filter=9 channel=91
    -6, -8, 0, -11, -12, 0, 0, -1, -8,
    -- layer=1 filter=9 channel=92
    0, -1, 8, -2, 8, 1, -9, 7, 9,
    -- layer=1 filter=9 channel=93
    -10, -9, -2, -8, -5, 4, -10, -4, -7,
    -- layer=1 filter=9 channel=94
    0, -1, 0, 5, 1, 2, -8, 3, 2,
    -- layer=1 filter=9 channel=95
    0, -3, -6, -10, 6, -5, 7, -1, 5,
    -- layer=1 filter=9 channel=96
    -6, 0, -1, 0, 2, -9, -3, 1, 3,
    -- layer=1 filter=9 channel=97
    -2, 3, -7, -4, -8, 3, -3, -4, 3,
    -- layer=1 filter=9 channel=98
    -6, 7, -4, -2, -9, 4, -10, -10, -9,
    -- layer=1 filter=9 channel=99
    5, -3, 8, -1, -8, -4, 3, 4, 6,
    -- layer=1 filter=9 channel=100
    -2, -7, -5, -4, -7, 3, -12, 4, -1,
    -- layer=1 filter=9 channel=101
    4, 6, 2, -10, 0, 4, 6, 6, -1,
    -- layer=1 filter=9 channel=102
    2, 2, 6, -10, -5, -2, -12, -9, -8,
    -- layer=1 filter=9 channel=103
    5, -4, 5, -6, 4, 5, -4, -1, -2,
    -- layer=1 filter=9 channel=104
    0, -9, 2, -10, -4, -3, -10, -11, 4,
    -- layer=1 filter=9 channel=105
    -8, 6, -4, -11, 6, -2, 1, -1, -7,
    -- layer=1 filter=9 channel=106
    7, 5, 0, -5, 4, -9, 0, -7, 9,
    -- layer=1 filter=9 channel=107
    -1, -2, -6, 1, 3, 3, 1, 5, -4,
    -- layer=1 filter=9 channel=108
    0, 6, 7, 6, -2, 0, -10, -7, -3,
    -- layer=1 filter=9 channel=109
    -4, -8, 0, 4, -4, 0, 7, 0, -3,
    -- layer=1 filter=9 channel=110
    -5, 0, -10, -8, -2, -9, -7, -5, -5,
    -- layer=1 filter=9 channel=111
    8, -6, -5, 7, -7, -5, -3, -1, -2,
    -- layer=1 filter=9 channel=112
    2, -8, -6, 0, 7, -1, 0, -3, -10,
    -- layer=1 filter=9 channel=113
    -6, -3, 5, 1, 0, -3, 7, 3, -6,
    -- layer=1 filter=9 channel=114
    1, 4, 0, 0, -10, -1, -1, 1, -2,
    -- layer=1 filter=9 channel=115
    2, -9, -8, -4, -8, -10, 0, 0, -10,
    -- layer=1 filter=9 channel=116
    10, -1, 3, 8, -10, 1, 0, 1, 4,
    -- layer=1 filter=9 channel=117
    -8, 9, 2, -6, 4, 0, -6, -8, -10,
    -- layer=1 filter=9 channel=118
    -7, 4, -7, -3, -9, 0, -9, -8, 0,
    -- layer=1 filter=9 channel=119
    -6, -9, -5, 7, 6, -7, 4, 2, 3,
    -- layer=1 filter=9 channel=120
    2, 6, 7, -7, -13, 0, 7, -1, -1,
    -- layer=1 filter=9 channel=121
    -2, 2, -9, -6, -11, -1, 0, -9, 0,
    -- layer=1 filter=9 channel=122
    -3, 0, 6, 3, 9, 3, -3, -7, 4,
    -- layer=1 filter=9 channel=123
    2, 8, -3, -12, -5, -1, -10, 0, 7,
    -- layer=1 filter=9 channel=124
    0, -9, -6, -5, 11, 3, 4, 0, 0,
    -- layer=1 filter=9 channel=125
    2, 2, 3, -10, -7, 8, 5, 5, 2,
    -- layer=1 filter=9 channel=126
    8, 6, 8, -10, -5, 2, 1, -4, -3,
    -- layer=1 filter=9 channel=127
    -4, 5, 5, 7, 6, 9, -10, 0, 0,
    -- layer=1 filter=10 channel=0
    4, 15, 5, 0, -8, 10, 0, -15, -5,
    -- layer=1 filter=10 channel=1
    25, 41, 31, 8, 15, -1, -19, 12, -22,
    -- layer=1 filter=10 channel=2
    -74, -75, -29, -4, -11, -26, 0, 2, -8,
    -- layer=1 filter=10 channel=3
    0, -2, -4, -6, -2, -4, 11, -3, 7,
    -- layer=1 filter=10 channel=4
    3, -7, 13, -4, -2, 8, -2, -6, 5,
    -- layer=1 filter=10 channel=5
    -11, 5, -13, 13, 32, 0, 17, 20, -25,
    -- layer=1 filter=10 channel=6
    28, 33, 27, 4, 0, 3, -32, -55, -21,
    -- layer=1 filter=10 channel=7
    2, -26, -33, 5, 10, 1, -1, -8, 18,
    -- layer=1 filter=10 channel=8
    24, 37, 5, -18, -13, -13, -4, 16, -19,
    -- layer=1 filter=10 channel=9
    29, -18, -24, 3, -35, 23, -35, -39, -32,
    -- layer=1 filter=10 channel=10
    20, -1, -23, 0, 35, 36, 3, 3, 29,
    -- layer=1 filter=10 channel=11
    -20, -25, 1, 3, 7, -5, 21, 22, -3,
    -- layer=1 filter=10 channel=12
    -2, -23, -28, 25, 38, -56, -51, -22, 18,
    -- layer=1 filter=10 channel=13
    9, 35, 34, -18, -17, 10, -14, -60, -25,
    -- layer=1 filter=10 channel=14
    -21, -47, -23, 2, 49, -15, -22, -2, 40,
    -- layer=1 filter=10 channel=15
    -36, 14, 31, -13, -7, -46, 18, 15, 2,
    -- layer=1 filter=10 channel=16
    -6, 2, -10, -5, -25, -16, 5, 18, -36,
    -- layer=1 filter=10 channel=17
    25, 36, 13, -21, -24, -16, -18, -25, -24,
    -- layer=1 filter=10 channel=18
    22, -9, 20, 3, 53, 1, -27, 1, 5,
    -- layer=1 filter=10 channel=19
    27, 10, -17, 54, 40, 47, 14, 31, -26,
    -- layer=1 filter=10 channel=20
    11, 41, 16, -12, -23, 11, -42, -40, -41,
    -- layer=1 filter=10 channel=21
    29, 34, 48, -9, -9, -10, -54, -57, -44,
    -- layer=1 filter=10 channel=22
    31, 54, 34, -29, -20, -6, -46, -43, -41,
    -- layer=1 filter=10 channel=23
    -12, -6, 23, 7, -4, 3, 0, 21, 8,
    -- layer=1 filter=10 channel=24
    10, 16, 9, -7, -18, 13, 0, -20, -35,
    -- layer=1 filter=10 channel=25
    -11, -13, -20, -20, -8, 11, 16, 14, -13,
    -- layer=1 filter=10 channel=26
    -21, -9, 12, -2, -11, -7, 20, -26, -29,
    -- layer=1 filter=10 channel=27
    -27, -31, -1, -21, -10, 0, -1, 22, 24,
    -- layer=1 filter=10 channel=28
    9, -14, -2, -28, -12, -11, -11, -19, 7,
    -- layer=1 filter=10 channel=29
    -19, -5, 13, -26, 9, 9, -1, -8, -2,
    -- layer=1 filter=10 channel=30
    18, -6, -11, 10, 59, 21, -26, -28, 2,
    -- layer=1 filter=10 channel=31
    17, -1, 4, 15, 53, 1, -34, -16, 0,
    -- layer=1 filter=10 channel=32
    0, -24, 10, 32, 4, 8, 27, -11, -13,
    -- layer=1 filter=10 channel=33
    12, 5, 6, 1, -7, -9, -9, 4, -15,
    -- layer=1 filter=10 channel=34
    6, 5, 6, 12, -1, -5, 1, -11, -10,
    -- layer=1 filter=10 channel=35
    -11, -3, -18, -2, -16, -8, -6, 4, -2,
    -- layer=1 filter=10 channel=36
    -11, -17, -6, 2, 11, -6, 30, 22, 11,
    -- layer=1 filter=10 channel=37
    -11, 6, -14, 34, 14, 13, 19, 14, -31,
    -- layer=1 filter=10 channel=38
    40, 36, 18, -21, -3, 9, -58, -53, -42,
    -- layer=1 filter=10 channel=39
    3, -16, 0, -21, -18, -17, 2, 9, 0,
    -- layer=1 filter=10 channel=40
    29, 9, 0, -1, 13, 2, -54, -52, -25,
    -- layer=1 filter=10 channel=41
    0, -59, -17, 7, 2, 13, 27, -27, -15,
    -- layer=1 filter=10 channel=42
    -90, -46, -29, -2, 11, -38, -25, -16, -12,
    -- layer=1 filter=10 channel=43
    21, 19, 5, -24, -19, -32, -1, 12, -33,
    -- layer=1 filter=10 channel=44
    -12, 14, 18, 16, 0, -3, 19, -9, 11,
    -- layer=1 filter=10 channel=45
    17, 42, 32, -6, 12, -3, -22, -15, -25,
    -- layer=1 filter=10 channel=46
    22, -2, 9, 79, 75, -3, -18, 15, -3,
    -- layer=1 filter=10 channel=47
    5, 3, 37, 25, 3, 35, -4, -9, -24,
    -- layer=1 filter=10 channel=48
    45, 35, 14, -9, 0, 18, -50, -48, -25,
    -- layer=1 filter=10 channel=49
    32, 33, 4, 13, 0, 22, -27, -49, -28,
    -- layer=1 filter=10 channel=50
    1, 0, -1, -16, -12, 4, -9, -18, -12,
    -- layer=1 filter=10 channel=51
    39, 22, 13, -3, 9, 10, -51, -57, -16,
    -- layer=1 filter=10 channel=52
    -13, -15, -13, -18, 1, -12, -19, -12, 0,
    -- layer=1 filter=10 channel=53
    -5, 2, 4, 7, 4, -2, -13, -5, -1,
    -- layer=1 filter=10 channel=54
    -28, -32, -57, 7, 4, 12, 28, 18, -19,
    -- layer=1 filter=10 channel=55
    -22, -35, -24, -1, -1, -12, 36, 43, 6,
    -- layer=1 filter=10 channel=56
    8, 1, 2, -5, -1, -8, -5, 0, -8,
    -- layer=1 filter=10 channel=57
    13, 11, 1, 12, 20, 27, -9, -24, 8,
    -- layer=1 filter=10 channel=58
    31, 1, -33, -7, 12, 38, -7, -15, 17,
    -- layer=1 filter=10 channel=59
    12, -10, 5, -11, -8, 0, -4, 4, -6,
    -- layer=1 filter=10 channel=60
    9, 1, 4, 13, -5, 0, 0, -9, 11,
    -- layer=1 filter=10 channel=61
    7, 4, 1, 0, -5, -2, -6, -2, 5,
    -- layer=1 filter=10 channel=62
    14, 34, 0, -10, 5, 12, 11, 22, -27,
    -- layer=1 filter=10 channel=63
    -7, -14, 0, 7, 13, -14, 8, 8, -4,
    -- layer=1 filter=10 channel=64
    24, 4, 26, -7, -10, 10, -30, -30, -25,
    -- layer=1 filter=10 channel=65
    30, 31, 24, -16, -16, 11, -39, -35, -15,
    -- layer=1 filter=10 channel=66
    -12, -6, 7, 4, 9, -10, 13, 17, 15,
    -- layer=1 filter=10 channel=67
    72, 68, 58, 47, 56, 68, -38, -54, -6,
    -- layer=1 filter=10 channel=68
    -36, -2, 20, 7, -6, -13, 6, -19, 4,
    -- layer=1 filter=10 channel=69
    -10, 14, -4, -18, -11, -15, 21, 23, -20,
    -- layer=1 filter=10 channel=70
    40, 28, -10, 28, 38, 19, -3, 2, -9,
    -- layer=1 filter=10 channel=71
    12, 5, 6, 1, 16, -4, -9, -2, 5,
    -- layer=1 filter=10 channel=72
    2, -14, -10, 25, 22, -2, -17, -7, -23,
    -- layer=1 filter=10 channel=73
    -4, -5, -1, 0, 8, -7, -4, 1, 0,
    -- layer=1 filter=10 channel=74
    0, -23, 24, 2, 29, 2, -42, -44, -3,
    -- layer=1 filter=10 channel=75
    13, -47, 13, 10, 69, -49, -36, 10, 38,
    -- layer=1 filter=10 channel=76
    0, -1, 4, 7, 6, 0, 7, -30, -26,
    -- layer=1 filter=10 channel=77
    45, 66, 45, -8, -1, 15, -21, -37, -36,
    -- layer=1 filter=10 channel=78
    1, -6, -13, -16, 9, 1, 8, -5, 0,
    -- layer=1 filter=10 channel=79
    13, 21, -4, -20, -8, -4, 12, 16, -25,
    -- layer=1 filter=10 channel=80
    3, 0, -6, -6, -3, -3, 2, 14, 4,
    -- layer=1 filter=10 channel=81
    28, 25, 21, -19, -19, 0, -2, -16, -15,
    -- layer=1 filter=10 channel=82
    48, 56, 41, -16, -10, 3, -56, -70, -49,
    -- layer=1 filter=10 channel=83
    -1, 39, 21, -5, -5, -6, -10, -18, -14,
    -- layer=1 filter=10 channel=84
    31, -13, 34, 17, 25, -10, -11, -13, -11,
    -- layer=1 filter=10 channel=85
    21, 13, 11, 13, 5, 43, 23, 16, -6,
    -- layer=1 filter=10 channel=86
    -15, -14, -12, 0, 5, -15, 5, 25, 10,
    -- layer=1 filter=10 channel=87
    -4, -15, -45, 41, 19, 25, -34, 8, -40,
    -- layer=1 filter=10 channel=88
    33, 34, 22, 0, 0, 11, -39, -34, -22,
    -- layer=1 filter=10 channel=89
    16, 37, 34, -7, 0, -16, -64, -59, -45,
    -- layer=1 filter=10 channel=90
    -20, 13, 10, -15, -7, -7, 34, 5, 6,
    -- layer=1 filter=10 channel=91
    12, 30, 16, 2, -6, 4, -58, -69, -37,
    -- layer=1 filter=10 channel=92
    -62, -8, 33, 35, 8, 23, 50, 7, -9,
    -- layer=1 filter=10 channel=93
    23, 19, 16, -13, -22, -9, -29, -30, -25,
    -- layer=1 filter=10 channel=94
    10, 0, -5, 1, 9, -5, -12, -14, -5,
    -- layer=1 filter=10 channel=95
    34, -14, 12, 37, 43, -1, -21, -5, 22,
    -- layer=1 filter=10 channel=96
    18, 3, 0, 1, -13, -7, 4, -6, -6,
    -- layer=1 filter=10 channel=97
    6, 20, 7, -6, -26, -8, -10, -7, -4,
    -- layer=1 filter=10 channel=98
    46, 55, 7, -26, 3, -8, -4, -1, -34,
    -- layer=1 filter=10 channel=99
    17, -2, 7, -24, 13, 32, -28, -36, 2,
    -- layer=1 filter=10 channel=100
    -7, -40, 2, 27, 26, -8, 4, 14, 12,
    -- layer=1 filter=10 channel=101
    25, 36, 17, -4, 7, 9, -55, -72, -23,
    -- layer=1 filter=10 channel=102
    10, 8, 1, 12, 21, 20, -50, -45, -14,
    -- layer=1 filter=10 channel=103
    2, 0, 11, 8, 26, 16, 9, 18, 5,
    -- layer=1 filter=10 channel=104
    9, -1, 9, 4, -12, 26, -2, 0, -7,
    -- layer=1 filter=10 channel=105
    2, 11, 8, -14, -10, 2, 1, -11, -7,
    -- layer=1 filter=10 channel=106
    19, 30, 32, -12, -2, -5, -30, -60, -36,
    -- layer=1 filter=10 channel=107
    -6, -8, -8, 8, -8, 11, -1, 4, 1,
    -- layer=1 filter=10 channel=108
    -9, -14, -11, -7, -19, -2, 29, 3, -17,
    -- layer=1 filter=10 channel=109
    -2, 7, -1, -5, 8, -2, 4, -5, 7,
    -- layer=1 filter=10 channel=110
    9, 13, -6, -2, -3, 5, -9, -18, 1,
    -- layer=1 filter=10 channel=111
    36, -6, 1, -15, 38, 14, -47, -47, 0,
    -- layer=1 filter=10 channel=112
    44, 28, 30, 16, 9, -23, -19, -7, 9,
    -- layer=1 filter=10 channel=113
    11, 7, 8, 4, 16, -11, -25, -32, -23,
    -- layer=1 filter=10 channel=114
    -40, -29, -27, -8, -39, -25, 18, 44, -18,
    -- layer=1 filter=10 channel=115
    1, -17, -8, -12, 2, 7, 8, -7, 22,
    -- layer=1 filter=10 channel=116
    -9, 3, -3, 6, 8, 1, -10, 8, 7,
    -- layer=1 filter=10 channel=117
    76, 55, 33, 20, 37, 19, -19, -10, 35,
    -- layer=1 filter=10 channel=118
    18, -9, 6, -9, 40, 16, -19, -36, -11,
    -- layer=1 filter=10 channel=119
    -15, -3, 6, 9, 3, 11, 30, -19, -18,
    -- layer=1 filter=10 channel=120
    31, 30, 9, -3, 0, 3, -32, -49, -26,
    -- layer=1 filter=10 channel=121
    -3, -13, -29, 23, 74, 12, -1, 15, 26,
    -- layer=1 filter=10 channel=122
    -3, 7, -2, 9, -9, -3, 9, 4, 2,
    -- layer=1 filter=10 channel=123
    -25, -47, -39, 13, 39, 9, -6, 27, 23,
    -- layer=1 filter=10 channel=124
    -7, -2, -3, 3, -8, -19, 8, -4, -10,
    -- layer=1 filter=10 channel=125
    44, 29, 14, 23, 43, 38, -19, -37, -23,
    -- layer=1 filter=10 channel=126
    71, 106, 50, 49, 34, 31, -25, -28, -42,
    -- layer=1 filter=10 channel=127
    21, -12, 1, 14, 43, 0, -21, -5, 17,
    -- layer=1 filter=11 channel=0
    6, -13, 0, -1, -8, -11, -12, 0, -9,
    -- layer=1 filter=11 channel=1
    29, -1, 8, -4, -10, 16, 39, -5, -14,
    -- layer=1 filter=11 channel=2
    -12, -7, -20, -27, -26, -17, 29, 18, 11,
    -- layer=1 filter=11 channel=3
    1, -1, -2, 4, 0, -2, 6, 12, 5,
    -- layer=1 filter=11 channel=4
    5, 7, 0, 7, 2, -1, -5, 5, 4,
    -- layer=1 filter=11 channel=5
    31, 18, 29, -1, 21, 22, 24, -8, -21,
    -- layer=1 filter=11 channel=6
    -40, -50, -33, -76, -75, -87, -49, -27, -9,
    -- layer=1 filter=11 channel=7
    -15, -12, 9, 12, -31, 21, 16, -17, 20,
    -- layer=1 filter=11 channel=8
    21, 9, 15, 0, 21, 30, 34, 16, 1,
    -- layer=1 filter=11 channel=9
    -63, -48, 0, 24, 6, 4, -33, -17, -4,
    -- layer=1 filter=11 channel=10
    -15, -17, 23, 28, -21, -4, -4, -8, 30,
    -- layer=1 filter=11 channel=11
    15, 17, 2, 16, 5, -7, -13, 7, 0,
    -- layer=1 filter=11 channel=12
    -41, -7, -10, 0, -34, -45, -22, 18, 14,
    -- layer=1 filter=11 channel=13
    -34, -22, -28, -32, -15, -27, 1, 0, -9,
    -- layer=1 filter=11 channel=14
    -36, -15, 3, 18, -30, 0, 16, 17, 26,
    -- layer=1 filter=11 channel=15
    -35, -46, -25, -19, -26, -7, 27, -15, -10,
    -- layer=1 filter=11 channel=16
    4, -3, -15, 5, 15, 10, 20, -7, -9,
    -- layer=1 filter=11 channel=17
    1, -4, 4, -20, 0, -2, -18, -7, 8,
    -- layer=1 filter=11 channel=18
    14, 24, 37, 36, -1, -3, 14, 38, 12,
    -- layer=1 filter=11 channel=19
    6, 3, 35, 70, 44, 25, -5, 9, 8,
    -- layer=1 filter=11 channel=20
    -28, -12, -29, -33, -9, -6, -13, -16, -23,
    -- layer=1 filter=11 channel=21
    -42, -28, -53, -43, -30, -27, -4, -10, -25,
    -- layer=1 filter=11 channel=22
    -7, -25, -31, -23, -16, -10, 37, 22, 13,
    -- layer=1 filter=11 channel=23
    -11, -26, 19, -12, -30, 17, 24, -15, 11,
    -- layer=1 filter=11 channel=24
    -10, -19, -13, -12, 1, 12, -21, -20, -25,
    -- layer=1 filter=11 channel=25
    -20, -27, -8, 20, -2, 16, 5, -27, 1,
    -- layer=1 filter=11 channel=26
    -14, 0, 0, -20, 7, 0, 17, -5, 7,
    -- layer=1 filter=11 channel=27
    -32, -37, -24, -19, -41, -39, -22, -18, -36,
    -- layer=1 filter=11 channel=28
    -24, -18, -21, 7, -23, 0, 8, -6, 24,
    -- layer=1 filter=11 channel=29
    -39, -43, -31, -35, -29, -45, -12, -28, -20,
    -- layer=1 filter=11 channel=30
    13, 22, 51, 31, 17, -7, 2, 30, 30,
    -- layer=1 filter=11 channel=31
    -22, -14, -17, 12, -20, -41, 0, 21, -1,
    -- layer=1 filter=11 channel=32
    -10, 9, 24, -10, 0, -30, 6, -14, -12,
    -- layer=1 filter=11 channel=33
    -4, 6, -7, 0, 6, -3, 11, 2, 0,
    -- layer=1 filter=11 channel=34
    0, -6, 6, 6, -9, -6, -4, -11, 7,
    -- layer=1 filter=11 channel=35
    -5, -5, -5, 0, -2, 0, -5, -3, -14,
    -- layer=1 filter=11 channel=36
    23, 14, 18, 14, 12, 8, 0, 7, 7,
    -- layer=1 filter=11 channel=37
    29, 24, 12, 29, 28, 35, 9, -19, -9,
    -- layer=1 filter=11 channel=38
    -19, -26, -25, -15, -26, -35, -19, -13, -9,
    -- layer=1 filter=11 channel=39
    -5, -14, -6, -5, -6, -3, 3, -8, 2,
    -- layer=1 filter=11 channel=40
    -37, -10, -26, 6, -26, -28, 20, 34, -1,
    -- layer=1 filter=11 channel=41
    -2, -29, 18, 4, -10, -21, 7, -27, -13,
    -- layer=1 filter=11 channel=42
    -24, -38, -28, 11, -14, -34, 33, -5, -7,
    -- layer=1 filter=11 channel=43
    17, -9, -6, -11, -10, 18, 21, 4, -10,
    -- layer=1 filter=11 channel=44
    -16, 8, 11, -18, -1, -3, 4, 1, 3,
    -- layer=1 filter=11 channel=45
    -27, -29, -12, -45, -14, -16, -10, -16, -14,
    -- layer=1 filter=11 channel=46
    17, 15, 53, 51, 49, 42, 22, 13, 18,
    -- layer=1 filter=11 channel=47
    -15, -49, 25, 10, -39, -2, 27, -40, -7,
    -- layer=1 filter=11 channel=48
    -20, -27, -14, -13, -29, -17, -18, -10, 0,
    -- layer=1 filter=11 channel=49
    -14, -13, -5, -14, -32, -16, -18, -9, -9,
    -- layer=1 filter=11 channel=50
    -2, -13, 9, -4, -12, 3, -19, -27, 4,
    -- layer=1 filter=11 channel=51
    -21, -29, -10, -21, -52, -32, -7, -33, -1,
    -- layer=1 filter=11 channel=52
    8, -7, 0, 5, 5, 4, 18, 12, 29,
    -- layer=1 filter=11 channel=53
    0, -4, -1, -8, -9, -17, -15, -9, -19,
    -- layer=1 filter=11 channel=54
    -7, -15, -16, 22, -4, 13, -1, -27, 5,
    -- layer=1 filter=11 channel=55
    19, 15, 0, 11, 13, 6, 5, 3, 0,
    -- layer=1 filter=11 channel=56
    -4, -9, 1, 6, -9, -9, -1, 4, 4,
    -- layer=1 filter=11 channel=57
    -17, -28, 5, 15, -26, -22, 5, -18, 19,
    -- layer=1 filter=11 channel=58
    -34, -60, 14, 21, -45, 13, 28, -58, 21,
    -- layer=1 filter=11 channel=59
    4, 4, -4, -7, 3, 0, 9, -2, -7,
    -- layer=1 filter=11 channel=60
    2, 17, 5, 17, 5, 8, 12, 13, 11,
    -- layer=1 filter=11 channel=61
    -2, -6, -2, -8, 0, -2, 0, 11, 8,
    -- layer=1 filter=11 channel=62
    29, 14, 3, 25, 21, 33, 22, 7, -12,
    -- layer=1 filter=11 channel=63
    8, 5, 7, 16, -2, -10, 6, 14, -8,
    -- layer=1 filter=11 channel=64
    0, -5, -10, -11, -12, -13, 0, 1, -7,
    -- layer=1 filter=11 channel=65
    -19, -5, -23, -16, -9, -4, -17, -18, -27,
    -- layer=1 filter=11 channel=66
    9, -2, -6, -6, -2, 3, -3, -14, -5,
    -- layer=1 filter=11 channel=67
    -12, -8, 1, -11, -13, -11, -25, -24, -16,
    -- layer=1 filter=11 channel=68
    -7, 3, -3, -27, 7, -4, 5, 18, 19,
    -- layer=1 filter=11 channel=69
    6, -8, -15, -7, 12, 13, 15, 1, -20,
    -- layer=1 filter=11 channel=70
    16, 13, 26, -25, -33, -27, -40, -19, -33,
    -- layer=1 filter=11 channel=71
    -7, -8, -1, -13, -2, 5, -8, -17, -8,
    -- layer=1 filter=11 channel=72
    0, 0, 34, 31, 0, -22, -5, 8, 16,
    -- layer=1 filter=11 channel=73
    -5, -8, -5, -6, 8, 3, 6, 0, 5,
    -- layer=1 filter=11 channel=74
    -29, 10, -10, -4, -21, -36, -20, 4, 0,
    -- layer=1 filter=11 channel=75
    1, 21, 28, 11, 1, -40, 16, 44, 19,
    -- layer=1 filter=11 channel=76
    3, 15, -2, 7, 6, -18, 1, 0, 3,
    -- layer=1 filter=11 channel=77
    -1, 14, 2, -14, -10, -6, -13, -3, -10,
    -- layer=1 filter=11 channel=78
    1, 10, -7, 6, -3, 4, -2, -2, 6,
    -- layer=1 filter=11 channel=79
    16, -1, -3, 20, 14, 26, 3, -4, -18,
    -- layer=1 filter=11 channel=80
    -7, 0, 10, -3, -3, -8, 11, 0, -3,
    -- layer=1 filter=11 channel=81
    -4, -27, -23, -13, 0, 2, 4, -13, -11,
    -- layer=1 filter=11 channel=82
    -9, -20, -13, -37, -34, -24, 0, -18, -19,
    -- layer=1 filter=11 channel=83
    -2, -19, -2, -29, -1, -2, -3, 12, -7,
    -- layer=1 filter=11 channel=84
    1, 17, 27, 15, 6, -8, 14, 40, 22,
    -- layer=1 filter=11 channel=85
    -12, -53, 15, 10, -23, 26, 27, -51, 24,
    -- layer=1 filter=11 channel=86
    8, 8, 8, -6, 9, -4, -13, -9, -7,
    -- layer=1 filter=11 channel=87
    -41, -13, 36, 43, -1, -8, -36, -15, 12,
    -- layer=1 filter=11 channel=88
    -3, -14, -8, -7, -8, -17, -15, -5, -13,
    -- layer=1 filter=11 channel=89
    -26, -20, -17, -41, -38, -34, 6, 0, -15,
    -- layer=1 filter=11 channel=90
    -26, -12, -17, -43, 18, -9, -8, 1, -11,
    -- layer=1 filter=11 channel=91
    -20, -23, -15, -21, -56, -49, -18, -13, -19,
    -- layer=1 filter=11 channel=92
    -50, -32, -8, -28, -50, -15, -5, -17, 0,
    -- layer=1 filter=11 channel=93
    0, -14, -10, -9, -7, 1, -10, -23, -9,
    -- layer=1 filter=11 channel=94
    2, -2, 11, -2, -3, 1, -5, -2, 11,
    -- layer=1 filter=11 channel=95
    13, 21, 39, 39, 8, 1, 22, 51, 20,
    -- layer=1 filter=11 channel=96
    0, -10, -7, 5, -4, 7, -5, 2, -8,
    -- layer=1 filter=11 channel=97
    -5, 1, 5, 3, 9, 12, 0, -12, -1,
    -- layer=1 filter=11 channel=98
    20, 2, 0, -15, -11, -4, 27, 0, 5,
    -- layer=1 filter=11 channel=99
    -28, -34, -26, 18, -8, -7, 0, 47, 32,
    -- layer=1 filter=11 channel=100
    1, 17, 13, -3, -10, -23, 0, -4, -11,
    -- layer=1 filter=11 channel=101
    -4, -7, -15, -35, -39, -39, -4, -7, -8,
    -- layer=1 filter=11 channel=102
    -9, 0, 4, -4, -20, -13, -5, -13, 0,
    -- layer=1 filter=11 channel=103
    -3, -4, 9, 3, -8, 1, 8, 4, 3,
    -- layer=1 filter=11 channel=104
    -30, -25, 1, -2, -16, -1, -10, -15, -14,
    -- layer=1 filter=11 channel=105
    1, 4, -1, 11, 6, 4, -12, 1, 3,
    -- layer=1 filter=11 channel=106
    -43, -4, -18, -45, -35, -45, -16, -9, -12,
    -- layer=1 filter=11 channel=107
    5, 7, 3, -24, -6, -19, -7, 0, -12,
    -- layer=1 filter=11 channel=108
    -24, -31, 4, -22, -1, -8, 4, -17, -12,
    -- layer=1 filter=11 channel=109
    5, -1, -11, 9, -7, 10, -7, -6, 3,
    -- layer=1 filter=11 channel=110
    -1, -2, -1, 2, 4, -11, -6, 5, -10,
    -- layer=1 filter=11 channel=111
    17, 2, 37, 24, -7, -9, 12, 40, 29,
    -- layer=1 filter=11 channel=112
    14, 20, 0, 15, -17, 2, 22, 52, 18,
    -- layer=1 filter=11 channel=113
    0, -24, -38, 4, -23, -65, 26, -18, -21,
    -- layer=1 filter=11 channel=114
    7, 1, -10, -5, 7, 12, 18, -8, -14,
    -- layer=1 filter=11 channel=115
    11, 1, 16, 16, -5, 8, -5, -6, 13,
    -- layer=1 filter=11 channel=116
    2, 9, -9, -11, 3, 0, -6, -5, -6,
    -- layer=1 filter=11 channel=117
    39, 15, 37, 45, 2, 18, 46, 54, 54,
    -- layer=1 filter=11 channel=118
    0, 6, 15, 15, 11, -17, -5, 27, 10,
    -- layer=1 filter=11 channel=119
    -11, 2, -1, -24, 28, -20, 9, -13, -11,
    -- layer=1 filter=11 channel=120
    -5, -15, -17, -22, -22, -21, 6, -39, -15,
    -- layer=1 filter=11 channel=121
    -18, 12, 18, 21, 8, -13, 6, 31, 12,
    -- layer=1 filter=11 channel=122
    -1, 0, -4, 9, -8, 6, 10, -1, 7,
    -- layer=1 filter=11 channel=123
    -10, 10, 5, 22, 12, -4, 0, 21, 0,
    -- layer=1 filter=11 channel=124
    2, 3, 4, -10, -11, 3, -11, -3, -12,
    -- layer=1 filter=11 channel=125
    39, 22, 29, -28, -10, -55, -30, -58, -30,
    -- layer=1 filter=11 channel=126
    23, 10, 41, 1, 5, -1, 67, 46, 41,
    -- layer=1 filter=11 channel=127
    10, 32, 41, 36, 0, -17, 19, 38, 15,
    -- layer=1 filter=12 channel=0
    1, -6, 0, 6, -12, 4, -9, -11, 0,
    -- layer=1 filter=12 channel=1
    5, 5, 1, -3, -2, -3, -9, 2, -5,
    -- layer=1 filter=12 channel=2
    2, -13, 2, -3, 3, -1, 6, -5, 2,
    -- layer=1 filter=12 channel=3
    -5, -4, 10, -9, 5, 10, -5, 3, 7,
    -- layer=1 filter=12 channel=4
    2, 5, 5, 2, 1, -2, -3, 3, -9,
    -- layer=1 filter=12 channel=5
    -1, 5, -2, 3, -8, 7, -9, 7, 6,
    -- layer=1 filter=12 channel=6
    -2, 1, -7, -8, -3, 2, -6, 7, 3,
    -- layer=1 filter=12 channel=7
    -8, -1, 6, -10, -2, 0, -8, 1, 6,
    -- layer=1 filter=12 channel=8
    2, -1, 0, -8, -8, 6, -2, 0, -5,
    -- layer=1 filter=12 channel=9
    -8, 4, -5, 4, 9, -9, 0, -7, -4,
    -- layer=1 filter=12 channel=10
    9, 0, 6, -8, 9, 0, 3, -4, 7,
    -- layer=1 filter=12 channel=11
    -1, -9, -8, -3, 0, -6, 0, -9, -5,
    -- layer=1 filter=12 channel=12
    0, 2, 10, 9, 4, 5, 1, -4, -4,
    -- layer=1 filter=12 channel=13
    1, 0, -6, 0, -12, -5, -4, 4, -5,
    -- layer=1 filter=12 channel=14
    0, 5, -3, 9, 0, 0, -7, -1, 6,
    -- layer=1 filter=12 channel=15
    0, -5, 6, -5, -11, -3, 7, 8, 6,
    -- layer=1 filter=12 channel=16
    0, -3, 2, -6, -11, -5, -6, -4, -11,
    -- layer=1 filter=12 channel=17
    8, -2, -7, 8, 3, -11, 0, 6, 7,
    -- layer=1 filter=12 channel=18
    -1, -1, 4, 6, 6, -8, -7, -7, 10,
    -- layer=1 filter=12 channel=19
    3, 2, -11, -4, 2, 5, -7, 0, 0,
    -- layer=1 filter=12 channel=20
    5, 1, -10, -6, 6, 3, 0, 2, 5,
    -- layer=1 filter=12 channel=21
    1, 7, -4, -8, -2, 3, 0, -10, -9,
    -- layer=1 filter=12 channel=22
    2, -5, 7, 3, 3, 6, -6, 8, 3,
    -- layer=1 filter=12 channel=23
    8, -9, -5, 7, -6, -1, -10, -1, 4,
    -- layer=1 filter=12 channel=24
    -5, 1, -5, -5, -8, 0, -11, 4, 0,
    -- layer=1 filter=12 channel=25
    -3, 6, 4, 0, -1, 7, -4, 8, 4,
    -- layer=1 filter=12 channel=26
    0, -4, 5, 0, 1, 0, -6, -7, 9,
    -- layer=1 filter=12 channel=27
    0, -5, -6, -10, -4, 8, 0, 8, 0,
    -- layer=1 filter=12 channel=28
    -6, 2, -7, -9, 0, -12, -1, -2, 2,
    -- layer=1 filter=12 channel=29
    8, 9, 8, 7, 3, 4, -2, 6, -1,
    -- layer=1 filter=12 channel=30
    1, -4, -3, 5, 0, 9, -5, -10, -5,
    -- layer=1 filter=12 channel=31
    7, -7, -8, 1, -3, -2, -13, -11, 2,
    -- layer=1 filter=12 channel=32
    -7, -8, 5, -3, -7, -2, 0, 5, -10,
    -- layer=1 filter=12 channel=33
    5, 7, -6, 3, -9, -3, 3, -1, -8,
    -- layer=1 filter=12 channel=34
    3, 0, -4, -7, -7, 4, 6, -5, 1,
    -- layer=1 filter=12 channel=35
    0, -4, 8, 8, -2, -1, 8, -7, -9,
    -- layer=1 filter=12 channel=36
    3, -4, -5, 6, -6, -5, -5, -1, -3,
    -- layer=1 filter=12 channel=37
    -3, -3, -2, 6, -2, 5, 6, 9, 0,
    -- layer=1 filter=12 channel=38
    -5, -12, -11, -2, 0, -4, -8, 1, 8,
    -- layer=1 filter=12 channel=39
    -4, -11, 4, 7, 6, -6, -2, -11, -1,
    -- layer=1 filter=12 channel=40
    -1, -8, 0, -3, -4, -6, 7, -7, 2,
    -- layer=1 filter=12 channel=41
    -1, -10, 4, -11, -4, -3, -1, -11, -1,
    -- layer=1 filter=12 channel=42
    2, 5, 0, -4, -8, 5, -3, -7, 5,
    -- layer=1 filter=12 channel=43
    -11, 4, -3, 7, 3, 0, 1, 0, 0,
    -- layer=1 filter=12 channel=44
    2, -6, 5, 6, 0, -9, -1, -10, 6,
    -- layer=1 filter=12 channel=45
    5, 5, 1, 4, 8, -3, -7, -1, -5,
    -- layer=1 filter=12 channel=46
    -7, 0, -8, -3, 4, 7, 1, -1, -5,
    -- layer=1 filter=12 channel=47
    9, 7, -7, 9, -7, 6, -9, 2, 7,
    -- layer=1 filter=12 channel=48
    -7, -11, -2, 0, -7, -6, 0, -11, -3,
    -- layer=1 filter=12 channel=49
    -6, 6, -6, -5, -11, 4, -2, -5, -1,
    -- layer=1 filter=12 channel=50
    -1, -4, 8, -8, -9, -6, 0, -4, -8,
    -- layer=1 filter=12 channel=51
    -11, 1, 3, 0, -11, -3, -6, -11, -12,
    -- layer=1 filter=12 channel=52
    -9, -7, -4, 5, -6, 7, -7, 3, -3,
    -- layer=1 filter=12 channel=53
    -9, -5, -10, 0, -2, -9, 4, 7, 0,
    -- layer=1 filter=12 channel=54
    -5, 0, -6, 2, -1, 4, -2, -8, 0,
    -- layer=1 filter=12 channel=55
    8, 9, 2, 3, -10, -5, 9, 1, -6,
    -- layer=1 filter=12 channel=56
    -4, -3, 7, 1, 5, -7, -8, -1, 4,
    -- layer=1 filter=12 channel=57
    -3, 7, -2, -2, -11, -1, 1, 5, 1,
    -- layer=1 filter=12 channel=58
    -3, -9, 5, 6, -4, -9, -6, 8, -3,
    -- layer=1 filter=12 channel=59
    -1, 0, -8, 8, 0, -2, -1, -8, 8,
    -- layer=1 filter=12 channel=60
    9, -6, 10, -6, 0, 4, -4, -3, -7,
    -- layer=1 filter=12 channel=61
    -7, 5, -8, -5, -7, -7, -6, -3, -5,
    -- layer=1 filter=12 channel=62
    -9, 1, 9, 1, -8, -2, -7, 10, -7,
    -- layer=1 filter=12 channel=63
    -11, 3, -9, 0, -1, -11, 5, -5, 7,
    -- layer=1 filter=12 channel=64
    5, 4, -10, 7, 0, 3, 6, -6, -3,
    -- layer=1 filter=12 channel=65
    1, -8, 6, -11, -2, 8, 5, -8, -6,
    -- layer=1 filter=12 channel=66
    7, 2, -11, 2, 4, 0, 4, -9, 7,
    -- layer=1 filter=12 channel=67
    4, 4, 8, -1, 0, 4, 9, -1, -6,
    -- layer=1 filter=12 channel=68
    -4, 2, -8, -8, 6, 0, -10, -8, 7,
    -- layer=1 filter=12 channel=69
    6, -10, 5, -6, 3, 9, 0, 1, 0,
    -- layer=1 filter=12 channel=70
    -3, 8, 8, -4, -3, -7, -1, 0, 0,
    -- layer=1 filter=12 channel=71
    -4, 5, -8, -4, -5, -11, -6, -5, -2,
    -- layer=1 filter=12 channel=72
    6, 1, -2, -5, 3, -5, 1, 2, -5,
    -- layer=1 filter=12 channel=73
    -7, 3, 1, 0, 7, -5, 1, 5, 9,
    -- layer=1 filter=12 channel=74
    1, 8, 6, 0, 0, -12, -4, -2, -10,
    -- layer=1 filter=12 channel=75
    -4, 0, 1, 3, -8, 0, -9, -9, 5,
    -- layer=1 filter=12 channel=76
    6, 0, 6, -10, 1, 3, -6, 0, 5,
    -- layer=1 filter=12 channel=77
    -10, -5, -1, -3, 2, 6, -4, 3, 2,
    -- layer=1 filter=12 channel=78
    5, 7, 0, -7, -10, 7, -7, -5, -8,
    -- layer=1 filter=12 channel=79
    5, -8, -5, -6, -9, -6, -4, -8, 0,
    -- layer=1 filter=12 channel=80
    7, -3, 0, -6, -2, 0, -6, -1, 9,
    -- layer=1 filter=12 channel=81
    4, 0, 8, 6, 0, -7, -6, -6, -8,
    -- layer=1 filter=12 channel=82
    -8, 4, 7, 7, -6, -11, 6, -4, 7,
    -- layer=1 filter=12 channel=83
    1, 0, -5, 0, -8, 0, -8, 6, 1,
    -- layer=1 filter=12 channel=84
    -1, -11, 3, -2, 4, 0, -3, -3, -2,
    -- layer=1 filter=12 channel=85
    -11, -10, 0, 5, -4, 6, 1, 7, 7,
    -- layer=1 filter=12 channel=86
    -5, -3, -10, -3, -10, -3, 8, 7, -11,
    -- layer=1 filter=12 channel=87
    5, -1, -2, -5, -10, -9, 2, 0, -8,
    -- layer=1 filter=12 channel=88
    2, -12, -12, 0, -7, 1, 0, -9, 1,
    -- layer=1 filter=12 channel=89
    6, -7, -2, -11, 7, -6, -6, -2, 0,
    -- layer=1 filter=12 channel=90
    -4, 0, 1, 7, 1, 7, -11, 6, -3,
    -- layer=1 filter=12 channel=91
    -4, -2, 8, 3, 0, 6, -10, 0, 3,
    -- layer=1 filter=12 channel=92
    -8, 8, -1, -4, 3, -4, -9, 1, -4,
    -- layer=1 filter=12 channel=93
    -2, -5, 0, 6, -1, 5, 6, -4, -11,
    -- layer=1 filter=12 channel=94
    -3, -12, -4, 5, -11, 0, 8, -4, 0,
    -- layer=1 filter=12 channel=95
    0, -9, -8, -4, -4, -9, -4, -6, -8,
    -- layer=1 filter=12 channel=96
    1, 3, -10, 8, 8, -12, -1, -12, 0,
    -- layer=1 filter=12 channel=97
    0, -6, -12, -5, -8, 3, 7, -8, 3,
    -- layer=1 filter=12 channel=98
    9, -9, 4, 0, 2, 4, 7, 5, -9,
    -- layer=1 filter=12 channel=99
    -11, -12, -3, -1, -8, -7, 5, -3, 1,
    -- layer=1 filter=12 channel=100
    3, -10, -9, -3, -2, 3, -1, 0, 1,
    -- layer=1 filter=12 channel=101
    3, -1, 8, -5, -8, -4, 7, -7, -8,
    -- layer=1 filter=12 channel=102
    -8, -2, -3, -9, -10, 6, -10, 4, 5,
    -- layer=1 filter=12 channel=103
    4, -2, 5, -7, 0, 1, -7, 1, 9,
    -- layer=1 filter=12 channel=104
    -8, -11, 2, -5, 5, 5, -2, 0, 3,
    -- layer=1 filter=12 channel=105
    5, -1, -11, -9, -8, 1, -8, 4, -5,
    -- layer=1 filter=12 channel=106
    6, -7, 0, -12, 0, -10, -6, 1, -4,
    -- layer=1 filter=12 channel=107
    0, -4, 11, 8, 5, 4, 9, -1, 9,
    -- layer=1 filter=12 channel=108
    -2, -7, -7, -7, -9, -10, -7, 3, 2,
    -- layer=1 filter=12 channel=109
    -5, 7, -3, 10, 6, 1, 9, 3, -6,
    -- layer=1 filter=12 channel=110
    -1, 0, 6, 0, 9, 0, -3, 1, 7,
    -- layer=1 filter=12 channel=111
    0, 6, -2, 5, 7, 2, 1, -7, -1,
    -- layer=1 filter=12 channel=112
    0, -1, 4, 1, 0, 5, -8, -2, -1,
    -- layer=1 filter=12 channel=113
    -7, -2, 3, 6, -7, -6, 3, -10, 6,
    -- layer=1 filter=12 channel=114
    1, 8, 5, 5, -8, 4, 4, -4, -4,
    -- layer=1 filter=12 channel=115
    -10, -8, 7, -10, 2, -10, 3, 8, -4,
    -- layer=1 filter=12 channel=116
    -5, -5, -3, 0, -5, -9, 8, 1, -5,
    -- layer=1 filter=12 channel=117
    -1, -2, 7, 0, -4, -7, -5, -1, -2,
    -- layer=1 filter=12 channel=118
    4, -6, 0, 2, -6, -9, 7, -6, 0,
    -- layer=1 filter=12 channel=119
    -13, -7, -1, 6, -9, -2, 5, 5, -7,
    -- layer=1 filter=12 channel=120
    -3, 6, -6, -4, 6, -2, 10, 2, -3,
    -- layer=1 filter=12 channel=121
    -7, -1, -6, -5, 0, 0, -2, 0, -9,
    -- layer=1 filter=12 channel=122
    -3, 10, -6, -8, 10, 1, -7, 5, 4,
    -- layer=1 filter=12 channel=123
    3, -12, -7, -11, 3, -1, 4, -9, -1,
    -- layer=1 filter=12 channel=124
    -2, 9, -1, 4, 3, -4, 0, 0, -9,
    -- layer=1 filter=12 channel=125
    8, -5, 8, -2, 8, 4, 5, -11, -1,
    -- layer=1 filter=12 channel=126
    4, 5, -7, -5, 2, 0, -6, -3, 0,
    -- layer=1 filter=12 channel=127
    8, -2, 0, 0, 7, -8, 0, 0, -2,
    -- layer=1 filter=13 channel=0
    -10, 4, -11, -4, -1, 6, -3, -11, 4,
    -- layer=1 filter=13 channel=1
    5, -9, 5, -1, -4, 7, -10, -11, 0,
    -- layer=1 filter=13 channel=2
    -3, -4, -2, 2, 1, 1, 4, -8, -9,
    -- layer=1 filter=13 channel=3
    -11, 5, -9, 4, -6, 4, 5, 5, -5,
    -- layer=1 filter=13 channel=4
    -3, -5, 0, 4, 6, 0, -6, 0, -2,
    -- layer=1 filter=13 channel=5
    -4, 11, -7, -7, 0, 0, 8, -4, 4,
    -- layer=1 filter=13 channel=6
    1, -5, -7, -3, -9, -10, -11, 4, 6,
    -- layer=1 filter=13 channel=7
    -2, -14, 3, -10, 9, -1, -5, -4, -3,
    -- layer=1 filter=13 channel=8
    -10, 0, 0, -3, 0, -15, 7, -10, -4,
    -- layer=1 filter=13 channel=9
    0, 2, 6, 5, -2, -5, 3, -3, 9,
    -- layer=1 filter=13 channel=10
    4, -14, 1, 0, 3, -7, -8, -9, -5,
    -- layer=1 filter=13 channel=11
    6, -6, -4, -3, 9, 6, -1, -15, -4,
    -- layer=1 filter=13 channel=12
    7, 1, -13, 2, 5, -1, 0, 0, 1,
    -- layer=1 filter=13 channel=13
    -12, 7, -11, -11, -10, -8, -3, 2, 3,
    -- layer=1 filter=13 channel=14
    -2, -3, -3, 3, 2, 0, -5, 6, -16,
    -- layer=1 filter=13 channel=15
    2, -11, -6, 1, -6, -1, -4, -6, 2,
    -- layer=1 filter=13 channel=16
    -8, -9, -7, -5, -5, -4, 1, 7, -3,
    -- layer=1 filter=13 channel=17
    -3, -4, -9, 0, 6, -6, -11, 4, -7,
    -- layer=1 filter=13 channel=18
    -4, -2, -1, 4, 4, -8, -10, -6, 5,
    -- layer=1 filter=13 channel=19
    -11, -3, 3, 0, -4, 2, 2, -11, 4,
    -- layer=1 filter=13 channel=20
    -12, 0, -1, -1, 6, -1, -11, -11, -6,
    -- layer=1 filter=13 channel=21
    3, -3, -2, 4, -7, 0, 8, -10, -11,
    -- layer=1 filter=13 channel=22
    -6, 1, -1, -13, 3, -5, -5, 6, 0,
    -- layer=1 filter=13 channel=23
    0, -8, -5, -6, -5, -12, -9, 6, -6,
    -- layer=1 filter=13 channel=24
    -6, -13, -16, -11, -7, -8, 1, 0, -7,
    -- layer=1 filter=13 channel=25
    -6, -4, -1, -11, 7, -16, -9, -2, -9,
    -- layer=1 filter=13 channel=26
    -4, -1, -14, -15, -2, -14, -5, -14, -5,
    -- layer=1 filter=13 channel=27
    -7, -8, 6, 2, -1, -8, -9, -3, 3,
    -- layer=1 filter=13 channel=28
    -2, 6, -10, -12, 4, -2, -3, -4, -3,
    -- layer=1 filter=13 channel=29
    -2, 0, 5, -9, -5, -9, -10, -2, 1,
    -- layer=1 filter=13 channel=30
    -1, 0, 0, 5, -1, 8, 0, -12, -5,
    -- layer=1 filter=13 channel=31
    -5, -6, -11, -2, -2, 1, 0, -11, -13,
    -- layer=1 filter=13 channel=32
    -9, -9, -11, -12, -3, 5, -6, -1, -1,
    -- layer=1 filter=13 channel=33
    -7, 6, -1, 5, 10, 0, 6, -4, -2,
    -- layer=1 filter=13 channel=34
    1, 3, -4, -8, 5, -10, -5, 3, 6,
    -- layer=1 filter=13 channel=35
    7, 1, -5, -3, 1, -2, -12, -9, -12,
    -- layer=1 filter=13 channel=36
    -3, -5, 6, 2, -1, 4, -6, -7, 6,
    -- layer=1 filter=13 channel=37
    -6, -2, 3, -13, -4, 0, -3, 3, -7,
    -- layer=1 filter=13 channel=38
    -12, 3, -14, 0, 1, -9, 2, 2, 5,
    -- layer=1 filter=13 channel=39
    5, -8, -4, -7, -3, 6, -2, 0, 0,
    -- layer=1 filter=13 channel=40
    -2, 1, -12, -5, -5, -11, -15, -14, 1,
    -- layer=1 filter=13 channel=41
    -10, -3, 5, -10, 6, 5, -9, -12, 6,
    -- layer=1 filter=13 channel=42
    1, -2, 1, 4, -7, 0, 8, 7, -3,
    -- layer=1 filter=13 channel=43
    -7, 3, 1, -16, -9, -13, 6, -11, -11,
    -- layer=1 filter=13 channel=44
    0, 6, -7, 6, -8, 2, -9, -11, -4,
    -- layer=1 filter=13 channel=45
    5, 4, 8, 1, -13, -8, -8, -12, -5,
    -- layer=1 filter=13 channel=46
    -12, 0, -10, -18, -13, -6, 5, 13, 11,
    -- layer=1 filter=13 channel=47
    1, -1, -8, -5, 2, -16, -5, -2, -16,
    -- layer=1 filter=13 channel=48
    6, -8, 1, 1, 8, 6, 7, -9, 7,
    -- layer=1 filter=13 channel=49
    -5, 3, -7, -5, 6, -10, 0, -9, -1,
    -- layer=1 filter=13 channel=50
    -9, -1, -5, 0, -3, 5, -4, 6, -11,
    -- layer=1 filter=13 channel=51
    2, 7, 3, -10, -12, -11, 1, -4, -14,
    -- layer=1 filter=13 channel=52
    -7, 7, -4, -4, 1, 4, 0, 0, 9,
    -- layer=1 filter=13 channel=53
    0, -5, 7, 2, -9, 7, -4, -5, -11,
    -- layer=1 filter=13 channel=54
    3, -11, -16, -8, -9, -13, -3, -5, -2,
    -- layer=1 filter=13 channel=55
    -10, 4, -1, 4, 1, -7, -15, 2, -12,
    -- layer=1 filter=13 channel=56
    4, 2, 4, 4, -4, 1, 4, -6, -5,
    -- layer=1 filter=13 channel=57
    2, -13, -12, -2, -10, -10, -9, -8, 1,
    -- layer=1 filter=13 channel=58
    -1, 2, 1, 7, -4, 1, -3, 3, -11,
    -- layer=1 filter=13 channel=59
    2, 8, 3, -3, 3, -5, -11, 5, -7,
    -- layer=1 filter=13 channel=60
    -1, -7, 1, -2, 8, -11, 11, -5, -2,
    -- layer=1 filter=13 channel=61
    -6, 1, -1, 7, 7, 0, 1, 7, 0,
    -- layer=1 filter=13 channel=62
    -7, 1, -5, 1, -4, -4, -8, -6, 2,
    -- layer=1 filter=13 channel=63
    6, 0, 0, -4, 0, -11, -13, -4, 3,
    -- layer=1 filter=13 channel=64
    -10, -9, 0, 1, -6, 2, 8, 0, 1,
    -- layer=1 filter=13 channel=65
    2, 3, 5, -10, -10, -2, -4, -1, -9,
    -- layer=1 filter=13 channel=66
    -5, -10, -10, -12, -9, -1, -11, -5, 2,
    -- layer=1 filter=13 channel=67
    7, 2, 5, -1, -8, 0, -6, 8, 8,
    -- layer=1 filter=13 channel=68
    0, 6, -2, 8, 2, -4, 0, -12, -5,
    -- layer=1 filter=13 channel=69
    -9, -4, 1, -13, -15, -14, 0, 8, 6,
    -- layer=1 filter=13 channel=70
    0, -5, -9, -8, 1, -1, 1, -8, 0,
    -- layer=1 filter=13 channel=71
    -7, -6, -12, -1, -8, -3, -5, 6, -3,
    -- layer=1 filter=13 channel=72
    0, -3, -4, -2, -7, -11, -8, -15, 0,
    -- layer=1 filter=13 channel=73
    1, -5, 5, 1, -10, -8, -9, -8, -2,
    -- layer=1 filter=13 channel=74
    0, -12, 6, 0, -8, 1, 4, 0, -9,
    -- layer=1 filter=13 channel=75
    -6, 4, 0, 0, 9, 0, -6, 8, 0,
    -- layer=1 filter=13 channel=76
    -9, 6, -9, 1, 0, -6, -7, 1, -11,
    -- layer=1 filter=13 channel=77
    -6, 0, 3, -7, 0, -8, -4, -1, -4,
    -- layer=1 filter=13 channel=78
    0, -2, -8, -2, 0, -6, 4, 6, 4,
    -- layer=1 filter=13 channel=79
    -9, -3, -4, -3, 0, -3, -4, -10, -10,
    -- layer=1 filter=13 channel=80
    2, 5, -8, -3, -7, 4, 0, 1, 9,
    -- layer=1 filter=13 channel=81
    -12, 0, -11, 0, -12, 2, -2, -6, -4,
    -- layer=1 filter=13 channel=82
    -4, 0, -9, -9, 2, -12, 0, 0, 0,
    -- layer=1 filter=13 channel=83
    0, 6, 5, 4, -2, 2, -9, 6, 7,
    -- layer=1 filter=13 channel=84
    8, -9, -5, 11, 8, 7, 2, 0, 3,
    -- layer=1 filter=13 channel=85
    7, -3, 3, -6, 5, -11, -11, -11, -6,
    -- layer=1 filter=13 channel=86
    -6, -3, -11, 0, -6, -10, 1, -11, -1,
    -- layer=1 filter=13 channel=87
    -10, 4, 0, 1, -4, 3, -2, -3, -3,
    -- layer=1 filter=13 channel=88
    4, -10, -10, 1, 0, -7, -8, -9, -12,
    -- layer=1 filter=13 channel=89
    -10, -9, 8, 0, -3, -7, -5, -5, 4,
    -- layer=1 filter=13 channel=90
    -6, 7, -8, -9, -12, -9, -10, 3, -7,
    -- layer=1 filter=13 channel=91
    -5, -14, -8, -3, -1, -10, 0, -11, -11,
    -- layer=1 filter=13 channel=92
    6, -9, 7, -2, -18, 8, -2, 5, 1,
    -- layer=1 filter=13 channel=93
    -12, 0, -4, -4, -13, -10, -9, -10, 4,
    -- layer=1 filter=13 channel=94
    -5, -2, -4, -3, 7, -3, 2, 2, 2,
    -- layer=1 filter=13 channel=95
    0, -5, 0, -8, -1, -10, -3, -7, -2,
    -- layer=1 filter=13 channel=96
    4, 8, -11, -3, -10, 1, 3, 7, 6,
    -- layer=1 filter=13 channel=97
    -1, -13, -4, 4, 5, 6, -9, 2, -10,
    -- layer=1 filter=13 channel=98
    4, -11, -10, -9, -3, -4, -5, -2, -7,
    -- layer=1 filter=13 channel=99
    0, 4, 4, -5, -1, 0, -13, 1, -10,
    -- layer=1 filter=13 channel=100
    -11, 2, 7, 2, -10, -13, 0, 4, -11,
    -- layer=1 filter=13 channel=101
    -7, 0, 3, -6, 7, -4, -4, 0, -2,
    -- layer=1 filter=13 channel=102
    -12, -9, -1, 2, -4, 0, -11, 0, 2,
    -- layer=1 filter=13 channel=103
    -7, 4, -3, -1, 6, 2, 3, -4, 4,
    -- layer=1 filter=13 channel=104
    7, -2, 5, 6, -7, 2, -8, -9, -10,
    -- layer=1 filter=13 channel=105
    -12, -5, -4, -2, -6, -9, 2, -8, 2,
    -- layer=1 filter=13 channel=106
    -10, -8, -14, -11, 1, -10, -8, 2, -13,
    -- layer=1 filter=13 channel=107
    5, 4, 2, -12, -2, 5, 7, 3, 5,
    -- layer=1 filter=13 channel=108
    5, -6, 6, -7, 2, -13, 2, 0, 7,
    -- layer=1 filter=13 channel=109
    3, 3, 10, 7, 1, 5, -3, -8, 5,
    -- layer=1 filter=13 channel=110
    -9, -5, -12, 7, 5, 6, 5, -6, -4,
    -- layer=1 filter=13 channel=111
    6, 1, -5, -10, -4, 2, -3, -15, -5,
    -- layer=1 filter=13 channel=112
    -12, 2, 3, 1, 2, 2, -13, 3, 0,
    -- layer=1 filter=13 channel=113
    -4, -11, -12, -2, -4, -1, -3, -5, -14,
    -- layer=1 filter=13 channel=114
    -4, 8, 2, -9, -7, 3, -2, -4, 5,
    -- layer=1 filter=13 channel=115
    -9, 6, -3, 3, -9, 0, 2, 6, -2,
    -- layer=1 filter=13 channel=116
    5, -8, -7, -2, -9, -3, -8, 3, -8,
    -- layer=1 filter=13 channel=117
    -1, 2, 9, -9, 6, -8, -19, -10, 3,
    -- layer=1 filter=13 channel=118
    7, 5, 6, -8, -11, -10, 1, -3, -3,
    -- layer=1 filter=13 channel=119
    -10, -10, -6, 10, 0, 7, 4, -8, -2,
    -- layer=1 filter=13 channel=120
    3, -3, 2, -8, 5, -3, -10, -6, -7,
    -- layer=1 filter=13 channel=121
    -11, -7, -11, 0, 4, -7, -4, -7, -6,
    -- layer=1 filter=13 channel=122
    6, 1, 4, 9, 5, 0, 3, -7, -9,
    -- layer=1 filter=13 channel=123
    -4, -4, 2, -5, -5, 0, 2, -4, -13,
    -- layer=1 filter=13 channel=124
    -9, -4, -10, 0, 0, 4, 6, 7, -10,
    -- layer=1 filter=13 channel=125
    -8, 2, -16, -1, -6, -1, 7, -2, -10,
    -- layer=1 filter=13 channel=126
    3, 4, -10, -2, 6, -9, -11, -8, 3,
    -- layer=1 filter=13 channel=127
    0, -11, -7, 2, 0, 2, 2, -3, -5,
    -- layer=1 filter=14 channel=0
    7, 11, 5, 3, -7, -17, -13, -12, 3,
    -- layer=1 filter=14 channel=1
    13, -25, -36, -12, 11, 17, 13, 21, 12,
    -- layer=1 filter=14 channel=2
    -1, -23, -8, -10, -2, -1, -1, 2, -11,
    -- layer=1 filter=14 channel=3
    10, -11, 15, -2, -13, -5, 7, 1, -8,
    -- layer=1 filter=14 channel=4
    -13, -4, -3, -13, -12, -6, 5, -11, -2,
    -- layer=1 filter=14 channel=5
    -2, -82, -57, 22, 41, 22, 23, 13, 4,
    -- layer=1 filter=14 channel=6
    22, 30, 36, -30, -42, -34, -75, -66, -34,
    -- layer=1 filter=14 channel=7
    40, 6, -7, -25, -19, 13, -25, -31, -33,
    -- layer=1 filter=14 channel=8
    -22, -76, -87, 14, 33, 40, 38, 46, 12,
    -- layer=1 filter=14 channel=9
    -21, 6, 16, 2, -36, -26, -32, -27, -78,
    -- layer=1 filter=14 channel=10
    39, 33, 18, -24, -3, 4, -24, -58, -49,
    -- layer=1 filter=14 channel=11
    -9, 20, 13, -11, 10, 0, -18, -13, 1,
    -- layer=1 filter=14 channel=12
    -19, 0, -13, 11, 16, -14, -4, 6, -15,
    -- layer=1 filter=14 channel=13
    -8, 16, 4, 9, -5, -8, 4, 15, 4,
    -- layer=1 filter=14 channel=14
    36, 17, 11, 25, 36, 7, 13, -11, -54,
    -- layer=1 filter=14 channel=15
    4, -25, -35, 10, 30, 2, 28, 9, 3,
    -- layer=1 filter=14 channel=16
    -26, -75, -73, 12, 43, 41, 26, 47, 20,
    -- layer=1 filter=14 channel=17
    -19, 0, -13, -10, -4, -3, 9, 23, 3,
    -- layer=1 filter=14 channel=18
    0, 22, 13, 20, 21, 12, -14, -44, -49,
    -- layer=1 filter=14 channel=19
    7, 7, 12, 61, 56, 58, 21, 5, -36,
    -- layer=1 filter=14 channel=20
    -5, -19, -12, -8, -19, 0, 16, 23, 16,
    -- layer=1 filter=14 channel=21
    19, 5, 2, -28, -7, -11, 0, 0, 6,
    -- layer=1 filter=14 channel=22
    -13, -17, -29, -17, -14, 5, 28, 34, 32,
    -- layer=1 filter=14 channel=23
    23, -5, 48, 3, -5, 22, -32, -16, -34,
    -- layer=1 filter=14 channel=24
    -31, 2, 4, 13, -2, 11, 12, 10, 1,
    -- layer=1 filter=14 channel=25
    40, -16, -6, -17, 18, 25, 13, 17, -23,
    -- layer=1 filter=14 channel=26
    -24, 5, 8, 35, 20, 1, -8, 10, 1,
    -- layer=1 filter=14 channel=27
    -10, -12, -3, -30, -18, 0, -17, -5, -12,
    -- layer=1 filter=14 channel=28
    40, 15, -6, -22, 0, 8, 0, 3, -11,
    -- layer=1 filter=14 channel=29
    -3, -35, -11, -35, -33, -34, -13, -11, -4,
    -- layer=1 filter=14 channel=30
    5, 17, 18, 22, 34, 5, -13, -34, -55,
    -- layer=1 filter=14 channel=31
    0, 0, -9, 2, 1, -2, -43, -55, -72,
    -- layer=1 filter=14 channel=32
    14, 28, 47, 16, 22, -2, -63, -65, -44,
    -- layer=1 filter=14 channel=33
    18, 16, -3, 3, -4, -14, -21, -18, -11,
    -- layer=1 filter=14 channel=34
    18, 33, 22, 38, 13, 0, -21, -29, -27,
    -- layer=1 filter=14 channel=35
    8, -16, -21, 12, -10, -17, -5, -6, 5,
    -- layer=1 filter=14 channel=36
    -4, -1, 18, -8, -6, 5, -5, -5, -18,
    -- layer=1 filter=14 channel=37
    -15, -62, -29, 21, 34, 22, 24, 15, -16,
    -- layer=1 filter=14 channel=38
    6, 22, 12, -25, -15, -10, -9, -16, -8,
    -- layer=1 filter=14 channel=39
    -21, -17, -10, -15, -6, 9, 9, 9, 7,
    -- layer=1 filter=14 channel=40
    7, 19, 6, -19, -21, -18, -43, -63, -52,
    -- layer=1 filter=14 channel=41
    -11, 29, 56, 21, 17, -11, -64, -49, -68,
    -- layer=1 filter=14 channel=42
    -26, -23, -18, 6, -17, 3, 4, -4, -9,
    -- layer=1 filter=14 channel=43
    -20, -67, -72, 0, 13, 29, 24, 21, 7,
    -- layer=1 filter=14 channel=44
    1, 43, 17, -6, 5, -32, -53, -35, -15,
    -- layer=1 filter=14 channel=45
    -11, -6, -6, 2, -6, -16, -1, 18, 10,
    -- layer=1 filter=14 channel=46
    51, 2, -44, 44, 25, 6, 13, 2, 3,
    -- layer=1 filter=14 channel=47
    38, -5, 60, 9, -6, -14, -70, -66, -98,
    -- layer=1 filter=14 channel=48
    2, 22, 15, -12, -26, -22, -7, -7, 5,
    -- layer=1 filter=14 channel=49
    8, 4, 19, 1, -3, -13, -23, -27, -27,
    -- layer=1 filter=14 channel=50
    -16, -13, 7, -13, -30, -11, -34, -31, -22,
    -- layer=1 filter=14 channel=51
    28, 32, 5, -19, -30, -4, -4, -12, -13,
    -- layer=1 filter=14 channel=52
    8, 12, -2, 3, -3, 11, 1, 2, 2,
    -- layer=1 filter=14 channel=53
    -4, 22, -19, -2, 13, 4, 16, 3, 9,
    -- layer=1 filter=14 channel=54
    14, -8, -4, 12, 22, 32, 16, 2, -40,
    -- layer=1 filter=14 channel=55
    -3, -11, -6, 2, 8, -2, -6, 6, 10,
    -- layer=1 filter=14 channel=56
    0, -1, 7, -2, 0, -2, 0, 0, -10,
    -- layer=1 filter=14 channel=57
    22, 9, 0, -22, -17, 2, -19, -42, -50,
    -- layer=1 filter=14 channel=58
    57, -7, 59, -28, -10, 5, -43, -53, -77,
    -- layer=1 filter=14 channel=59
    -10, 0, -10, -9, -3, -7, 17, 1, 0,
    -- layer=1 filter=14 channel=60
    10, 8, 1, 14, 7, 0, -6, -3, 0,
    -- layer=1 filter=14 channel=61
    -8, -3, 0, -2, -9, -2, 3, -7, -21,
    -- layer=1 filter=14 channel=62
    -13, -69, -54, 32, 39, 52, 44, 35, 0,
    -- layer=1 filter=14 channel=63
    -2, 28, 22, 8, -5, -10, -29, -39, -20,
    -- layer=1 filter=14 channel=64
    19, -3, 14, 8, -9, 5, -3, 1, 4,
    -- layer=1 filter=14 channel=65
    -3, 1, 4, -23, -7, -9, 0, 3, 18,
    -- layer=1 filter=14 channel=66
    10, 5, 13, -4, -14, 0, -3, 2, -13,
    -- layer=1 filter=14 channel=67
    9, 12, 25, -38, -28, -19, -56, -45, -54,
    -- layer=1 filter=14 channel=68
    0, 58, 27, -2, 9, -38, -66, -58, -29,
    -- layer=1 filter=14 channel=69
    -42, -69, -53, 15, 34, 18, 33, 38, -5,
    -- layer=1 filter=14 channel=70
    52, 51, 17, 7, 29, 27, 0, -47, -66,
    -- layer=1 filter=14 channel=71
    3, -14, -23, -9, 10, 0, 8, 8, 8,
    -- layer=1 filter=14 channel=72
    -2, 0, 6, 24, 7, 18, -12, -23, -16,
    -- layer=1 filter=14 channel=73
    -5, 6, 5, -18, -12, 2, -13, 1, -15,
    -- layer=1 filter=14 channel=74
    5, 32, 6, -5, 32, -5, -62, -86, -64,
    -- layer=1 filter=14 channel=75
    3, -17, -28, 6, 5, -3, -18, -30, -35,
    -- layer=1 filter=14 channel=76
    3, 22, 35, -6, 16, -23, -31, -34, -21,
    -- layer=1 filter=14 channel=77
    -10, 10, -9, -21, -14, -17, -13, -9, 0,
    -- layer=1 filter=14 channel=78
    11, 0, 7, -16, -22, -13, 9, -20, -27,
    -- layer=1 filter=14 channel=79
    -36, -80, -58, 11, 22, 39, 39, 29, 5,
    -- layer=1 filter=14 channel=80
    5, 15, -3, -12, 13, -5, 3, 4, 15,
    -- layer=1 filter=14 channel=81
    -23, -19, -28, -6, -6, -6, 10, 18, 13,
    -- layer=1 filter=14 channel=82
    26, 12, 26, 0, -29, -22, -9, -4, 9,
    -- layer=1 filter=14 channel=83
    -9, 7, -11, 20, 11, -3, -5, 21, -1,
    -- layer=1 filter=14 channel=84
    6, 30, 44, 24, 48, 1, -32, -45, -24,
    -- layer=1 filter=14 channel=85
    34, 29, 53, 51, -2, 23, -49, -41, -75,
    -- layer=1 filter=14 channel=86
    -14, -18, -3, -4, 17, 13, 6, 0, 17,
    -- layer=1 filter=14 channel=87
    -1, -1, -11, 24, -5, 4, -23, -35, -39,
    -- layer=1 filter=14 channel=88
    3, 0, 9, 2, -17, 0, 7, 6, 2,
    -- layer=1 filter=14 channel=89
    16, 30, 14, -12, -30, -21, -14, -15, -4,
    -- layer=1 filter=14 channel=90
    -16, 16, 2, 8, 20, -5, -7, 0, -2,
    -- layer=1 filter=14 channel=91
    30, 26, 12, 0, -20, -9, -5, -22, -12,
    -- layer=1 filter=14 channel=92
    -53, 21, -25, -8, -23, -29, -34, -66, -45,
    -- layer=1 filter=14 channel=93
    8, 13, 9, -14, -3, 2, 16, 16, 3,
    -- layer=1 filter=14 channel=94
    -2, 5, 0, -8, -15, -3, 4, -8, 4,
    -- layer=1 filter=14 channel=95
    33, 25, 29, 26, 47, 22, -41, -31, -54,
    -- layer=1 filter=14 channel=96
    -2, 4, -10, -6, -8, -15, -41, -30, -13,
    -- layer=1 filter=14 channel=97
    -1, 2, -2, -6, -8, -6, 15, 13, 10,
    -- layer=1 filter=14 channel=98
    -23, -39, -49, 4, -2, 24, 28, 32, 17,
    -- layer=1 filter=14 channel=99
    51, 90, 48, -9, 5, -5, -56, -67, -43,
    -- layer=1 filter=14 channel=100
    2, 28, 20, 2, 18, -5, -28, -29, -9,
    -- layer=1 filter=14 channel=101
    36, 37, 21, -7, -23, -26, -12, -21, 6,
    -- layer=1 filter=14 channel=102
    10, 28, 10, -12, -22, -18, -2, -17, -1,
    -- layer=1 filter=14 channel=103
    -4, 10, 19, 3, 0, 9, 6, -11, -13,
    -- layer=1 filter=14 channel=104
    32, 4, 29, 28, 12, 19, -34, -36, -34,
    -- layer=1 filter=14 channel=105
    12, 9, -1, -7, -14, -8, 3, -11, 5,
    -- layer=1 filter=14 channel=106
    17, 28, 27, -3, -15, -31, -38, -36, -19,
    -- layer=1 filter=14 channel=107
    -9, -19, -20, -5, -16, -12, -9, 1, -17,
    -- layer=1 filter=14 channel=108
    3, 21, 24, 17, 5, -18, -17, -13, -12,
    -- layer=1 filter=14 channel=109
    -8, -3, 3, 9, -6, -6, 3, 8, 6,
    -- layer=1 filter=14 channel=110
    4, 14, -3, 6, -18, -8, -3, 6, -8,
    -- layer=1 filter=14 channel=111
    16, 27, 27, 21, 39, 2, 1, -51, -36,
    -- layer=1 filter=14 channel=112
    21, 19, 23, 29, 30, 7, -35, -17, -11,
    -- layer=1 filter=14 channel=113
    25, 14, -4, 10, -14, -3, 5, -28, -26,
    -- layer=1 filter=14 channel=114
    -9, -56, -45, 10, 31, 27, 14, 22, 17,
    -- layer=1 filter=14 channel=115
    -5, -10, -4, -29, -8, 1, 1, -1, -2,
    -- layer=1 filter=14 channel=116
    7, 3, 4, 0, 1, 8, -10, 10, 0,
    -- layer=1 filter=14 channel=117
    45, 53, 21, 68, 50, 40, 15, 16, 9,
    -- layer=1 filter=14 channel=118
    3, 20, 13, -1, 19, 0, -52, -58, -68,
    -- layer=1 filter=14 channel=119
    -17, 40, 40, 26, 22, -18, -42, -37, -68,
    -- layer=1 filter=14 channel=120
    14, 10, 3, -19, -9, -6, 23, 12, 2,
    -- layer=1 filter=14 channel=121
    13, 15, 0, 24, 23, 21, -4, 4, -42,
    -- layer=1 filter=14 channel=122
    -1, -9, -8, 5, 8, 0, 2, -7, 8,
    -- layer=1 filter=14 channel=123
    6, -11, -18, 6, 21, 19, -24, -11, -32,
    -- layer=1 filter=14 channel=124
    1, -4, -19, -9, 0, 4, -3, 8, -12,
    -- layer=1 filter=14 channel=125
    57, 62, 52, 24, 23, 26, -24, -57, -53,
    -- layer=1 filter=14 channel=126
    -12, 34, -3, 25, 1, 24, 17, 27, -7,
    -- layer=1 filter=14 channel=127
    12, 16, 27, 27, 45, 17, -23, -31, -39,
    -- layer=1 filter=15 channel=0
    -15, -20, -7, -11, -11, 1, -6, -2, -1,
    -- layer=1 filter=15 channel=1
    4, -5, -10, 12, 11, -23, 2, -3, 11,
    -- layer=1 filter=15 channel=2
    8, 16, -2, 21, 0, 9, 5, 4, -16,
    -- layer=1 filter=15 channel=3
    -14, 4, -12, 1, -5, -11, -18, -5, 0,
    -- layer=1 filter=15 channel=4
    9, -1, 0, -2, -7, -6, 11, 6, 11,
    -- layer=1 filter=15 channel=5
    8, -18, -22, 15, 10, -34, -3, 8, 5,
    -- layer=1 filter=15 channel=6
    -21, -24, -33, -5, -23, -15, -35, -22, -31,
    -- layer=1 filter=15 channel=7
    32, 38, 41, 15, 56, 5, 12, 35, 22,
    -- layer=1 filter=15 channel=8
    11, -19, -16, -3, 0, -36, 3, -15, 9,
    -- layer=1 filter=15 channel=9
    -17, -23, 20, -11, -4, -60, 17, -45, -19,
    -- layer=1 filter=15 channel=10
    30, 27, 37, -1, 38, 14, 7, 22, 25,
    -- layer=1 filter=15 channel=11
    -36, -13, -14, -5, -12, 5, 13, 13, 6,
    -- layer=1 filter=15 channel=12
    1, -51, -17, -2, -49, -29, -11, 2, 34,
    -- layer=1 filter=15 channel=13
    -1, -11, 3, -1, -17, 15, -10, -9, 3,
    -- layer=1 filter=15 channel=14
    3, -3, 4, -16, -43, -8, -29, -11, -11,
    -- layer=1 filter=15 channel=15
    19, -15, -8, -13, -1, -15, 11, 7, 9,
    -- layer=1 filter=15 channel=16
    21, -11, -21, 18, 9, -26, 18, 0, 20,
    -- layer=1 filter=15 channel=17
    -6, 8, -7, -10, -1, 1, 1, -4, 3,
    -- layer=1 filter=15 channel=18
    -16, -14, -49, 16, -30, -25, -27, -34, -15,
    -- layer=1 filter=15 channel=19
    -20, -18, -8, 5, -5, -37, 21, 7, 47,
    -- layer=1 filter=15 channel=20
    -9, 4, 1, -7, 5, 6, 2, 7, 9,
    -- layer=1 filter=15 channel=21
    6, -11, -14, 0, 1, 0, -10, 1, -8,
    -- layer=1 filter=15 channel=22
    -2, -5, 2, -20, 10, -9, 8, 0, 4,
    -- layer=1 filter=15 channel=23
    31, 49, 38, 54, 78, 54, 36, 46, 72,
    -- layer=1 filter=15 channel=24
    6, -16, -14, 7, -26, -16, 1, -14, 5,
    -- layer=1 filter=15 channel=25
    26, 20, 15, -2, 33, -17, 15, 26, 25,
    -- layer=1 filter=15 channel=26
    -9, 0, 0, -3, -17, 16, -2, -26, 26,
    -- layer=1 filter=15 channel=27
    -54, -50, -15, -47, -41, -15, -24, -46, -19,
    -- layer=1 filter=15 channel=28
    10, 5, 14, -7, 24, 5, 7, 25, -6,
    -- layer=1 filter=15 channel=29
    13, 17, 39, 11, -5, 13, 5, -2, 8,
    -- layer=1 filter=15 channel=30
    -30, 10, -45, 4, -10, -25, -2, -43, -7,
    -- layer=1 filter=15 channel=31
    -19, -6, -2, 6, -25, 14, -25, 7, 0,
    -- layer=1 filter=15 channel=32
    -4, 40, 6, 7, 7, 33, -17, -17, 31,
    -- layer=1 filter=15 channel=33
    -1, -9, -17, 14, 7, -14, -3, -5, -17,
    -- layer=1 filter=15 channel=34
    -16, -44, -8, -54, 7, 10, -11, 9, -8,
    -- layer=1 filter=15 channel=35
    -11, -9, 4, 9, -2, -5, 7, -4, 1,
    -- layer=1 filter=15 channel=36
    -28, -10, -16, -19, -15, 8, 8, 16, 1,
    -- layer=1 filter=15 channel=37
    8, -5, -9, 17, -2, -35, 4, -4, 8,
    -- layer=1 filter=15 channel=38
    -2, 6, 12, 11, 9, 1, 9, 4, 6,
    -- layer=1 filter=15 channel=39
    3, -16, -3, -6, -12, -2, -1, -5, 0,
    -- layer=1 filter=15 channel=40
    2, 3, -3, 3, -7, -18, -10, -7, -31,
    -- layer=1 filter=15 channel=41
    -6, 54, 31, -9, 24, 17, -17, 8, 21,
    -- layer=1 filter=15 channel=42
    13, 41, -7, 5, 11, 35, 11, -8, 6,
    -- layer=1 filter=15 channel=43
    12, 9, -9, 9, 7, -21, -3, 2, 5,
    -- layer=1 filter=15 channel=44
    0, 11, 0, -6, -11, 17, 8, -20, 18,
    -- layer=1 filter=15 channel=45
    9, -14, -23, 11, -16, 7, 12, -11, 18,
    -- layer=1 filter=15 channel=46
    -17, -37, -76, -6, -34, -65, 9, -1, 8,
    -- layer=1 filter=15 channel=47
    33, 67, 34, 27, 56, 42, 0, 27, 45,
    -- layer=1 filter=15 channel=48
    -14, -5, -2, -2, 6, -12, -1, -11, -7,
    -- layer=1 filter=15 channel=49
    26, 4, -15, -3, -3, 0, -8, -1, -7,
    -- layer=1 filter=15 channel=50
    -11, -12, -10, -15, -16, -13, 0, -1, -10,
    -- layer=1 filter=15 channel=51
    4, -2, 19, -1, 2, -10, -4, 11, -16,
    -- layer=1 filter=15 channel=52
    7, 7, 6, 5, 11, -4, 5, 4, 12,
    -- layer=1 filter=15 channel=53
    -1, 17, 26, 7, 11, 11, 23, 3, 11,
    -- layer=1 filter=15 channel=54
    13, 34, 11, 17, 19, -18, 18, 16, 50,
    -- layer=1 filter=15 channel=55
    -2, 9, 12, -4, 3, 27, 5, 0, 13,
    -- layer=1 filter=15 channel=56
    7, -2, 11, 5, 8, 6, 7, 3, 5,
    -- layer=1 filter=15 channel=57
    18, 15, 15, -13, 8, -7, -2, 36, 2,
    -- layer=1 filter=15 channel=58
    37, 83, 53, 62, 97, 76, 21, 76, 85,
    -- layer=1 filter=15 channel=59
    5, 9, 9, -9, 0, 13, 5, -2, 0,
    -- layer=1 filter=15 channel=60
    -6, 2, 11, -16, -9, 4, 6, -1, -2,
    -- layer=1 filter=15 channel=61
    -8, -6, -10, -5, -10, 4, 0, -11, -7,
    -- layer=1 filter=15 channel=62
    1, -10, -8, 17, -7, -28, 11, -5, 8,
    -- layer=1 filter=15 channel=63
    -28, -22, -18, -16, -26, 7, -4, -2, 15,
    -- layer=1 filter=15 channel=64
    3, -10, 13, -6, -2, 7, 10, 10, -3,
    -- layer=1 filter=15 channel=65
    -10, -7, -2, -3, -12, 3, 8, 6, -17,
    -- layer=1 filter=15 channel=66
    -19, -8, -9, -10, 2, 9, -12, 7, 1,
    -- layer=1 filter=15 channel=67
    -6, -34, 3, -6, -26, -12, -6, -12, 29,
    -- layer=1 filter=15 channel=68
    18, 37, 15, 13, -1, 18, 17, 0, 32,
    -- layer=1 filter=15 channel=69
    19, -1, -9, 5, -9, -1, 15, 7, 17,
    -- layer=1 filter=15 channel=70
    -62, -74, -38, -50, -37, -18, -54, -31, -18,
    -- layer=1 filter=15 channel=71
    0, -1, -8, -5, -14, 0, 1, 8, -3,
    -- layer=1 filter=15 channel=72
    -42, -12, -50, 18, -18, -46, 19, -35, -3,
    -- layer=1 filter=15 channel=73
    5, -10, 0, -9, -7, 4, 3, 2, 12,
    -- layer=1 filter=15 channel=74
    -27, 2, 6, 32, 31, 9, 26, 15, 21,
    -- layer=1 filter=15 channel=75
    -39, -28, -37, 16, -38, -25, -35, -38, -13,
    -- layer=1 filter=15 channel=76
    -11, 21, -20, 0, -33, 4, 0, -16, 23,
    -- layer=1 filter=15 channel=77
    -14, -5, -6, 0, 0, -16, -4, -17, -11,
    -- layer=1 filter=15 channel=78
    -10, 1, 4, -14, 14, 5, 0, -3, -9,
    -- layer=1 filter=15 channel=79
    14, -6, -18, 11, 2, -18, 4, -10, 15,
    -- layer=1 filter=15 channel=80
    -7, 1, -7, -11, 1, 9, -3, 0, -7,
    -- layer=1 filter=15 channel=81
    -7, -19, -20, -12, -11, -2, -13, -17, -14,
    -- layer=1 filter=15 channel=82
    -5, -16, -3, 1, -15, 1, -2, -14, -10,
    -- layer=1 filter=15 channel=83
    -5, -7, -7, -8, -36, -15, -5, -3, 5,
    -- layer=1 filter=15 channel=84
    -5, 0, -17, 14, -26, 3, 0, -20, 18,
    -- layer=1 filter=15 channel=85
    9, 65, 26, 43, 60, 48, 12, 30, 67,
    -- layer=1 filter=15 channel=86
    -6, -5, 10, 3, 15, 7, 8, 12, 17,
    -- layer=1 filter=15 channel=87
    0, -4, 0, 16, -21, -31, 16, 4, 1,
    -- layer=1 filter=15 channel=88
    4, -7, -9, 3, -3, -3, 11, -1, -6,
    -- layer=1 filter=15 channel=89
    3, -9, -19, 0, -16, -6, -11, -12, 5,
    -- layer=1 filter=15 channel=90
    3, 0, 8, 1, 0, 13, 5, -5, 34,
    -- layer=1 filter=15 channel=91
    -2, 7, -3, -1, 2, -9, 2, 2, -7,
    -- layer=1 filter=15 channel=92
    5, -32, -29, -55, -26, -50, -34, -17, 0,
    -- layer=1 filter=15 channel=93
    -5, 0, 0, -5, 7, -2, -1, -2, 0,
    -- layer=1 filter=15 channel=94
    -6, -18, 6, -19, 1, -3, 0, 0, 2,
    -- layer=1 filter=15 channel=95
    -16, -15, -17, 13, -44, -8, -11, -38, 12,
    -- layer=1 filter=15 channel=96
    -9, -13, -17, 6, -6, -5, -8, -5, -10,
    -- layer=1 filter=15 channel=97
    -16, 0, 9, -12, 1, -1, -5, 9, 3,
    -- layer=1 filter=15 channel=98
    8, -9, 3, 0, 5, -15, 6, -5, 2,
    -- layer=1 filter=15 channel=99
    29, 38, 46, 17, 37, 40, 40, 51, -2,
    -- layer=1 filter=15 channel=100
    -25, -13, -5, -14, -31, -13, -5, 8, 20,
    -- layer=1 filter=15 channel=101
    10, -8, 6, 0, -1, -2, -7, -8, 0,
    -- layer=1 filter=15 channel=102
    -15, -8, 5, -19, -4, -10, -17, 4, 0,
    -- layer=1 filter=15 channel=103
    -27, -16, -7, -9, -23, -19, -30, -10, -11,
    -- layer=1 filter=15 channel=104
    -11, 23, 20, 25, 48, 44, -12, -3, 50,
    -- layer=1 filter=15 channel=105
    -11, -8, 3, -18, 4, 3, 7, 8, 3,
    -- layer=1 filter=15 channel=106
    -4, -7, -7, 0, -19, 14, 1, -27, 16,
    -- layer=1 filter=15 channel=107
    -16, 0, -6, -14, 1, -3, -6, -2, -11,
    -- layer=1 filter=15 channel=108
    2, 19, 14, -8, -11, 36, -21, -22, 26,
    -- layer=1 filter=15 channel=109
    -3, -4, -7, -1, -7, -1, 7, 0, 5,
    -- layer=1 filter=15 channel=110
    1, 2, -6, -6, 0, -3, -11, -11, -7,
    -- layer=1 filter=15 channel=111
    -4, 0, -45, 9, -7, -10, -18, -19, -4,
    -- layer=1 filter=15 channel=112
    6, -9, -37, 21, -31, -3, -18, -6, 30,
    -- layer=1 filter=15 channel=113
    -27, 2, 6, -14, -3, 9, -27, 10, 1,
    -- layer=1 filter=15 channel=114
    6, -47, -35, -11, -31, -64, -2, -13, -19,
    -- layer=1 filter=15 channel=115
    2, 6, 10, -9, 6, -14, 7, 30, -5,
    -- layer=1 filter=15 channel=116
    1, 1, 0, 10, 1, 8, 4, -7, -1,
    -- layer=1 filter=15 channel=117
    14, -45, -50, -1, -37, -16, -5, -13, -17,
    -- layer=1 filter=15 channel=118
    -1, 11, -23, 21, 0, -9, -7, -19, 2,
    -- layer=1 filter=15 channel=119
    16, 25, 9, 13, 11, 37, -18, -1, 29,
    -- layer=1 filter=15 channel=120
    3, -4, -2, -20, 4, -15, -5, -6, -7,
    -- layer=1 filter=15 channel=121
    -23, -24, -16, -8, -26, -15, 10, -10, 1,
    -- layer=1 filter=15 channel=122
    -8, 10, -7, -2, 4, -7, 3, 1, -3,
    -- layer=1 filter=15 channel=123
    -40, -32, -8, -7, -19, -14, -4, -7, -1,
    -- layer=1 filter=15 channel=124
    -2, -3, 10, -3, 13, 0, 16, -5, -1,
    -- layer=1 filter=15 channel=125
    -40, -41, -26, -11, -7, -10, -33, -25, -7,
    -- layer=1 filter=15 channel=126
    -17, -29, -8, -17, -15, -28, -12, -35, -39,
    -- layer=1 filter=15 channel=127
    -15, 11, -40, 15, -23, -5, -1, -46, 8,
    -- layer=1 filter=16 channel=0
    6, -5, 4, 7, 4, 5, -7, 4, 1,
    -- layer=1 filter=16 channel=1
    7, -8, 7, 4, -9, 7, 0, -9, 4,
    -- layer=1 filter=16 channel=2
    1, -3, 4, 5, 0, 16, 1, 6, -1,
    -- layer=1 filter=16 channel=3
    -8, -3, 0, -9, -9, 2, -7, -3, 2,
    -- layer=1 filter=16 channel=4
    -2, 5, 1, 4, -1, 4, 5, -10, 9,
    -- layer=1 filter=16 channel=5
    -11, -10, -18, 13, 9, 5, 3, -12, -1,
    -- layer=1 filter=16 channel=6
    -2, -10, -4, 8, 7, -4, 0, 4, -7,
    -- layer=1 filter=16 channel=7
    -13, -9, 10, 8, -5, 6, -9, 1, 0,
    -- layer=1 filter=16 channel=8
    -6, -6, 1, 6, 0, 2, -4, -10, -2,
    -- layer=1 filter=16 channel=9
    -12, -11, 0, -3, 9, -5, -5, -16, -6,
    -- layer=1 filter=16 channel=10
    0, 0, 14, -3, 1, 3, -11, 5, -10,
    -- layer=1 filter=16 channel=11
    -2, -11, -15, -13, 2, -10, -9, -3, 3,
    -- layer=1 filter=16 channel=12
    -2, -8, 0, -5, 11, 0, -8, 8, 0,
    -- layer=1 filter=16 channel=13
    1, 0, 0, 6, -2, -3, -8, -10, -9,
    -- layer=1 filter=16 channel=14
    -5, -5, 6, -5, 3, 4, 5, 9, -4,
    -- layer=1 filter=16 channel=15
    5, 9, 0, -2, -10, 8, -14, 0, 0,
    -- layer=1 filter=16 channel=16
    1, 0, -6, -7, 0, 5, -10, 2, 1,
    -- layer=1 filter=16 channel=17
    2, 0, 0, -6, 4, 7, -7, 6, -12,
    -- layer=1 filter=16 channel=18
    -2, -5, 8, -3, 7, -13, 0, 7, 0,
    -- layer=1 filter=16 channel=19
    2, -11, -4, 6, 7, 6, 0, 6, -6,
    -- layer=1 filter=16 channel=20
    6, -12, 1, -9, 3, -8, -4, -6, 4,
    -- layer=1 filter=16 channel=21
    0, 4, -3, -10, 3, -6, -4, -13, -9,
    -- layer=1 filter=16 channel=22
    -2, 3, -8, 4, 4, 7, -6, 0, -9,
    -- layer=1 filter=16 channel=23
    -4, 1, -12, 6, -2, 6, -1, -9, 3,
    -- layer=1 filter=16 channel=24
    0, 4, -10, -2, 4, -6, 6, -11, -2,
    -- layer=1 filter=16 channel=25
    -5, -1, -5, -9, 8, -3, -13, 5, -2,
    -- layer=1 filter=16 channel=26
    3, 3, 0, -3, -1, -6, -8, 2, -4,
    -- layer=1 filter=16 channel=27
    -9, 0, -6, -5, 4, -6, -2, -13, -4,
    -- layer=1 filter=16 channel=28
    -11, -10, -3, 4, 0, 5, 7, -1, 5,
    -- layer=1 filter=16 channel=29
    0, -1, 9, 8, -1, 1, 5, -7, 4,
    -- layer=1 filter=16 channel=30
    -15, -5, -7, 13, 11, 7, 4, -5, 12,
    -- layer=1 filter=16 channel=31
    -12, -2, 1, -6, -7, 0, 7, -7, -4,
    -- layer=1 filter=16 channel=32
    -7, -5, -6, -5, 7, 2, 4, -10, 5,
    -- layer=1 filter=16 channel=33
    -7, 8, -1, 0, -2, 0, -5, -4, -3,
    -- layer=1 filter=16 channel=34
    1, 2, 2, -9, 5, 1, -5, 0, -7,
    -- layer=1 filter=16 channel=35
    3, 4, -1, -3, 2, 5, -7, -8, -3,
    -- layer=1 filter=16 channel=36
    -13, 0, 0, -9, -6, -5, 0, -7, 3,
    -- layer=1 filter=16 channel=37
    -1, -6, -13, 0, -2, -6, -7, -2, 1,
    -- layer=1 filter=16 channel=38
    7, 6, -4, 5, 5, -7, 0, -7, -10,
    -- layer=1 filter=16 channel=39
    7, 2, -11, -11, 5, 6, 1, -7, -7,
    -- layer=1 filter=16 channel=40
    1, -10, -5, 10, 4, 1, -9, 7, -3,
    -- layer=1 filter=16 channel=41
    -8, 6, 8, 5, -10, -8, 0, 8, -6,
    -- layer=1 filter=16 channel=42
    9, 0, 3, -8, 0, 0, -1, -2, 6,
    -- layer=1 filter=16 channel=43
    2, -5, 3, 2, 0, -8, -7, -3, 0,
    -- layer=1 filter=16 channel=44
    -4, 3, 1, -12, -2, 0, 7, -11, -11,
    -- layer=1 filter=16 channel=45
    -6, -2, 1, 2, 5, 6, -11, 1, 3,
    -- layer=1 filter=16 channel=46
    -10, -4, -6, -6, -3, -13, -7, 1, 4,
    -- layer=1 filter=16 channel=47
    -2, -10, -21, 5, 0, 0, -6, -13, -1,
    -- layer=1 filter=16 channel=48
    -12, -6, -4, -12, -3, -13, -4, 4, -9,
    -- layer=1 filter=16 channel=49
    -14, -9, -1, 2, -4, 2, 0, -7, 1,
    -- layer=1 filter=16 channel=50
    -4, 7, -6, -6, -5, -11, -6, 8, -2,
    -- layer=1 filter=16 channel=51
    -6, -5, -7, 5, -14, 3, 3, 2, -4,
    -- layer=1 filter=16 channel=52
    5, -14, 0, 2, -9, -9, -1, -7, -10,
    -- layer=1 filter=16 channel=53
    0, 0, -10, 3, -6, 0, -8, 9, 0,
    -- layer=1 filter=16 channel=54
    3, -2, -8, 1, -3, -5, -11, -4, -11,
    -- layer=1 filter=16 channel=55
    -4, -18, -3, 0, -7, 0, 4, 0, -6,
    -- layer=1 filter=16 channel=56
    -8, 3, 6, -8, -8, 3, -1, 1, 8,
    -- layer=1 filter=16 channel=57
    -2, -11, 1, 4, 0, 6, -13, 2, -7,
    -- layer=1 filter=16 channel=58
    -5, -15, -1, -1, -4, -2, 4, -5, 3,
    -- layer=1 filter=16 channel=59
    4, 3, -2, -4, -5, 2, 3, -10, 3,
    -- layer=1 filter=16 channel=60
    -5, 6, 1, 5, -3, 6, -7, -4, -4,
    -- layer=1 filter=16 channel=61
    -10, 0, -4, 0, 3, 9, -8, -2, 0,
    -- layer=1 filter=16 channel=62
    -11, -8, 0, 6, 7, -4, -4, -1, -5,
    -- layer=1 filter=16 channel=63
    3, 1, -2, -5, 1, -4, 0, -8, 6,
    -- layer=1 filter=16 channel=64
    5, -1, -4, 0, 0, -11, -6, -5, -12,
    -- layer=1 filter=16 channel=65
    -13, -7, -8, 2, -10, 5, -8, -4, 0,
    -- layer=1 filter=16 channel=66
    -3, -2, 0, -14, -14, -7, -2, -3, -8,
    -- layer=1 filter=16 channel=67
    1, -4, -4, -1, -4, -6, -6, 1, -11,
    -- layer=1 filter=16 channel=68
    -2, -4, -4, -5, 0, 3, -7, 1, -12,
    -- layer=1 filter=16 channel=69
    -13, -14, -6, 2, 8, -7, 3, -5, -4,
    -- layer=1 filter=16 channel=70
    4, -2, 13, 0, 0, -5, -3, -5, 14,
    -- layer=1 filter=16 channel=71
    0, 6, -2, 7, 1, 5, -12, -11, 5,
    -- layer=1 filter=16 channel=72
    -8, -5, -2, -1, 0, -14, -12, -5, -9,
    -- layer=1 filter=16 channel=73
    -6, -9, 8, 6, -4, 2, -3, -7, 2,
    -- layer=1 filter=16 channel=74
    0, -4, -3, 6, 3, 2, 0, -2, 7,
    -- layer=1 filter=16 channel=75
    -5, -7, 9, 16, -7, 6, -9, -7, -4,
    -- layer=1 filter=16 channel=76
    -8, 0, 3, -5, -1, -7, 2, 0, 2,
    -- layer=1 filter=16 channel=77
    7, 7, 5, 1, -3, 5, 6, 5, -3,
    -- layer=1 filter=16 channel=78
    2, 5, -4, 8, -11, 2, 8, 2, 5,
    -- layer=1 filter=16 channel=79
    -5, -6, -2, 3, 7, -1, 1, 3, -2,
    -- layer=1 filter=16 channel=80
    7, -6, 4, -4, 6, 6, 6, 0, -8,
    -- layer=1 filter=16 channel=81
    -6, 0, -8, 0, -11, -1, -6, 0, -5,
    -- layer=1 filter=16 channel=82
    1, -8, -8, -8, 1, -2, 0, 0, 0,
    -- layer=1 filter=16 channel=83
    -7, 2, -9, -10, -2, 3, 0, -9, -7,
    -- layer=1 filter=16 channel=84
    0, -7, 7, 12, 4, 2, -5, -10, 3,
    -- layer=1 filter=16 channel=85
    3, -2, 3, -3, -6, 0, -9, 3, 0,
    -- layer=1 filter=16 channel=86
    -7, 5, 3, 0, -10, -2, 0, -3, -12,
    -- layer=1 filter=16 channel=87
    -6, -10, 0, -11, -6, 6, -3, 0, -8,
    -- layer=1 filter=16 channel=88
    -13, -14, -6, -13, -9, -8, -1, 5, -7,
    -- layer=1 filter=16 channel=89
    -3, 2, -14, 0, -6, -7, 2, -4, -14,
    -- layer=1 filter=16 channel=90
    3, 6, -8, -3, -2, -8, 4, -7, -3,
    -- layer=1 filter=16 channel=91
    2, -10, 0, 3, -4, -6, -11, -12, -15,
    -- layer=1 filter=16 channel=92
    2, -1, 4, -11, -2, -3, -3, -4, -7,
    -- layer=1 filter=16 channel=93
    -1, 1, -2, -11, -3, 0, -11, 4, -9,
    -- layer=1 filter=16 channel=94
    7, 5, -8, 5, -2, 3, -7, 7, -11,
    -- layer=1 filter=16 channel=95
    -16, 5, 0, -2, -4, 6, -14, -4, -3,
    -- layer=1 filter=16 channel=96
    -6, -2, 0, -13, 0, -4, 0, 0, -5,
    -- layer=1 filter=16 channel=97
    0, -7, -11, -12, -3, -4, -10, 0, 0,
    -- layer=1 filter=16 channel=98
    -8, -7, -12, 1, 12, -8, 0, -12, 0,
    -- layer=1 filter=16 channel=99
    -5, 1, -5, -4, 6, -3, 6, 5, -1,
    -- layer=1 filter=16 channel=100
    0, 6, -10, -12, -9, -9, -9, -10, 6,
    -- layer=1 filter=16 channel=101
    -11, 2, -4, -9, -8, -5, 6, -13, 0,
    -- layer=1 filter=16 channel=102
    1, -5, 6, -11, -2, -8, -3, -1, 0,
    -- layer=1 filter=16 channel=103
    -8, -7, -3, -7, -7, -8, -5, -13, -2,
    -- layer=1 filter=16 channel=104
    -1, -5, -12, 2, 0, 4, 1, -2, -4,
    -- layer=1 filter=16 channel=105
    -14, 0, 3, -12, 1, -8, 4, -9, -13,
    -- layer=1 filter=16 channel=106
    -12, -8, -9, -9, 0, 0, -5, -6, -7,
    -- layer=1 filter=16 channel=107
    -5, -1, 7, 6, 8, -6, 0, -11, -5,
    -- layer=1 filter=16 channel=108
    -14, 9, -12, -13, 0, -1, -8, -3, 6,
    -- layer=1 filter=16 channel=109
    -3, -8, 4, 1, -8, 9, -4, -9, -3,
    -- layer=1 filter=16 channel=110
    -10, -2, 0, 0, -7, -12, 5, -3, 5,
    -- layer=1 filter=16 channel=111
    -15, -5, 10, 0, -8, -6, 0, 9, 7,
    -- layer=1 filter=16 channel=112
    -10, 4, -7, -6, -10, -2, 7, -5, 8,
    -- layer=1 filter=16 channel=113
    1, 1, -6, 0, 6, 6, 3, -9, -9,
    -- layer=1 filter=16 channel=114
    0, -5, -7, 11, -5, -2, -9, -13, 1,
    -- layer=1 filter=16 channel=115
    1, -3, -5, 0, 3, -5, -10, 6, 3,
    -- layer=1 filter=16 channel=116
    8, 4, 9, -5, 9, -9, -6, 5, -9,
    -- layer=1 filter=16 channel=117
    -11, -6, 4, 9, 0, 3, 3, -7, -12,
    -- layer=1 filter=16 channel=118
    1, -5, 0, 4, -3, -4, 0, 4, 4,
    -- layer=1 filter=16 channel=119
    -5, 3, -2, -5, -2, -3, 6, -9, -4,
    -- layer=1 filter=16 channel=120
    6, -14, -8, -6, 3, -6, -16, 0, -16,
    -- layer=1 filter=16 channel=121
    -1, -4, 11, -8, -10, -5, -8, 2, -10,
    -- layer=1 filter=16 channel=122
    7, 0, 2, -4, 5, -4, -2, -7, 9,
    -- layer=1 filter=16 channel=123
    0, 4, 0, -3, 1, -4, -7, -11, 2,
    -- layer=1 filter=16 channel=124
    -4, -1, 4, 0, 0, -9, -4, -8, 1,
    -- layer=1 filter=16 channel=125
    -7, -12, -12, -3, -1, 9, -6, 0, -1,
    -- layer=1 filter=16 channel=126
    0, 0, -7, -4, 0, 1, -12, -7, -8,
    -- layer=1 filter=16 channel=127
    1, -13, -5, 4, -1, -1, -4, 12, 2,
    -- layer=1 filter=17 channel=0
    -24, -22, -8, -24, -24, -13, 3, 2, -11,
    -- layer=1 filter=17 channel=1
    3, 4, 0, -23, -3, 38, -1, -30, -13,
    -- layer=1 filter=17 channel=2
    18, 2, -13, 30, 15, 1, 23, 0, 15,
    -- layer=1 filter=17 channel=3
    -9, 4, -15, -1, 4, -5, -8, 8, 0,
    -- layer=1 filter=17 channel=4
    -5, 4, -7, -9, -2, 3, -2, -1, 4,
    -- layer=1 filter=17 channel=5
    -15, -1, -21, -19, 0, 14, 1, -60, 26,
    -- layer=1 filter=17 channel=6
    -5, -15, -7, -35, -39, -28, -66, -41, -35,
    -- layer=1 filter=17 channel=7
    9, 2, 8, 0, 16, -7, 17, 31, 15,
    -- layer=1 filter=17 channel=8
    10, -7, -6, -23, 22, 45, 7, -34, 25,
    -- layer=1 filter=17 channel=9
    5, -19, -33, -4, -14, -10, 1, -12, 19,
    -- layer=1 filter=17 channel=10
    9, 13, -11, 29, 23, 0, 22, 40, 9,
    -- layer=1 filter=17 channel=11
    -32, -35, -36, -32, -34, -46, -9, -27, -14,
    -- layer=1 filter=17 channel=12
    0, -3, -59, 32, 48, 23, -15, -26, -4,
    -- layer=1 filter=17 channel=13
    -3, 24, -5, 4, -8, 14, -15, -19, -2,
    -- layer=1 filter=17 channel=14
    35, 14, -13, -11, 0, -14, 48, 27, -40,
    -- layer=1 filter=17 channel=15
    -10, -7, -22, -50, -60, -36, -17, -50, -59,
    -- layer=1 filter=17 channel=16
    21, 6, 3, -14, 24, 25, 16, -30, 37,
    -- layer=1 filter=17 channel=17
    -20, -10, -20, 3, 14, 9, -8, 6, 19,
    -- layer=1 filter=17 channel=18
    16, 8, -20, 5, 10, 12, 19, -2, 15,
    -- layer=1 filter=17 channel=19
    -22, -8, -12, 9, -24, -38, -21, -17, 8,
    -- layer=1 filter=17 channel=20
    -6, 2, 11, -5, 10, 14, 7, -6, 9,
    -- layer=1 filter=17 channel=21
    5, 0, 25, 0, 0, 3, 22, 7, -3,
    -- layer=1 filter=17 channel=22
    2, -4, 1, -25, -13, 5, 3, -6, 4,
    -- layer=1 filter=17 channel=23
    13, -51, 5, -48, -22, -28, -44, -61, -20,
    -- layer=1 filter=17 channel=24
    -13, 19, -14, 3, -11, -12, -9, -17, 15,
    -- layer=1 filter=17 channel=25
    18, 6, -2, 21, 41, -2, 9, 28, 41,
    -- layer=1 filter=17 channel=26
    7, 20, -17, -12, -18, -17, -2, -24, 4,
    -- layer=1 filter=17 channel=27
    -49, -3, -39, -29, -18, -25, -48, -39, -46,
    -- layer=1 filter=17 channel=28
    17, 9, 16, 17, 32, 8, 19, 10, 1,
    -- layer=1 filter=17 channel=29
    -29, -12, -30, -5, -25, -19, -21, -41, -31,
    -- layer=1 filter=17 channel=30
    14, 32, -1, 5, 0, 24, 4, 15, 20,
    -- layer=1 filter=17 channel=31
    0, -44, -31, -10, 9, -16, -11, -12, 8,
    -- layer=1 filter=17 channel=32
    -15, 8, -42, -24, -30, -28, -48, -30, -9,
    -- layer=1 filter=17 channel=33
    -43, -26, -22, -9, -16, -16, -24, -8, -1,
    -- layer=1 filter=17 channel=34
    -59, -37, -13, -41, -19, -20, -43, -41, -8,
    -- layer=1 filter=17 channel=35
    8, 8, 12, 2, 0, 10, 8, 0, 15,
    -- layer=1 filter=17 channel=36
    -52, -40, -55, -51, -60, -59, -40, -46, -43,
    -- layer=1 filter=17 channel=37
    -8, -5, 1, 9, 5, -3, -12, -44, 22,
    -- layer=1 filter=17 channel=38
    13, 14, 9, 7, 5, 15, 0, -2, -2,
    -- layer=1 filter=17 channel=39
    -10, -20, -15, -9, -15, 3, -3, -12, -11,
    -- layer=1 filter=17 channel=40
    22, -10, -7, -19, -18, -14, -8, -18, -14,
    -- layer=1 filter=17 channel=41
    -10, 2, -30, -38, -48, -30, -43, -82, 12,
    -- layer=1 filter=17 channel=42
    5, -11, 0, 8, 3, -6, 7, 7, -14,
    -- layer=1 filter=17 channel=43
    8, 3, -7, 8, 30, 21, 6, -34, 25,
    -- layer=1 filter=17 channel=44
    -9, 3, -47, -33, -15, -19, -23, -17, -6,
    -- layer=1 filter=17 channel=45
    -2, 22, 8, -8, -3, 0, 11, -26, -12,
    -- layer=1 filter=17 channel=46
    -35, 4, 6, 32, 6, -70, 4, -13, -21,
    -- layer=1 filter=17 channel=47
    1, -19, -32, -47, -33, -23, -61, -41, -39,
    -- layer=1 filter=17 channel=48
    4, 11, 3, 7, 9, -2, -7, 11, -7,
    -- layer=1 filter=17 channel=49
    3, 7, 0, -4, -20, -18, -14, -11, -11,
    -- layer=1 filter=17 channel=50
    -16, -14, -15, -19, -12, -1, 1, -5, -4,
    -- layer=1 filter=17 channel=51
    9, 5, 9, 16, 13, -7, -7, 14, -1,
    -- layer=1 filter=17 channel=52
    -1, 0, -5, -3, -9, -4, -5, 12, 2,
    -- layer=1 filter=17 channel=53
    11, 1, 2, 11, 3, 3, 5, 17, 2,
    -- layer=1 filter=17 channel=54
    18, 13, -10, 32, 36, -9, 1, 14, 39,
    -- layer=1 filter=17 channel=55
    -38, -40, -59, -30, -49, -35, -20, -24, -43,
    -- layer=1 filter=17 channel=56
    8, 0, 8, 9, 2, -13, 0, 5, 2,
    -- layer=1 filter=17 channel=57
    20, 13, -19, 33, 12, 0, 10, 32, 0,
    -- layer=1 filter=17 channel=58
    0, -2, -6, -29, -6, -27, -60, 4, -14,
    -- layer=1 filter=17 channel=59
    13, 13, 9, -6, -2, 9, 12, -4, 0,
    -- layer=1 filter=17 channel=60
    -4, 9, -4, 0, -5, 8, -5, 19, -3,
    -- layer=1 filter=17 channel=61
    -7, 4, 2, 0, 9, -13, 3, 3, -5,
    -- layer=1 filter=17 channel=62
    18, 15, 7, 5, 45, 34, 16, -11, 49,
    -- layer=1 filter=17 channel=63
    -30, -42, -48, -59, -32, -30, -20, -19, -29,
    -- layer=1 filter=17 channel=64
    -11, -2, -4, -11, -5, 15, -17, -5, 3,
    -- layer=1 filter=17 channel=65
    -2, 0, 14, -5, -4, 4, 0, 2, 0,
    -- layer=1 filter=17 channel=66
    -44, -45, -17, -36, -22, -26, -7, -12, -2,
    -- layer=1 filter=17 channel=67
    -4, -6, -11, -19, -42, -27, -26, -31, -34,
    -- layer=1 filter=17 channel=68
    -15, -1, -51, -26, -20, -29, -25, -6, -8,
    -- layer=1 filter=17 channel=69
    31, 6, 2, -13, -4, -8, 23, -33, 11,
    -- layer=1 filter=17 channel=70
    -22, -40, -13, -36, -60, -56, -78, -63, -33,
    -- layer=1 filter=17 channel=71
    5, -4, 17, 5, 8, -17, 3, 6, 7,
    -- layer=1 filter=17 channel=72
    8, 6, -5, 20, 21, -28, -21, -20, 34,
    -- layer=1 filter=17 channel=73
    -7, -7, 6, -1, -7, -1, 4, 8, -4,
    -- layer=1 filter=17 channel=74
    29, -16, -15, 14, -15, -12, -33, -14, 5,
    -- layer=1 filter=17 channel=75
    30, 18, 0, 17, 66, -17, 16, -3, 11,
    -- layer=1 filter=17 channel=76
    -11, -8, -37, -23, -10, -30, -41, 5, 2,
    -- layer=1 filter=17 channel=77
    -6, 6, 1, -13, -8, 11, -11, 3, -1,
    -- layer=1 filter=17 channel=78
    4, -13, -11, -1, -10, -3, 23, -2, 3,
    -- layer=1 filter=17 channel=79
    9, 19, 9, -6, 34, 21, 2, -19, 32,
    -- layer=1 filter=17 channel=80
    -11, -1, -3, 5, 2, -4, 4, 0, -1,
    -- layer=1 filter=17 channel=81
    -12, -16, -7, -12, -3, -10, -23, -17, -3,
    -- layer=1 filter=17 channel=82
    3, 7, 15, -5, 6, 9, -5, 8, -5,
    -- layer=1 filter=17 channel=83
    0, -8, -3, -10, -12, 26, -2, -27, -21,
    -- layer=1 filter=17 channel=84
    7, 23, -27, -8, -13, 27, -25, 9, 36,
    -- layer=1 filter=17 channel=85
    -7, -15, -22, -28, 6, -28, -62, -20, -3,
    -- layer=1 filter=17 channel=86
    -26, -24, -22, -19, -15, -4, -8, -4, 1,
    -- layer=1 filter=17 channel=87
    -48, -9, -25, -8, -25, -12, -28, -25, -23,
    -- layer=1 filter=17 channel=88
    11, 2, -12, -12, -12, -15, -6, 7, -15,
    -- layer=1 filter=17 channel=89
    9, 2, 5, -14, -16, 2, -9, 8, -7,
    -- layer=1 filter=17 channel=90
    -15, -1, -34, -27, -25, -30, -19, -26, -23,
    -- layer=1 filter=17 channel=91
    18, 23, 18, 0, 11, 8, 1, 21, 21,
    -- layer=1 filter=17 channel=92
    -62, -66, -66, -30, -76, -68, -10, -21, -32,
    -- layer=1 filter=17 channel=93
    0, 3, 17, 9, 11, 6, 5, 14, 19,
    -- layer=1 filter=17 channel=94
    -17, -21, -14, -7, -24, -7, -2, -6, -6,
    -- layer=1 filter=17 channel=95
    20, -8, -33, -3, 3, 29, 11, 15, 19,
    -- layer=1 filter=17 channel=96
    0, -5, -3, -1, 0, 0, 2, 1, -4,
    -- layer=1 filter=17 channel=97
    -23, -16, -12, -5, -2, 8, 5, -1, 11,
    -- layer=1 filter=17 channel=98
    17, 0, -2, 6, 20, 24, 0, -14, 17,
    -- layer=1 filter=17 channel=99
    20, -1, -34, 15, -14, -15, 31, 11, -11,
    -- layer=1 filter=17 channel=100
    -30, -30, -35, -46, -13, -45, -34, -38, -27,
    -- layer=1 filter=17 channel=101
    11, 20, 26, 10, 9, 6, 8, 14, 10,
    -- layer=1 filter=17 channel=102
    2, -3, -5, -21, -22, 0, -7, 12, 15,
    -- layer=1 filter=17 channel=103
    -29, -32, -20, -26, -10, -17, -6, 1, -16,
    -- layer=1 filter=17 channel=104
    2, -19, -40, -45, -1, -36, -42, -45, -15,
    -- layer=1 filter=17 channel=105
    -26, -8, -18, -3, 0, -5, -12, 15, 1,
    -- layer=1 filter=17 channel=106
    -5, 16, 9, 0, -8, 5, -21, -9, 0,
    -- layer=1 filter=17 channel=107
    17, 10, 3, -3, -3, -10, -4, -4, 7,
    -- layer=1 filter=17 channel=108
    -14, -3, -31, -29, -55, -13, -10, -58, -18,
    -- layer=1 filter=17 channel=109
    -8, -1, 4, -3, -5, 0, -2, -7, -4,
    -- layer=1 filter=17 channel=110
    8, -7, 3, -8, -5, -5, 2, -4, -7,
    -- layer=1 filter=17 channel=111
    30, 23, -17, 9, -11, 41, 9, 24, 28,
    -- layer=1 filter=17 channel=112
    34, 7, -11, -5, -27, 37, -11, 25, -13,
    -- layer=1 filter=17 channel=113
    -53, -41, -26, -5, -3, -39, -19, -13, -33,
    -- layer=1 filter=17 channel=114
    -32, -26, -53, -64, -79, -54, -42, -87, -38,
    -- layer=1 filter=17 channel=115
    -4, -8, -14, 6, 4, -11, 8, 17, 14,
    -- layer=1 filter=17 channel=116
    -6, 0, 0, -3, 4, 2, -10, 3, 3,
    -- layer=1 filter=17 channel=117
    69, 55, -13, 10, -31, 40, 25, 66, 0,
    -- layer=1 filter=17 channel=118
    14, 25, -8, 17, -16, 17, -20, -12, 23,
    -- layer=1 filter=17 channel=119
    -24, 10, -42, -27, -40, -41, -45, -33, 0,
    -- layer=1 filter=17 channel=120
    6, 0, 13, 0, 16, 6, -11, 11, 8,
    -- layer=1 filter=17 channel=121
    -8, 12, -6, -14, 1, -20, 40, 6, -30,
    -- layer=1 filter=17 channel=122
    3, 1, -3, -2, -8, 0, -3, 7, -7,
    -- layer=1 filter=17 channel=123
    -23, -17, -36, -36, 22, -36, 0, -22, -48,
    -- layer=1 filter=17 channel=124
    -19, -1, 2, -10, -13, -18, -12, -20, -18,
    -- layer=1 filter=17 channel=125
    2, -13, -4, -20, -35, -41, -44, -33, -61,
    -- layer=1 filter=17 channel=126
    -5, -12, 11, -12, 20, 35, 3, -24, 12,
    -- layer=1 filter=17 channel=127
    19, 21, -5, 9, 25, 31, 5, -5, 37,
    -- layer=1 filter=18 channel=0
    -45, -50, -26, -39, -38, -53, -62, -52, -21,
    -- layer=1 filter=18 channel=1
    -42, -39, -47, -58, -39, -81, -39, -19, 35,
    -- layer=1 filter=18 channel=2
    36, 43, 21, 33, 34, 37, 52, 45, 21,
    -- layer=1 filter=18 channel=3
    -9, 0, -5, 6, 6, 0, -5, -3, -6,
    -- layer=1 filter=18 channel=4
    -1, -5, -6, -8, -7, -9, -8, -19, -8,
    -- layer=1 filter=18 channel=5
    -50, -43, -68, -104, -129, -60, -1, -1, 65,
    -- layer=1 filter=18 channel=6
    -9, -2, 28, -30, -16, -16, -13, -13, -37,
    -- layer=1 filter=18 channel=7
    -35, -39, 7, -76, -123, -31, -51, 15, 58,
    -- layer=1 filter=18 channel=8
    -33, -85, -89, -74, -128, -64, -32, -2, 66,
    -- layer=1 filter=18 channel=9
    30, -12, 20, 17, 41, 24, 58, 59, 19,
    -- layer=1 filter=18 channel=10
    -21, -30, 12, -50, -82, -2, -34, 41, 66,
    -- layer=1 filter=18 channel=11
    -61, -84, -50, -81, -70, -64, -69, -78, -51,
    -- layer=1 filter=18 channel=12
    9, 31, 11, -7, -18, 8, 32, -10, -9,
    -- layer=1 filter=18 channel=13
    -3, 0, 25, 5, 3, 20, 8, 14, 9,
    -- layer=1 filter=18 channel=14
    -16, 8, 39, -7, -46, 10, -50, -37, -37,
    -- layer=1 filter=18 channel=15
    -10, -71, -31, -53, -59, -22, -32, -43, -4,
    -- layer=1 filter=18 channel=16
    -46, -78, -105, -104, -123, -29, -13, 7, 68,
    -- layer=1 filter=18 channel=17
    -38, -12, -33, -19, -16, -31, -22, -10, 57,
    -- layer=1 filter=18 channel=18
    -23, -20, 6, -67, -56, -27, -30, 0, -49,
    -- layer=1 filter=18 channel=19
    -3, -77, -36, -78, -78, 19, 20, 40, 66,
    -- layer=1 filter=18 channel=20
    -16, 3, 5, -18, -16, 7, -5, 14, 44,
    -- layer=1 filter=18 channel=21
    17, 8, 9, 24, 10, 6, 4, 12, 14,
    -- layer=1 filter=18 channel=22
    -47, -41, -31, -34, -43, -25, -21, -16, 38,
    -- layer=1 filter=18 channel=23
    -14, -57, 4, -136, -108, 23, -54, 18, 28,
    -- layer=1 filter=18 channel=24
    23, 5, 13, 8, 11, 26, 4, 21, 16,
    -- layer=1 filter=18 channel=25
    -24, -61, -10, -54, -116, -10, -7, 38, 89,
    -- layer=1 filter=18 channel=26
    -45, -86, -11, -113, -64, -37, -53, -44, -42,
    -- layer=1 filter=18 channel=27
    14, -1, -5, 18, 25, 0, 27, 24, 26,
    -- layer=1 filter=18 channel=28
    -16, -37, -28, -36, -105, -23, -18, 2, 57,
    -- layer=1 filter=18 channel=29
    2, -21, -17, 8, -9, -8, -8, 7, 6,
    -- layer=1 filter=18 channel=30
    -8, -15, 0, -58, -35, -33, -21, -41, -67,
    -- layer=1 filter=18 channel=31
    6, 18, 21, 19, 1, -1, 32, 2, -23,
    -- layer=1 filter=18 channel=32
    -43, -78, 4, -153, -59, -51, -39, -54, -39,
    -- layer=1 filter=18 channel=33
    36, 6, 32, -21, -11, 22, 35, 36, 49,
    -- layer=1 filter=18 channel=34
    4, -9, -6, -22, -30, -21, -20, -24, -17,
    -- layer=1 filter=18 channel=35
    6, 3, 5, -13, 4, 10, 0, -3, 5,
    -- layer=1 filter=18 channel=36
    -66, -77, -47, -86, -64, -82, -31, -60, -33,
    -- layer=1 filter=18 channel=37
    -16, -57, -51, -111, -124, -18, 8, 33, 75,
    -- layer=1 filter=18 channel=38
    5, 27, 19, 11, 22, 20, 7, 23, 28,
    -- layer=1 filter=18 channel=39
    -10, -13, -11, 5, 13, -26, -36, -34, -5,
    -- layer=1 filter=18 channel=40
    -17, -11, 11, -24, -22, -6, 0, -14, -34,
    -- layer=1 filter=18 channel=41
    -17, -54, 21, -76, -13, 11, 5, 30, 26,
    -- layer=1 filter=18 channel=42
    37, 40, 18, 45, 45, 40, 57, 52, 33,
    -- layer=1 filter=18 channel=43
    -20, -70, -81, -83, -118, -43, -13, -17, 60,
    -- layer=1 filter=18 channel=44
    -122, -120, -14, -152, -92, -82, -79, -69, -31,
    -- layer=1 filter=18 channel=45
    -5, 18, 15, -20, -7, 3, 1, 0, -7,
    -- layer=1 filter=18 channel=46
    13, 9, -3, -15, -30, 40, 42, 51, 63,
    -- layer=1 filter=18 channel=47
    0, 5, 32, -27, 12, 57, 32, 56, 61,
    -- layer=1 filter=18 channel=48
    3, 3, 4, 11, -2, -6, -11, 5, -9,
    -- layer=1 filter=18 channel=49
    39, 24, 41, 23, 33, 48, 42, 40, 35,
    -- layer=1 filter=18 channel=50
    31, 9, 22, 42, 13, 14, 36, 8, 9,
    -- layer=1 filter=18 channel=51
    18, 21, 23, 18, 9, 0, 4, 19, 24,
    -- layer=1 filter=18 channel=52
    -21, -7, -22, -9, -19, -6, -3, -6, 0,
    -- layer=1 filter=18 channel=53
    -8, -4, -5, 1, -12, -5, -5, -2, -3,
    -- layer=1 filter=18 channel=54
    21, -41, -9, -4, -55, 13, 17, 68, 101,
    -- layer=1 filter=18 channel=55
    8, 12, 12, -9, 2, 6, 1, 25, 14,
    -- layer=1 filter=18 channel=56
    -7, 5, -10, 0, -6, 3, -1, 6, -8,
    -- layer=1 filter=18 channel=57
    1, -28, -1, 0, -46, -13, -23, 27, 60,
    -- layer=1 filter=18 channel=58
    -6, -69, -7, -69, -40, 22, -23, 82, 82,
    -- layer=1 filter=18 channel=59
    2, -4, -9, -11, 1, -21, -14, -10, 1,
    -- layer=1 filter=18 channel=60
    -13, 0, -2, -11, -19, -29, 5, -20, -16,
    -- layer=1 filter=18 channel=61
    7, -1, 7, -6, 7, 5, -1, -10, 6,
    -- layer=1 filter=18 channel=62
    -45, -90, -93, -123, -146, -37, -6, 14, 79,
    -- layer=1 filter=18 channel=63
    -46, -42, -45, -16, -13, -8, -23, -21, -24,
    -- layer=1 filter=18 channel=64
    -4, 10, 6, -11, -16, -14, 3, -4, 25,
    -- layer=1 filter=18 channel=65
    0, 6, -9, 2, -4, -5, 0, -17, -4,
    -- layer=1 filter=18 channel=66
    -32, -27, -35, -14, -35, -29, -34, -54, -14,
    -- layer=1 filter=18 channel=67
    21, 25, 12, 15, 5, 16, 23, 21, 2,
    -- layer=1 filter=18 channel=68
    -122, -118, -5, -123, -70, -67, -74, -44, -50,
    -- layer=1 filter=18 channel=69
    -30, -52, -21, -81, -67, -27, -12, 1, 32,
    -- layer=1 filter=18 channel=70
    5, 16, 45, -36, -33, -25, -32, -42, -33,
    -- layer=1 filter=18 channel=71
    33, 25, 6, 17, 15, 11, 14, 15, 21,
    -- layer=1 filter=18 channel=72
    -3, -31, -4, -73, -56, -36, 17, 5, 25,
    -- layer=1 filter=18 channel=73
    5, -4, 4, -11, 0, -9, 3, 1, -5,
    -- layer=1 filter=18 channel=74
    -22, -28, 15, -74, -45, -33, 17, 0, -48,
    -- layer=1 filter=18 channel=75
    -6, 25, 17, 9, 4, 19, 26, 27, 4,
    -- layer=1 filter=18 channel=76
    -57, -68, -14, -80, -55, -67, -59, -60, -63,
    -- layer=1 filter=18 channel=77
    -5, 0, -1, -1, -8, -2, -24, -8, 0,
    -- layer=1 filter=18 channel=78
    -6, -20, -22, -22, 2, -3, -18, 20, 12,
    -- layer=1 filter=18 channel=79
    -31, -89, -88, -98, -137, -25, -5, 22, 74,
    -- layer=1 filter=18 channel=80
    -20, 9, 38, -9, 0, 11, 6, -21, 31,
    -- layer=1 filter=18 channel=81
    0, -5, -9, 0, 2, -7, -16, 7, 5,
    -- layer=1 filter=18 channel=82
    21, 11, 7, 11, 14, 5, 9, 9, 5,
    -- layer=1 filter=18 channel=83
    -62, -49, -75, -69, -34, -64, -44, -41, -18,
    -- layer=1 filter=18 channel=84
    -39, -45, 9, -67, -40, -61, -43, -23, -50,
    -- layer=1 filter=18 channel=85
    -2, -34, -26, -75, -22, 51, -30, 78, 90,
    -- layer=1 filter=18 channel=86
    -50, -33, -60, -70, -67, -43, -17, -7, 11,
    -- layer=1 filter=18 channel=87
    35, -4, 21, -15, 5, 19, 45, 83, 71,
    -- layer=1 filter=18 channel=88
    16, 26, 11, 15, 9, 26, 14, 9, 5,
    -- layer=1 filter=18 channel=89
    3, 5, 17, 2, 6, 1, 1, 7, -7,
    -- layer=1 filter=18 channel=90
    -103, -101, -37, -148, -100, -94, -82, -72, -35,
    -- layer=1 filter=18 channel=91
    6, 17, 20, 8, 8, 5, 7, 21, 20,
    -- layer=1 filter=18 channel=92
    -22, -30, -3, -48, -46, -29, 20, -13, 13,
    -- layer=1 filter=18 channel=93
    8, 14, 11, 7, 11, 0, 1, 5, 23,
    -- layer=1 filter=18 channel=94
    -7, 0, -4, -35, -25, -34, -5, -28, -16,
    -- layer=1 filter=18 channel=95
    -58, -47, -27, -64, -71, -50, -32, -80, -61,
    -- layer=1 filter=18 channel=96
    15, 0, -13, 21, 10, -8, 16, 9, 10,
    -- layer=1 filter=18 channel=97
    -20, -17, -23, -20, -27, -26, -28, -21, 2,
    -- layer=1 filter=18 channel=98
    -18, -77, -82, -44, -108, -45, -20, 15, 74,
    -- layer=1 filter=18 channel=99
    -28, -48, -15, -17, -40, -64, -46, -20, 12,
    -- layer=1 filter=18 channel=100
    -83, -84, -95, -77, -53, -62, -10, -40, 0,
    -- layer=1 filter=18 channel=101
    7, 21, 30, 1, 19, 14, 15, 19, 12,
    -- layer=1 filter=18 channel=102
    -57, -29, -17, -51, -50, -61, -48, -56, -64,
    -- layer=1 filter=18 channel=103
    -27, -73, -64, -63, -59, -43, -16, -65, -23,
    -- layer=1 filter=18 channel=104
    10, -8, -10, -80, -1, 21, -35, 5, 19,
    -- layer=1 filter=18 channel=105
    -21, -25, -19, -5, -24, -51, -25, -35, -13,
    -- layer=1 filter=18 channel=106
    0, 13, 26, -7, 4, 25, -1, 0, 5,
    -- layer=1 filter=18 channel=107
    10, 9, 15, 10, 6, 10, 0, -1, 0,
    -- layer=1 filter=18 channel=108
    -41, -59, 3, -108, -32, -36, -33, -22, -15,
    -- layer=1 filter=18 channel=109
    -2, -1, -1, 0, 0, 6, 5, -8, 6,
    -- layer=1 filter=18 channel=110
    -3, 12, -3, -16, -24, -12, -9, -7, 3,
    -- layer=1 filter=18 channel=111
    -27, -49, 8, -39, -37, -52, -45, -38, -62,
    -- layer=1 filter=18 channel=112
    -60, -57, -9, -8, -58, -27, -27, -38, -29,
    -- layer=1 filter=18 channel=113
    25, 29, 6, 30, 20, 30, 38, 51, 38,
    -- layer=1 filter=18 channel=114
    -58, -42, -63, -105, -108, -45, -26, -8, 16,
    -- layer=1 filter=18 channel=115
    -33, -12, 1, -32, -76, -27, -4, 3, 35,
    -- layer=1 filter=18 channel=116
    -2, 2, -2, -6, 9, 7, 0, -3, -4,
    -- layer=1 filter=18 channel=117
    -49, -60, 2, -49, -47, -63, -51, -29, -49,
    -- layer=1 filter=18 channel=118
    2, -27, 13, -64, -24, -41, -18, -21, -47,
    -- layer=1 filter=18 channel=119
    -57, -69, -18, -145, -70, -55, -74, -50, -39,
    -- layer=1 filter=18 channel=120
    8, 18, 10, 5, -1, 6, 5, 14, 41,
    -- layer=1 filter=18 channel=121
    0, -7, -32, -4, -7, 21, 29, 8, 3,
    -- layer=1 filter=18 channel=122
    -5, 2, 1, 3, 10, 6, 0, -7, 7,
    -- layer=1 filter=18 channel=123
    0, 1, -22, 0, -4, 1, 27, 20, -7,
    -- layer=1 filter=18 channel=124
    1, -12, 18, 6, 6, 0, -13, 3, 6,
    -- layer=1 filter=18 channel=125
    5, 17, 42, -22, -27, -20, -18, -15, -13,
    -- layer=1 filter=18 channel=126
    -43, -67, -73, -26, -51, -59, -65, -32, 62,
    -- layer=1 filter=18 channel=127
    10, -14, 1, -54, -25, -13, -10, -30, -61,
    -- layer=1 filter=19 channel=0
    3, 4, -10, -7, -5, -7, -10, 2, -1,
    -- layer=1 filter=19 channel=1
    -7, 0, 1, -7, -1, -9, 0, -2, -6,
    -- layer=1 filter=19 channel=2
    17, 9, -5, -5, -5, 1, -6, 6, 9,
    -- layer=1 filter=19 channel=3
    5, 8, -10, 4, -8, -8, 0, -5, 5,
    -- layer=1 filter=19 channel=4
    2, -5, -7, -3, 1, 2, 4, 3, 0,
    -- layer=1 filter=19 channel=5
    -10, -17, 2, -7, 1, 3, 0, -3, 1,
    -- layer=1 filter=19 channel=6
    7, 1, -4, -1, 0, 1, 0, 0, -4,
    -- layer=1 filter=19 channel=7
    3, -4, -9, -13, 2, 9, -1, -2, -2,
    -- layer=1 filter=19 channel=8
    7, -13, -13, -6, -10, 7, -10, -8, 0,
    -- layer=1 filter=19 channel=9
    -3, 0, 4, 2, 1, 0, 0, 7, -1,
    -- layer=1 filter=19 channel=10
    17, -1, 5, -8, 3, 3, -8, -10, -9,
    -- layer=1 filter=19 channel=11
    0, -11, -1, 3, -2, -4, -9, -3, -8,
    -- layer=1 filter=19 channel=12
    -3, -1, 0, -2, 1, -7, 1, 5, 0,
    -- layer=1 filter=19 channel=13
    1, -11, 3, -8, 2, 6, -5, -3, -9,
    -- layer=1 filter=19 channel=14
    5, 17, 3, 9, -7, -10, -3, -5, -11,
    -- layer=1 filter=19 channel=15
    -6, -10, -1, 4, -11, 6, -12, -5, 8,
    -- layer=1 filter=19 channel=16
    -11, -5, -1, -5, 4, -11, -15, -8, -6,
    -- layer=1 filter=19 channel=17
    -8, 1, 4, -8, -11, -8, -12, -2, -8,
    -- layer=1 filter=19 channel=18
    -2, 10, 1, -9, 0, -21, 7, 5, -13,
    -- layer=1 filter=19 channel=19
    5, -9, 7, 7, 0, -10, -11, 1, 1,
    -- layer=1 filter=19 channel=20
    -3, -12, 2, -14, -3, -1, 4, 1, -1,
    -- layer=1 filter=19 channel=21
    -1, -14, -17, -5, -6, -4, -1, 0, -9,
    -- layer=1 filter=19 channel=22
    0, 4, -9, -5, -6, 1, -7, 1, -5,
    -- layer=1 filter=19 channel=23
    -1, -2, -5, -9, 6, 4, 2, -2, -5,
    -- layer=1 filter=19 channel=24
    0, -10, -11, -9, 1, -4, -3, -3, -14,
    -- layer=1 filter=19 channel=25
    -1, -12, -1, -7, -13, -4, -1, -9, 0,
    -- layer=1 filter=19 channel=26
    -6, -8, -8, 3, -11, 3, -13, 2, 0,
    -- layer=1 filter=19 channel=27
    -1, 4, -10, 9, 0, 4, -5, -10, 3,
    -- layer=1 filter=19 channel=28
    -4, -16, 2, -16, -10, -12, -15, -6, -5,
    -- layer=1 filter=19 channel=29
    -4, 2, -6, 6, -5, 7, -4, 1, -6,
    -- layer=1 filter=19 channel=30
    -9, 2, 10, -12, 2, -6, -6, -7, -9,
    -- layer=1 filter=19 channel=31
    0, 2, 0, -12, 1, -7, 1, -3, -3,
    -- layer=1 filter=19 channel=32
    -10, 4, 2, -2, 1, 0, -12, -14, -2,
    -- layer=1 filter=19 channel=33
    -9, 2, -2, -1, 0, -7, -9, 11, -3,
    -- layer=1 filter=19 channel=34
    -4, -6, -3, -10, 3, 2, -3, 6, -5,
    -- layer=1 filter=19 channel=35
    8, 2, 7, 4, -8, -1, 0, -10, 8,
    -- layer=1 filter=19 channel=36
    -5, -2, -11, 2, -8, 3, -11, -1, -1,
    -- layer=1 filter=19 channel=37
    -3, -13, -15, -3, -7, 0, -5, 6, 0,
    -- layer=1 filter=19 channel=38
    -8, 0, 4, 0, -15, -4, -2, -9, -4,
    -- layer=1 filter=19 channel=39
    6, 7, -7, 0, 4, 6, 2, -10, -10,
    -- layer=1 filter=19 channel=40
    -5, -8, -2, 3, 4, 3, -8, -12, 9,
    -- layer=1 filter=19 channel=41
    3, 0, -7, -6, -7, -11, -6, -6, -3,
    -- layer=1 filter=19 channel=42
    -5, 0, 1, 9, -2, 0, -4, -1, -9,
    -- layer=1 filter=19 channel=43
    -2, -15, -13, -4, 7, -13, -6, -9, -14,
    -- layer=1 filter=19 channel=44
    -13, 8, -13, -8, -10, -7, -9, -14, -3,
    -- layer=1 filter=19 channel=45
    0, 5, -7, 2, -6, -3, -6, -15, 2,
    -- layer=1 filter=19 channel=46
    1, 3, 9, -2, -3, 4, -9, 2, -9,
    -- layer=1 filter=19 channel=47
    -4, -11, 2, -6, -6, -13, -18, -6, -13,
    -- layer=1 filter=19 channel=48
    -9, 4, -7, -11, -3, -5, 5, -3, -11,
    -- layer=1 filter=19 channel=49
    -7, 0, 5, 3, 0, 3, -1, -1, -5,
    -- layer=1 filter=19 channel=50
    -6, -8, -3, -2, -9, -8, -8, 1, 8,
    -- layer=1 filter=19 channel=51
    4, -6, -1, -2, -4, -13, -6, -15, -10,
    -- layer=1 filter=19 channel=52
    3, 4, 10, -8, 0, 8, 0, -5, 0,
    -- layer=1 filter=19 channel=53
    1, 0, -9, -12, 4, 8, -12, -4, -7,
    -- layer=1 filter=19 channel=54
    -3, -7, -6, 6, -8, -2, 4, -14, -13,
    -- layer=1 filter=19 channel=55
    0, -9, -11, -4, 7, -4, -3, -10, -12,
    -- layer=1 filter=19 channel=56
    -8, -3, 3, 4, -7, 5, -1, -9, -5,
    -- layer=1 filter=19 channel=57
    4, 1, -2, -6, 4, -11, -4, -6, -7,
    -- layer=1 filter=19 channel=58
    -7, -17, 17, -6, -9, 5, -13, -9, 0,
    -- layer=1 filter=19 channel=59
    -8, 8, 0, -7, 1, 8, -6, 3, 6,
    -- layer=1 filter=19 channel=60
    -1, 4, 0, 8, 3, 8, 2, -7, 1,
    -- layer=1 filter=19 channel=61
    -2, 8, 3, 0, -4, 0, -10, -8, -2,
    -- layer=1 filter=19 channel=62
    -3, -11, -16, -13, 2, -5, 0, -10, 0,
    -- layer=1 filter=19 channel=63
    -12, 6, 4, -6, 2, 2, -8, 3, 2,
    -- layer=1 filter=19 channel=64
    -10, -4, 0, -10, -5, 1, -14, 6, 0,
    -- layer=1 filter=19 channel=65
    4, 5, 2, 3, -9, -8, -8, 1, 1,
    -- layer=1 filter=19 channel=66
    -4, -10, -10, -7, -9, -6, 2, -10, -11,
    -- layer=1 filter=19 channel=67
    0, -9, -9, -10, -7, -16, -4, 1, -15,
    -- layer=1 filter=19 channel=68
    -11, 5, -9, -5, -7, -8, 5, -6, 2,
    -- layer=1 filter=19 channel=69
    -17, -12, 5, -3, -4, -2, -23, -4, -2,
    -- layer=1 filter=19 channel=70
    4, 3, 0, 2, 6, 2, -13, -1, -3,
    -- layer=1 filter=19 channel=71
    -14, -4, 3, 0, 5, -1, 2, -7, -9,
    -- layer=1 filter=19 channel=72
    -10, -4, 6, -15, -7, 6, -7, -11, 0,
    -- layer=1 filter=19 channel=73
    -4, -11, 3, 2, 6, -11, -5, -1, 7,
    -- layer=1 filter=19 channel=74
    -11, -8, -4, -9, 2, -13, -7, 4, -12,
    -- layer=1 filter=19 channel=75
    -7, -1, 6, 7, 12, -16, 0, 4, 10,
    -- layer=1 filter=19 channel=76
    1, -2, -12, -6, -1, 0, 4, 2, 8,
    -- layer=1 filter=19 channel=77
    3, 0, -7, -14, -1, -12, -9, -13, 6,
    -- layer=1 filter=19 channel=78
    -8, -8, -7, 3, 6, 2, 5, -8, 7,
    -- layer=1 filter=19 channel=79
    -6, -7, -3, -4, -14, 5, -13, -5, 1,
    -- layer=1 filter=19 channel=80
    -7, -9, 9, -7, -3, -10, 5, -10, 7,
    -- layer=1 filter=19 channel=81
    5, -8, -2, -6, 5, 4, -5, -11, 0,
    -- layer=1 filter=19 channel=82
    -3, 4, 0, 0, -14, 3, 3, -12, -3,
    -- layer=1 filter=19 channel=83
    2, 0, 6, 5, 3, 7, 6, 2, -9,
    -- layer=1 filter=19 channel=84
    -5, 12, 1, -7, 5, -10, 4, -9, -8,
    -- layer=1 filter=19 channel=85
    1, -10, 9, 1, 7, 3, 10, 7, -2,
    -- layer=1 filter=19 channel=86
    2, -5, 0, 6, 0, -7, -14, -13, 7,
    -- layer=1 filter=19 channel=87
    6, -5, -7, -2, -5, -4, -9, -6, -1,
    -- layer=1 filter=19 channel=88
    -13, -15, 2, -16, -1, -7, -15, 2, -8,
    -- layer=1 filter=19 channel=89
    -10, -9, -2, -3, -15, -4, 0, -5, 2,
    -- layer=1 filter=19 channel=90
    4, 8, -7, 0, -11, -3, -8, 2, -8,
    -- layer=1 filter=19 channel=91
    -5, -14, 0, -6, -5, 0, 0, -11, -13,
    -- layer=1 filter=19 channel=92
    7, -6, -4, -11, -12, 1, -2, -5, 1,
    -- layer=1 filter=19 channel=93
    -9, -11, -2, -10, -10, -12, 3, 2, 0,
    -- layer=1 filter=19 channel=94
    -1, -1, -2, -8, -4, 6, 1, -1, 0,
    -- layer=1 filter=19 channel=95
    2, 2, -10, -1, -10, -22, 2, -6, 0,
    -- layer=1 filter=19 channel=96
    2, -5, -2, -3, 6, 4, -10, -11, 6,
    -- layer=1 filter=19 channel=97
    5, 4, -5, -10, 2, -3, 2, 0, 0,
    -- layer=1 filter=19 channel=98
    -7, 1, -12, -9, -13, -14, 1, -13, -4,
    -- layer=1 filter=19 channel=99
    4, 7, -5, 3, -5, 0, 4, -8, -12,
    -- layer=1 filter=19 channel=100
    -6, 0, -5, 6, -9, 6, 4, 1, 4,
    -- layer=1 filter=19 channel=101
    3, -7, 6, 1, -3, -3, 4, 0, 5,
    -- layer=1 filter=19 channel=102
    -13, -11, -8, 5, 3, -10, 1, -8, 5,
    -- layer=1 filter=19 channel=103
    6, 0, 2, -6, 6, -9, -5, 6, -5,
    -- layer=1 filter=19 channel=104
    -12, 2, 0, -12, -3, -10, 7, 4, -7,
    -- layer=1 filter=19 channel=105
    -3, 4, -2, -13, 0, -8, -4, -12, 3,
    -- layer=1 filter=19 channel=106
    -3, -8, -8, 5, -3, 2, -8, -12, -10,
    -- layer=1 filter=19 channel=107
    -3, -1, 7, -6, 7, 8, -6, -6, -2,
    -- layer=1 filter=19 channel=108
    -2, -2, -10, -10, 13, -15, -7, -4, -11,
    -- layer=1 filter=19 channel=109
    -7, -4, 7, 1, -2, 6, -11, -7, 7,
    -- layer=1 filter=19 channel=110
    -8, 0, -13, -4, 0, -6, -1, -6, -1,
    -- layer=1 filter=19 channel=111
    -6, -5, -6, -9, 3, -7, -8, -7, -2,
    -- layer=1 filter=19 channel=112
    0, -2, 0, 2, -13, -3, 7, 6, -7,
    -- layer=1 filter=19 channel=113
    -2, 0, -2, 1, -10, -9, 1, -3, -4,
    -- layer=1 filter=19 channel=114
    -9, 0, -16, -3, -8, 5, -3, 7, -3,
    -- layer=1 filter=19 channel=115
    5, -3, -6, 2, -6, 1, -6, -8, -2,
    -- layer=1 filter=19 channel=116
    -8, 2, -9, -8, -9, 3, -3, 9, 2,
    -- layer=1 filter=19 channel=117
    -1, -2, -3, -3, 1, -15, -2, -11, 3,
    -- layer=1 filter=19 channel=118
    -5, -9, 0, -13, -2, -6, -7, -1, 3,
    -- layer=1 filter=19 channel=119
    1, -6, -4, -3, 14, -15, 5, 11, -9,
    -- layer=1 filter=19 channel=120
    -9, 1, -2, 2, 0, -5, -1, -2, 3,
    -- layer=1 filter=19 channel=121
    4, 10, 18, -12, 5, -17, 8, -9, -4,
    -- layer=1 filter=19 channel=122
    0, 10, 9, -6, 0, 1, 9, 1, 8,
    -- layer=1 filter=19 channel=123
    -9, -8, 0, -9, -16, 6, -3, 0, 7,
    -- layer=1 filter=19 channel=124
    -9, -3, 6, -9, -6, 2, -3, 8, -8,
    -- layer=1 filter=19 channel=125
    -4, -5, -1, 3, 2, 6, 6, 7, 1,
    -- layer=1 filter=19 channel=126
    4, 8, 0, 3, -2, -2, -9, -2, -7,
    -- layer=1 filter=19 channel=127
    9, -2, 9, -14, 0, -17, 8, 3, -2,
    -- layer=1 filter=20 channel=0
    -1, -3, 0, -19, -19, -10, -15, -3, -11,
    -- layer=1 filter=20 channel=1
    0, -13, 2, 0, -7, -12, -13, -15, -20,
    -- layer=1 filter=20 channel=2
    -16, -4, -20, -13, -3, -8, -12, -8, 1,
    -- layer=1 filter=20 channel=3
    7, 3, 9, 7, -3, -4, 9, 1, 7,
    -- layer=1 filter=20 channel=4
    -7, -1, -8, 1, -1, 6, 3, -10, 0,
    -- layer=1 filter=20 channel=5
    -12, -12, -7, -6, 5, -6, 0, -13, -8,
    -- layer=1 filter=20 channel=6
    -12, -17, -1, 0, 0, 3, -5, -14, -9,
    -- layer=1 filter=20 channel=7
    7, -14, 7, -7, -16, 3, -8, 3, -16,
    -- layer=1 filter=20 channel=8
    -2, 4, -5, 0, -1, 0, -12, -12, -19,
    -- layer=1 filter=20 channel=9
    -2, -2, -18, -3, -9, -3, -16, -5, -1,
    -- layer=1 filter=20 channel=10
    0, 3, 1, -9, -7, 0, -15, -6, 1,
    -- layer=1 filter=20 channel=11
    0, 0, -3, -17, -4, -4, -13, -14, -5,
    -- layer=1 filter=20 channel=12
    -2, -4, -1, -5, -5, -7, -10, 10, -10,
    -- layer=1 filter=20 channel=13
    -1, -2, -1, -9, -9, -17, -8, -3, -10,
    -- layer=1 filter=20 channel=14
    -4, -15, 3, 0, 0, 3, -4, 2, 3,
    -- layer=1 filter=20 channel=15
    0, 0, -1, 1, -8, -13, -6, 3, 0,
    -- layer=1 filter=20 channel=16
    7, -2, -1, 4, -7, -11, -15, -4, 0,
    -- layer=1 filter=20 channel=17
    -5, 0, -8, -15, -3, -16, -2, -13, -15,
    -- layer=1 filter=20 channel=18
    -8, -8, -8, -3, -2, -15, -5, -16, -13,
    -- layer=1 filter=20 channel=19
    -14, -22, -8, -11, 0, -3, -16, -15, -12,
    -- layer=1 filter=20 channel=20
    -16, 0, -9, -10, -22, -20, -16, -13, -11,
    -- layer=1 filter=20 channel=21
    -4, -12, -5, -11, -9, -8, 2, -19, -6,
    -- layer=1 filter=20 channel=22
    -2, -9, -9, -10, -2, -21, -1, -9, -10,
    -- layer=1 filter=20 channel=23
    -4, -1, -12, -10, -14, -3, 1, 0, -7,
    -- layer=1 filter=20 channel=24
    4, 0, -3, -7, 4, -8, -8, -7, -13,
    -- layer=1 filter=20 channel=25
    6, -4, 3, -6, -7, -9, -8, -9, -13,
    -- layer=1 filter=20 channel=26
    -8, 6, -6, -14, 5, -10, -21, -14, -6,
    -- layer=1 filter=20 channel=27
    -9, -8, -15, -3, -2, -13, -8, -6, -12,
    -- layer=1 filter=20 channel=28
    4, -4, -8, -13, 1, 2, -10, -18, -4,
    -- layer=1 filter=20 channel=29
    -16, 0, 0, 0, -7, -2, -12, 2, 4,
    -- layer=1 filter=20 channel=30
    -7, -7, -12, -5, -5, -6, -24, -5, -1,
    -- layer=1 filter=20 channel=31
    -11, -13, -4, 5, -10, -13, 0, -13, -10,
    -- layer=1 filter=20 channel=32
    -9, 0, -10, -7, 0, -6, -18, -4, 0,
    -- layer=1 filter=20 channel=33
    2, 1, 10, 7, 10, 2, -3, -5, -8,
    -- layer=1 filter=20 channel=34
    5, 3, -5, -16, 2, -7, -7, -12, -13,
    -- layer=1 filter=20 channel=35
    0, 0, -3, -4, -1, -3, 0, -1, -4,
    -- layer=1 filter=20 channel=36
    -9, -5, -4, -6, -16, -5, 3, -6, -6,
    -- layer=1 filter=20 channel=37
    7, 0, 4, 0, -13, -5, 4, -15, -7,
    -- layer=1 filter=20 channel=38
    -6, -13, -15, -8, 0, 0, -13, -8, -7,
    -- layer=1 filter=20 channel=39
    -10, -6, -4, -19, 0, -15, -9, -14, -17,
    -- layer=1 filter=20 channel=40
    -4, 1, -20, -11, 1, 0, -18, -7, -7,
    -- layer=1 filter=20 channel=41
    -4, 2, -8, -13, 1, 1, -6, 3, 2,
    -- layer=1 filter=20 channel=42
    -17, -10, -17, -16, -16, -8, -3, -3, -10,
    -- layer=1 filter=20 channel=43
    -8, -3, -2, -9, -7, 1, -15, -17, -1,
    -- layer=1 filter=20 channel=44
    -6, 1, -1, -8, 0, -5, -1, -7, 0,
    -- layer=1 filter=20 channel=45
    4, -7, -10, -15, 0, -6, -15, -8, -5,
    -- layer=1 filter=20 channel=46
    -11, 2, -10, -9, -18, -11, 4, -6, 0,
    -- layer=1 filter=20 channel=47
    -7, -7, -3, -16, 2, -18, -13, -4, -4,
    -- layer=1 filter=20 channel=48
    -8, -7, 0, -2, -14, -11, -11, -16, -9,
    -- layer=1 filter=20 channel=49
    -3, -5, -13, 1, 3, -11, -14, -16, 3,
    -- layer=1 filter=20 channel=50
    2, -10, 0, 4, -5, -5, -6, -8, 6,
    -- layer=1 filter=20 channel=51
    -3, -15, -13, -16, -7, 0, -11, -15, -6,
    -- layer=1 filter=20 channel=52
    -7, 0, -2, -7, 2, 0, -11, 1, -8,
    -- layer=1 filter=20 channel=53
    -7, -5, -3, -8, -1, -3, -6, -12, 4,
    -- layer=1 filter=20 channel=54
    7, -13, 7, 2, -8, -3, -17, -16, 4,
    -- layer=1 filter=20 channel=55
    0, 5, 0, -18, 3, -12, -9, -15, 0,
    -- layer=1 filter=20 channel=56
    5, 6, -12, -7, 5, -6, -11, -1, 6,
    -- layer=1 filter=20 channel=57
    -13, -11, -12, 0, -13, -9, -11, -10, -3,
    -- layer=1 filter=20 channel=58
    -5, -3, -1, 0, -9, -15, -1, -5, 2,
    -- layer=1 filter=20 channel=59
    -8, -10, 2, -4, 0, -3, 2, -1, -7,
    -- layer=1 filter=20 channel=60
    5, -3, -7, -9, -4, -5, 7, 7, 2,
    -- layer=1 filter=20 channel=61
    9, 3, -8, 7, 0, -5, -6, 10, -4,
    -- layer=1 filter=20 channel=62
    2, 3, -7, -4, -8, -1, -12, -19, -17,
    -- layer=1 filter=20 channel=63
    -2, 0, -10, 1, 2, 0, -18, -13, -11,
    -- layer=1 filter=20 channel=64
    -14, -18, -1, 0, -16, -15, 0, -13, -7,
    -- layer=1 filter=20 channel=65
    0, -11, 2, 1, -14, -7, -4, -17, -3,
    -- layer=1 filter=20 channel=66
    -11, -15, -6, -9, -11, -13, -15, -13, -1,
    -- layer=1 filter=20 channel=67
    6, -11, -5, -20, 0, -6, -13, -13, -3,
    -- layer=1 filter=20 channel=68
    -10, -11, -9, -15, -7, -4, -16, 0, -3,
    -- layer=1 filter=20 channel=69
    -12, 0, -3, 6, -6, -4, -5, -4, -13,
    -- layer=1 filter=20 channel=70
    -11, -18, -11, -9, -3, -5, -1, -4, 0,
    -- layer=1 filter=20 channel=71
    -8, 1, -13, -14, -6, -7, -3, -8, 3,
    -- layer=1 filter=20 channel=72
    -8, -4, -9, -7, -10, -16, -2, -11, -15,
    -- layer=1 filter=20 channel=73
    6, -5, 6, 0, -12, -9, -5, -6, -12,
    -- layer=1 filter=20 channel=74
    -6, -15, -10, -21, -14, -17, -15, -11, -13,
    -- layer=1 filter=20 channel=75
    -10, -8, 0, 2, -20, -11, -12, -5, -1,
    -- layer=1 filter=20 channel=76
    -4, 1, -17, -13, -3, -15, -10, -13, -14,
    -- layer=1 filter=20 channel=77
    -3, -7, -3, -18, -6, -11, -12, -12, -8,
    -- layer=1 filter=20 channel=78
    -1, -13, -1, -9, -1, -9, 0, -18, -12,
    -- layer=1 filter=20 channel=79
    -13, 7, 4, 2, -9, -10, -15, 1, -18,
    -- layer=1 filter=20 channel=80
    -9, -11, 5, 1, -4, -10, 1, 0, -6,
    -- layer=1 filter=20 channel=81
    -5, -11, 1, -18, -3, -11, -16, -5, -12,
    -- layer=1 filter=20 channel=82
    -2, -8, -2, -1, 0, -7, -2, 1, -2,
    -- layer=1 filter=20 channel=83
    -7, -6, -13, -3, -5, -17, -8, -7, -2,
    -- layer=1 filter=20 channel=84
    1, -10, -14, -16, -2, 3, -19, -12, -1,
    -- layer=1 filter=20 channel=85
    0, -21, -11, -13, -2, -3, -2, -7, -18,
    -- layer=1 filter=20 channel=86
    -12, -1, 7, -2, -14, -8, -14, -9, -9,
    -- layer=1 filter=20 channel=87
    0, 7, -2, -1, 2, -7, 3, -15, 0,
    -- layer=1 filter=20 channel=88
    -7, -10, -1, -2, -3, 8, 0, -18, -8,
    -- layer=1 filter=20 channel=89
    0, -14, -4, -8, -1, 0, -9, 0, -9,
    -- layer=1 filter=20 channel=90
    -17, 3, -8, -12, 1, -5, -12, -4, -10,
    -- layer=1 filter=20 channel=91
    2, -17, 0, 1, -12, -11, -21, 0, -8,
    -- layer=1 filter=20 channel=92
    0, 1, 0, -9, -7, -5, 2, 3, -1,
    -- layer=1 filter=20 channel=93
    -14, 3, -10, -8, -6, -2, -3, -8, -12,
    -- layer=1 filter=20 channel=94
    -10, -7, 1, -14, -17, -5, -14, -17, 0,
    -- layer=1 filter=20 channel=95
    -16, -8, 2, -4, 2, -8, -9, -3, -9,
    -- layer=1 filter=20 channel=96
    -6, -6, -2, -10, -17, 0, -13, -2, 4,
    -- layer=1 filter=20 channel=97
    -7, -3, -1, 2, -7, -5, -6, -2, -9,
    -- layer=1 filter=20 channel=98
    3, -11, 4, -15, -3, -7, -9, -19, -4,
    -- layer=1 filter=20 channel=99
    -1, -2, 4, -9, -5, -4, -4, -14, 0,
    -- layer=1 filter=20 channel=100
    -9, -13, 2, -8, -12, -1, -13, -1, 0,
    -- layer=1 filter=20 channel=101
    -15, -17, -6, -16, -7, -1, -2, -14, -9,
    -- layer=1 filter=20 channel=102
    -8, -2, -2, -17, -16, -18, -5, -9, -21,
    -- layer=1 filter=20 channel=103
    -20, -13, -13, -15, -8, -9, -9, 1, -4,
    -- layer=1 filter=20 channel=104
    -6, 2, -4, -2, -3, -15, -7, -21, -16,
    -- layer=1 filter=20 channel=105
    -1, -15, -16, -14, -18, 2, -11, -9, -1,
    -- layer=1 filter=20 channel=106
    -8, -8, -2, 0, -6, -18, -16, -9, -14,
    -- layer=1 filter=20 channel=107
    9, 0, 0, 1, -11, -2, 0, -2, -6,
    -- layer=1 filter=20 channel=108
    0, -1, -2, -4, 4, -17, -11, -8, 2,
    -- layer=1 filter=20 channel=109
    5, 10, 7, -4, 0, 0, 9, 0, 9,
    -- layer=1 filter=20 channel=110
    -11, -13, 3, 1, -16, -15, -5, -20, -14,
    -- layer=1 filter=20 channel=111
    -17, -11, 3, -3, -11, -7, -22, -3, -17,
    -- layer=1 filter=20 channel=112
    -13, -11, -4, 1, -14, -4, -15, 0, -21,
    -- layer=1 filter=20 channel=113
    -7, -7, 1, -7, -3, 3, -1, -9, -9,
    -- layer=1 filter=20 channel=114
    -13, -6, -7, -13, -1, -15, 0, -12, -12,
    -- layer=1 filter=20 channel=115
    -4, -12, 0, -16, -10, -1, -15, -12, -12,
    -- layer=1 filter=20 channel=116
    2, 6, -7, -3, 3, -2, -3, -10, -9,
    -- layer=1 filter=20 channel=117
    -8, 2, -1, 2, -14, -15, -10, -18, -17,
    -- layer=1 filter=20 channel=118
    0, -16, -9, -16, 5, -15, -10, -14, 0,
    -- layer=1 filter=20 channel=119
    -8, -7, 0, -6, -14, -3, -2, -10, -4,
    -- layer=1 filter=20 channel=120
    1, -14, 2, -4, -15, -13, -1, -17, 4,
    -- layer=1 filter=20 channel=121
    -1, -12, -8, -15, -16, -10, -14, 0, -3,
    -- layer=1 filter=20 channel=122
    4, -2, 9, 0, -8, 1, 3, -7, -9,
    -- layer=1 filter=20 channel=123
    -4, -4, -12, -6, 3, -2, -6, -1, -16,
    -- layer=1 filter=20 channel=124
    0, 6, 2, -5, -3, -10, -1, -4, 0,
    -- layer=1 filter=20 channel=125
    -2, -14, -11, 0, 4, 5, -18, -8, -9,
    -- layer=1 filter=20 channel=126
    3, 5, -9, -8, -11, -1, 0, -12, -19,
    -- layer=1 filter=20 channel=127
    -3, 0, 4, 4, -7, 0, -8, -1, -15,
    -- layer=1 filter=21 channel=0
    -25, -34, -34, -7, -21, -32, -29, -35, -11,
    -- layer=1 filter=21 channel=1
    -35, -16, -30, -33, -11, -23, -51, -33, -11,
    -- layer=1 filter=21 channel=2
    31, 16, -5, 23, 26, -42, 22, 40, -3,
    -- layer=1 filter=21 channel=3
    8, -8, 4, -5, 0, -6, 6, 0, -1,
    -- layer=1 filter=21 channel=4
    -2, -15, 2, 6, 4, -4, -7, 8, -8,
    -- layer=1 filter=21 channel=5
    -24, -10, 14, -12, -18, 25, -41, -40, -17,
    -- layer=1 filter=21 channel=6
    -6, 15, 0, 3, 9, -12, -11, -17, 0,
    -- layer=1 filter=21 channel=7
    8, -31, -13, -1, -27, 47, 32, -34, 78,
    -- layer=1 filter=21 channel=8
    -28, -17, 14, -31, -30, 20, -57, -65, -36,
    -- layer=1 filter=21 channel=9
    6, -27, -9, -4, 24, 32, 10, 22, 29,
    -- layer=1 filter=21 channel=10
    11, -11, -12, 4, -14, 60, 18, -46, 76,
    -- layer=1 filter=21 channel=11
    -43, -62, -61, -36, -28, -67, -22, 11, -37,
    -- layer=1 filter=21 channel=12
    13, 11, 0, 25, 21, -17, 15, 31, 41,
    -- layer=1 filter=21 channel=13
    -3, -8, 25, -15, -19, -4, -21, -1, -31,
    -- layer=1 filter=21 channel=14
    14, -13, -8, 17, -18, 3, 25, 3, 105,
    -- layer=1 filter=21 channel=15
    32, 18, 21, -12, 18, -28, -2, 0, -24,
    -- layer=1 filter=21 channel=16
    -11, -17, 35, -17, -37, 51, -44, -74, -11,
    -- layer=1 filter=21 channel=17
    -7, 0, -26, -47, -11, 5, -26, -10, -36,
    -- layer=1 filter=21 channel=18
    -58, -65, -20, -23, -41, -78, -24, -19, 18,
    -- layer=1 filter=21 channel=19
    -21, -52, 30, -38, -30, 29, -37, -65, 7,
    -- layer=1 filter=21 channel=20
    -3, 9, 9, -13, -4, 35, -33, -18, 8,
    -- layer=1 filter=21 channel=21
    -11, -21, -30, 2, -18, -9, -20, -21, 14,
    -- layer=1 filter=21 channel=22
    27, 23, 16, -13, 8, 30, -4, 1, 5,
    -- layer=1 filter=21 channel=23
    -15, -36, 4, -44, -13, 53, 31, -23, 47,
    -- layer=1 filter=21 channel=24
    -1, -22, 44, -6, -19, 0, -17, 4, -75,
    -- layer=1 filter=21 channel=25
    -3, -28, -10, 0, -43, 54, 11, -55, 72,
    -- layer=1 filter=21 channel=26
    -3, -27, 0, -34, -13, -22, -6, 15, -30,
    -- layer=1 filter=21 channel=27
    1, 3, -6, 26, -10, -24, 32, 8, 29,
    -- layer=1 filter=21 channel=28
    -2, -23, -29, -9, -26, 34, -14, -45, 54,
    -- layer=1 filter=21 channel=29
    -4, -15, -9, -50, -46, -5, -42, -47, 27,
    -- layer=1 filter=21 channel=30
    -31, -52, -19, -34, -34, -71, -34, -17, 22,
    -- layer=1 filter=21 channel=31
    3, 15, 13, 22, 10, -18, 35, 34, 47,
    -- layer=1 filter=21 channel=32
    -18, -26, -37, -43, -13, -18, -17, 0, -37,
    -- layer=1 filter=21 channel=33
    22, 18, -30, 24, 15, -16, 18, 23, -28,
    -- layer=1 filter=21 channel=34
    -17, -19, -14, -4, -11, -12, -2, 14, -19,
    -- layer=1 filter=21 channel=35
    2, 0, 6, 7, -3, -4, -1, -11, 0,
    -- layer=1 filter=21 channel=36
    -57, -71, -78, -34, -58, -85, -42, -19, -33,
    -- layer=1 filter=21 channel=37
    -3, -19, 20, -11, -41, 42, -42, -63, -8,
    -- layer=1 filter=21 channel=38
    -7, 8, 15, -9, -11, 28, -13, -16, 26,
    -- layer=1 filter=21 channel=39
    -16, -21, -2, -35, -25, -18, 0, -40, -28,
    -- layer=1 filter=21 channel=40
    4, 11, 8, -2, 14, 23, -23, 10, 72,
    -- layer=1 filter=21 channel=41
    -24, -28, 0, -50, 6, 0, -3, 36, -20,
    -- layer=1 filter=21 channel=42
    33, 24, 24, 9, 13, -5, 24, 27, 27,
    -- layer=1 filter=21 channel=43
    -3, -20, 14, -2, -16, 54, -36, -45, 37,
    -- layer=1 filter=21 channel=44
    -24, -41, -36, -38, -20, -32, -15, 3, -23,
    -- layer=1 filter=21 channel=45
    -9, -35, 0, -17, -4, -2, -37, -2, -49,
    -- layer=1 filter=21 channel=46
    -26, -17, 37, -26, -9, -11, -2, -27, 14,
    -- layer=1 filter=21 channel=47
    14, 6, 18, -35, 11, 29, 32, 0, 10,
    -- layer=1 filter=21 channel=48
    -56, -23, -3, -32, -46, 47, -37, -49, 43,
    -- layer=1 filter=21 channel=49
    -9, -5, -9, -7, 26, -32, 4, 26, -36,
    -- layer=1 filter=21 channel=50
    1, -15, 0, -10, -1, -18, -2, 9, 5,
    -- layer=1 filter=21 channel=51
    -16, -15, -19, -9, -5, 35, -16, -26, 53,
    -- layer=1 filter=21 channel=52
    6, 4, -4, -30, -10, -25, 32, 17, 9,
    -- layer=1 filter=21 channel=53
    3, 4, 0, -7, 4, 13, 6, 9, 2,
    -- layer=1 filter=21 channel=54
    1, -23, 19, -1, -23, 71, 20, -42, 62,
    -- layer=1 filter=21 channel=55
    -7, 4, -13, -16, 0, -59, -10, -2, -76,
    -- layer=1 filter=21 channel=56
    0, -6, -5, 5, 6, 2, -1, 0, 6,
    -- layer=1 filter=21 channel=57
    -10, -1, -19, 11, -9, 44, 12, -28, 57,
    -- layer=1 filter=21 channel=58
    9, -32, 3, -3, -21, 70, 54, -34, 61,
    -- layer=1 filter=21 channel=59
    -3, 5, 0, 2, 5, 5, 0, -3, -3,
    -- layer=1 filter=21 channel=60
    13, 30, -14, 8, 0, -24, 20, 37, 0,
    -- layer=1 filter=21 channel=61
    2, 9, -4, -4, 1, 0, 3, 8, -4,
    -- layer=1 filter=21 channel=62
    -16, -16, 41, -21, -38, 65, -26, -75, -4,
    -- layer=1 filter=21 channel=63
    -56, -75, -64, -56, -51, -72, -17, -9, -30,
    -- layer=1 filter=21 channel=64
    7, -6, -8, 0, 10, 3, -4, -6, 5,
    -- layer=1 filter=21 channel=65
    -46, -25, -23, -46, -32, 16, -35, -35, 26,
    -- layer=1 filter=21 channel=66
    -47, -39, -49, -31, -39, -31, 1, -13, -27,
    -- layer=1 filter=21 channel=67
    -51, -32, -27, 9, -28, -24, -23, -30, -14,
    -- layer=1 filter=21 channel=68
    -5, -34, -30, -19, -24, -27, -12, 16, -62,
    -- layer=1 filter=21 channel=69
    -5, -4, 53, -15, -7, 8, -24, -28, -57,
    -- layer=1 filter=21 channel=70
    -5, -6, -13, 18, 10, -13, 28, 22, 54,
    -- layer=1 filter=21 channel=71
    -16, -28, -4, 0, -23, 4, -13, -27, 22,
    -- layer=1 filter=21 channel=72
    -34, -70, 4, -32, -22, -33, -43, -30, -6,
    -- layer=1 filter=21 channel=73
    -5, 7, 0, 6, -10, 7, -8, -10, 7,
    -- layer=1 filter=21 channel=74
    -21, -35, -8, 14, 8, 4, -20, 15, -26,
    -- layer=1 filter=21 channel=75
    14, -26, 41, 1, -16, -31, 36, 20, 55,
    -- layer=1 filter=21 channel=76
    -42, -38, -61, -46, -23, 14, -28, 7, -27,
    -- layer=1 filter=21 channel=77
    -22, -32, -19, 6, -20, -4, -18, -28, 0,
    -- layer=1 filter=21 channel=78
    -11, 5, -33, -14, -4, 18, -19, 0, 19,
    -- layer=1 filter=21 channel=79
    -6, -35, 49, -15, -31, 56, -33, -72, -12,
    -- layer=1 filter=21 channel=80
    0, 12, 9, 3, 24, 29, -20, -8, 13,
    -- layer=1 filter=21 channel=81
    -17, -29, 2, -7, -18, 27, -18, -40, -20,
    -- layer=1 filter=21 channel=82
    -50, -39, -26, -32, -36, -4, -22, -35, 3,
    -- layer=1 filter=21 channel=83
    17, -30, -1, -20, -18, -3, -27, -3, -22,
    -- layer=1 filter=21 channel=84
    -44, -59, -14, -43, -12, -36, -48, -1, -23,
    -- layer=1 filter=21 channel=85
    7, -41, 27, -15, -8, 57, 32, 6, 58,
    -- layer=1 filter=21 channel=86
    -16, -24, -20, -38, -14, -24, -22, -24, -4,
    -- layer=1 filter=21 channel=87
    14, -38, 26, -30, 10, -14, -5, -23, -16,
    -- layer=1 filter=21 channel=88
    -11, -14, 7, 10, 1, -17, -9, 7, -34,
    -- layer=1 filter=21 channel=89
    -55, -39, -34, -50, -29, -47, -58, -41, -27,
    -- layer=1 filter=21 channel=90
    -3, -40, -30, -18, -22, -16, -13, -3, -24,
    -- layer=1 filter=21 channel=91
    -17, 1, 6, -11, -3, 10, -16, -18, 45,
    -- layer=1 filter=21 channel=92
    -8, 22, -21, -13, 21, 0, 0, 26, 21,
    -- layer=1 filter=21 channel=93
    -41, -37, -23, -10, -21, 9, -38, -31, 12,
    -- layer=1 filter=21 channel=94
    -28, -33, -44, -13, -30, -35, -18, -28, 15,
    -- layer=1 filter=21 channel=95
    -45, -57, 3, -36, -42, -76, -29, -21, 3,
    -- layer=1 filter=21 channel=96
    -5, 7, 10, 8, 6, -2, 38, 38, 41,
    -- layer=1 filter=21 channel=97
    -48, -48, -41, -54, -26, -22, -44, -47, -24,
    -- layer=1 filter=21 channel=98
    -7, -21, 22, -27, -21, 78, -20, -53, 19,
    -- layer=1 filter=21 channel=99
    -7, 26, -40, -3, 12, 13, -51, -10, 37,
    -- layer=1 filter=21 channel=100
    -71, -80, -35, -62, -47, -13, -18, -3, -14,
    -- layer=1 filter=21 channel=101
    -24, -23, -14, -14, -9, 1, -32, -11, 21,
    -- layer=1 filter=21 channel=102
    -22, -6, -16, -18, -12, -34, -44, -25, -12,
    -- layer=1 filter=21 channel=103
    -44, -46, -44, 6, -24, -30, -17, 22, -27,
    -- layer=1 filter=21 channel=104
    -18, -28, 2, -43, 11, 69, 0, 22, 73,
    -- layer=1 filter=21 channel=105
    -40, -26, -41, -21, -32, -8, -18, -50, 13,
    -- layer=1 filter=21 channel=106
    -1, -11, -17, -13, -5, -14, -23, 11, -39,
    -- layer=1 filter=21 channel=107
    -1, 7, -8, -2, 7, -11, -9, 0, -5,
    -- layer=1 filter=21 channel=108
    -15, -43, -29, -48, -4, -25, -27, 16, -30,
    -- layer=1 filter=21 channel=109
    4, 4, -4, -9, 6, 5, -8, -9, -5,
    -- layer=1 filter=21 channel=110
    -8, 13, 24, -13, -7, 0, -4, -10, 39,
    -- layer=1 filter=21 channel=111
    -53, -50, -19, -23, -9, -37, -36, -32, 11,
    -- layer=1 filter=21 channel=112
    -27, -15, -8, -14, -3, 6, -8, -18, -2,
    -- layer=1 filter=21 channel=113
    11, 5, 43, 16, 16, 45, 28, 20, 69,
    -- layer=1 filter=21 channel=114
    -32, 1, 39, -41, -24, 4, -49, -52, -78,
    -- layer=1 filter=21 channel=115
    -4, -17, -24, -18, -19, 36, 0, -63, 45,
    -- layer=1 filter=21 channel=116
    -4, 0, 1, 1, 9, -2, -9, 7, 2,
    -- layer=1 filter=21 channel=117
    -21, -2, -13, 30, 14, 65, -31, -41, 44,
    -- layer=1 filter=21 channel=118
    -48, -37, -19, -22, -27, -17, -42, 0, -6,
    -- layer=1 filter=21 channel=119
    -18, -51, -27, -52, -20, -17, -32, 2, -47,
    -- layer=1 filter=21 channel=120
    -25, -27, -18, 7, -18, 39, -15, -43, 33,
    -- layer=1 filter=21 channel=121
    -7, -42, -15, -27, -24, -89, 7, 0, 14,
    -- layer=1 filter=21 channel=122
    8, 4, 6, -2, 6, 2, -8, -1, -4,
    -- layer=1 filter=21 channel=123
    -5, -29, -12, -17, -7, -52, 17, -5, 19,
    -- layer=1 filter=21 channel=124
    0, 24, 9, 8, -7, -2, -10, 17, 0,
    -- layer=1 filter=21 channel=125
    -29, -5, -18, 15, 30, 73, 10, 11, 66,
    -- layer=1 filter=21 channel=126
    -11, -15, 1, -37, -17, 30, -31, -53, -14,
    -- layer=1 filter=21 channel=127
    -36, -43, -18, -46, -40, -56, -28, -5, 4,
    -- layer=1 filter=22 channel=0
    32, -18, -54, 40, 5, -48, 23, 5, -21,
    -- layer=1 filter=22 channel=1
    14, 13, -18, -16, -15, -11, -39, 3, 17,
    -- layer=1 filter=22 channel=2
    -44, -19, 27, -11, 33, 42, 6, 2, 55,
    -- layer=1 filter=22 channel=3
    -2, 0, 4, -1, 1, 10, -9, 1, 5,
    -- layer=1 filter=22 channel=4
    0, -9, -19, 12, -12, -13, -4, -8, -5,
    -- layer=1 filter=22 channel=5
    12, 26, -32, 1, -6, -4, -29, 9, 30,
    -- layer=1 filter=22 channel=6
    -75, 8, 52, -77, -11, 52, -11, 5, 35,
    -- layer=1 filter=22 channel=7
    -42, -49, 10, -55, -77, -21, -29, -72, -60,
    -- layer=1 filter=22 channel=8
    19, 26, -10, -9, -18, 0, -12, 30, 15,
    -- layer=1 filter=22 channel=9
    -17, -20, -6, -24, -12, -14, -15, -18, -10,
    -- layer=1 filter=22 channel=10
    -51, -71, -22, -72, -83, -32, -50, -44, -68,
    -- layer=1 filter=22 channel=11
    46, -4, -50, 59, -1, -52, 70, 3, -21,
    -- layer=1 filter=22 channel=12
    -4, -47, -10, -38, 2, 56, -12, 11, 13,
    -- layer=1 filter=22 channel=13
    6, 6, 26, -20, 14, 27, -24, 19, 13,
    -- layer=1 filter=22 channel=14
    -34, -15, 8, -38, -2, 36, -84, -57, -25,
    -- layer=1 filter=22 channel=15
    19, 31, 16, 16, 6, 24, -51, 46, 43,
    -- layer=1 filter=22 channel=16
    6, -3, -14, 0, -22, -13, -14, -4, -3,
    -- layer=1 filter=22 channel=17
    23, -18, -34, 31, 16, -36, 35, 25, -20,
    -- layer=1 filter=22 channel=18
    5, 21, 8, 1, -29, -9, 4, 0, -20,
    -- layer=1 filter=22 channel=19
    -73, -56, -38, -64, -70, -39, -25, -66, -77,
    -- layer=1 filter=22 channel=20
    9, 20, 27, -8, 6, 18, -11, 5, 5,
    -- layer=1 filter=22 channel=21
    -26, -1, 20, -29, -10, 22, -41, -13, 25,
    -- layer=1 filter=22 channel=22
    -18, 8, 8, -23, -4, 13, -20, 0, 9,
    -- layer=1 filter=22 channel=23
    -20, 8, -41, -33, -11, -34, 23, -25, -39,
    -- layer=1 filter=22 channel=24
    14, 20, 21, 1, 32, 25, -6, 26, 17,
    -- layer=1 filter=22 channel=25
    -56, -77, -21, -74, -98, -49, -38, -74, -63,
    -- layer=1 filter=22 channel=26
    21, 19, 7, 25, 28, 21, -6, 20, 16,
    -- layer=1 filter=22 channel=27
    12, -7, -42, 34, 8, -49, 25, 0, -12,
    -- layer=1 filter=22 channel=28
    -30, -83, -6, -40, -100, -55, -17, -59, -77,
    -- layer=1 filter=22 channel=29
    27, -1, -29, 20, -1, -18, 0, -11, -25,
    -- layer=1 filter=22 channel=30
    -40, -21, 18, 2, -50, 5, -6, -31, -39,
    -- layer=1 filter=22 channel=31
    -15, -19, 10, -38, -17, 30, 3, 18, 25,
    -- layer=1 filter=22 channel=32
    30, 27, 20, 36, 33, 29, 13, 20, 21,
    -- layer=1 filter=22 channel=33
    -14, 14, 45, -43, 5, 29, -22, -9, 44,
    -- layer=1 filter=22 channel=34
    -17, -5, 48, -21, -23, 28, -9, -7, 24,
    -- layer=1 filter=22 channel=35
    1, 0, -8, 3, -10, 10, -1, -10, 11,
    -- layer=1 filter=22 channel=36
    55, -5, -47, 71, 0, -66, 77, 22, -37,
    -- layer=1 filter=22 channel=37
    15, -2, -22, -11, -19, 0, -13, 9, 20,
    -- layer=1 filter=22 channel=38
    -6, 19, 38, -27, -1, 30, -24, 7, 9,
    -- layer=1 filter=22 channel=39
    5, -13, -54, 27, -22, -60, 19, 15, -19,
    -- layer=1 filter=22 channel=40
    -61, -21, 42, -62, -48, 38, -14, -6, 33,
    -- layer=1 filter=22 channel=41
    27, -31, 0, -15, -22, -45, 4, -37, -22,
    -- layer=1 filter=22 channel=42
    -31, -5, 3, -42, -1, 49, -50, 0, 27,
    -- layer=1 filter=22 channel=43
    -15, -24, -25, -20, -40, -40, -13, -22, -17,
    -- layer=1 filter=22 channel=44
    52, 34, 5, 31, 48, 10, 3, 39, 8,
    -- layer=1 filter=22 channel=45
    21, 15, 26, 8, 28, 20, -34, 13, 17,
    -- layer=1 filter=22 channel=46
    -65, -4, 13, 0, 16, 19, -52, -19, -1,
    -- layer=1 filter=22 channel=47
    -26, -12, 2, -49, -58, 6, -32, -38, 8,
    -- layer=1 filter=22 channel=48
    -39, -3, 20, -23, -14, 38, -6, -17, 8,
    -- layer=1 filter=22 channel=49
    -37, -10, 40, -67, -23, 27, -33, -17, 34,
    -- layer=1 filter=22 channel=50
    -5, -14, -10, -14, -3, -18, 5, -5, 3,
    -- layer=1 filter=22 channel=51
    -50, -14, 15, -54, -25, 18, -16, -28, -4,
    -- layer=1 filter=22 channel=52
    -9, -6, -9, 19, -10, -14, 20, -14, 10,
    -- layer=1 filter=22 channel=53
    -13, -9, -10, 0, 9, -7, -7, -22, -5,
    -- layer=1 filter=22 channel=54
    -72, -45, -37, -66, -85, -55, -36, -50, -69,
    -- layer=1 filter=22 channel=55
    35, -15, -42, 54, -13, -27, 59, 12, -7,
    -- layer=1 filter=22 channel=56
    6, -6, 5, 2, 3, -7, 8, 7, -8,
    -- layer=1 filter=22 channel=57
    -59, -49, 4, -68, -95, -24, -54, -45, -50,
    -- layer=1 filter=22 channel=58
    -137, -51, -53, -114, -119, -49, -34, -67, -90,
    -- layer=1 filter=22 channel=59
    34, 15, -28, 6, 7, 2, -16, 7, 19,
    -- layer=1 filter=22 channel=60
    17, -6, -41, -1, 21, 6, 30, 5, 5,
    -- layer=1 filter=22 channel=61
    -1, -10, 1, 8, -6, 0, -4, 8, -2,
    -- layer=1 filter=22 channel=62
    18, 28, -18, -10, -2, -6, -12, 21, 0,
    -- layer=1 filter=22 channel=63
    43, -2, -33, 53, -14, -60, 46, 6, -22,
    -- layer=1 filter=22 channel=64
    -6, 4, 13, -27, 1, -2, -13, -3, -3,
    -- layer=1 filter=22 channel=65
    -14, 0, 25, -11, -5, 20, -17, -9, 5,
    -- layer=1 filter=22 channel=66
    32, -15, -55, 40, 0, -53, 53, 6, -20,
    -- layer=1 filter=22 channel=67
    -60, -12, 46, -62, 14, 74, -33, 1, 55,
    -- layer=1 filter=22 channel=68
    70, 14, 0, 44, 53, 15, 23, 52, 12,
    -- layer=1 filter=22 channel=69
    18, 37, 25, -1, 14, 19, -45, 16, 28,
    -- layer=1 filter=22 channel=70
    -33, 11, 44, -65, -6, 40, -47, -2, 55,
    -- layer=1 filter=22 channel=71
    -9, 7, 5, -16, 17, 8, -3, 2, 3,
    -- layer=1 filter=22 channel=72
    -40, -19, -2, -28, -59, -21, -9, -21, -41,
    -- layer=1 filter=22 channel=73
    10, -6, -4, 7, 16, -9, -1, 9, -14,
    -- layer=1 filter=22 channel=74
    -3, -5, -5, 14, -13, -28, 16, -7, -62,
    -- layer=1 filter=22 channel=75
    -43, -21, 11, -45, -14, 72, -37, -19, 5,
    -- layer=1 filter=22 channel=76
    18, 10, -13, 28, 7, -25, 23, -2, -38,
    -- layer=1 filter=22 channel=77
    -8, -24, 9, -11, -11, 0, -13, 4, 1,
    -- layer=1 filter=22 channel=78
    0, -42, -24, 2, -36, -51, 6, -1, -31,
    -- layer=1 filter=22 channel=79
    -6, 27, 6, -12, 0, 13, -22, 20, 17,
    -- layer=1 filter=22 channel=80
    18, 1, -31, 8, 3, 7, -3, 6, 22,
    -- layer=1 filter=22 channel=81
    -16, -23, -5, 11, -32, -3, 21, 16, 6,
    -- layer=1 filter=22 channel=82
    -35, 4, 36, -42, 2, 42, -41, 0, 37,
    -- layer=1 filter=22 channel=83
    37, 2, -21, 14, 5, 1, -24, 18, 13,
    -- layer=1 filter=22 channel=84
    9, 26, 2, 27, 3, 6, 43, -1, -16,
    -- layer=1 filter=22 channel=85
    -54, -32, -12, -62, -33, -5, -20, -35, -43,
    -- layer=1 filter=22 channel=86
    36, 0, -48, 53, 0, -42, 46, 0, -37,
    -- layer=1 filter=22 channel=87
    -14, -47, -31, -1, -34, -13, -14, 20, -3,
    -- layer=1 filter=22 channel=88
    -38, 1, 28, -50, -1, 40, -38, -13, 16,
    -- layer=1 filter=22 channel=89
    -17, 14, 34, -35, 9, 29, -29, -9, 22,
    -- layer=1 filter=22 channel=90
    65, 36, 22, 48, 56, 25, 12, 40, 26,
    -- layer=1 filter=22 channel=91
    -23, -1, 27, -35, -4, 36, -25, -13, 11,
    -- layer=1 filter=22 channel=92
    2, -27, -9, 3, -32, 4, -29, -9, 6,
    -- layer=1 filter=22 channel=93
    9, 9, -2, 3, 2, 15, -6, 4, 10,
    -- layer=1 filter=22 channel=94
    22, -12, -47, 26, -21, -64, 30, -1, -51,
    -- layer=1 filter=22 channel=95
    10, 15, 18, 10, -7, 12, 30, -20, -43,
    -- layer=1 filter=22 channel=96
    17, -3, -26, 1, -29, -17, 2, -6, -7,
    -- layer=1 filter=22 channel=97
    31, -12, -17, 36, 0, -25, 22, 12, -5,
    -- layer=1 filter=22 channel=98
    -4, -21, -6, -32, -18, -11, -11, 4, 0,
    -- layer=1 filter=22 channel=99
    -13, -96, -80, -43, -65, -105, -13, -43, -108,
    -- layer=1 filter=22 channel=100
    42, -6, -38, 58, 1, -58, 59, 26, -26,
    -- layer=1 filter=22 channel=101
    -2, 14, 25, -11, 0, 18, -16, -3, 15,
    -- layer=1 filter=22 channel=102
    13, -10, -24, 11, -3, -28, 13, -4, -33,
    -- layer=1 filter=22 channel=103
    32, -5, -19, 32, 15, -39, 47, 17, -14,
    -- layer=1 filter=22 channel=104
    -20, -10, 15, -16, 9, 11, 13, -5, -4,
    -- layer=1 filter=22 channel=105
    27, -9, -33, 44, -3, -38, 37, 2, -33,
    -- layer=1 filter=22 channel=106
    8, 17, 37, 0, 22, 37, -19, 20, 21,
    -- layer=1 filter=22 channel=107
    5, 8, 18, -2, -2, 16, 9, 15, 6,
    -- layer=1 filter=22 channel=108
    44, 48, 37, 41, 63, 45, 0, 66, 42,
    -- layer=1 filter=22 channel=109
    -6, -4, 5, 10, -3, 9, 9, 5, 2,
    -- layer=1 filter=22 channel=110
    9, -10, -20, 5, -19, -26, 0, -3, -18,
    -- layer=1 filter=22 channel=111
    -9, 24, 21, 16, -37, 12, 4, -6, -37,
    -- layer=1 filter=22 channel=112
    -1, 14, -11, 7, -4, -4, -7, -15, -29,
    -- layer=1 filter=22 channel=113
    -30, -13, 17, -80, -50, 14, -60, -30, 17,
    -- layer=1 filter=22 channel=114
    5, 0, -36, 38, -26, -29, 3, 19, 19,
    -- layer=1 filter=22 channel=115
    25, -31, -60, 27, -20, -53, 34, 1, -34,
    -- layer=1 filter=22 channel=116
    6, 0, 9, 7, 9, -9, 6, -8, -6,
    -- layer=1 filter=22 channel=117
    10, -15, 7, -14, 4, 2, -38, -58, 5,
    -- layer=1 filter=22 channel=118
    14, 14, 16, 23, -8, -5, 22, -7, -18,
    -- layer=1 filter=22 channel=119
    52, 29, 37, 37, 43, 21, 21, 49, 33,
    -- layer=1 filter=22 channel=120
    -55, -13, 32, -43, -35, 34, -15, -23, 12,
    -- layer=1 filter=22 channel=121
    10, -11, -24, 1, 1, 0, 2, -18, -6,
    -- layer=1 filter=22 channel=122
    -8, 9, -2, 5, -2, 10, 2, 4, 6,
    -- layer=1 filter=22 channel=123
    26, -11, -9, 26, 0, -35, 34, 9, -21,
    -- layer=1 filter=22 channel=124
    5, 5, -2, 4, 0, 6, 3, 1, 2,
    -- layer=1 filter=22 channel=125
    -51, -4, 23, -96, -48, 26, -65, -42, 41,
    -- layer=1 filter=22 channel=126
    3, -38, -55, -38, -19, -9, -14, 24, 37,
    -- layer=1 filter=22 channel=127
    -8, 4, 15, 13, -15, -2, 13, -7, -36,
    -- layer=1 filter=23 channel=0
    16, -5, 1, -1, -2, 14, 3, 11, -8,
    -- layer=1 filter=23 channel=1
    1, -5, -13, -2, -6, 1, 18, -13, 5,
    -- layer=1 filter=23 channel=2
    11, 2, 13, -8, 18, 3, -8, 3, -6,
    -- layer=1 filter=23 channel=3
    -11, -3, -2, -11, 8, -8, -6, -7, -1,
    -- layer=1 filter=23 channel=4
    -4, 0, 2, -2, 2, 7, -9, -6, 0,
    -- layer=1 filter=23 channel=5
    -5, -18, -21, -7, -23, 0, 12, -20, 15,
    -- layer=1 filter=23 channel=6
    -25, -28, -4, -17, -24, -14, -38, -19, -9,
    -- layer=1 filter=23 channel=7
    -13, 0, -11, -4, 6, -1, 5, 6, 0,
    -- layer=1 filter=23 channel=8
    -4, -23, -19, -8, -10, 8, 4, -9, 13,
    -- layer=1 filter=23 channel=9
    7, -1, 31, -12, 1, -16, 3, -8, -1,
    -- layer=1 filter=23 channel=10
    -12, 9, -12, -3, -10, -17, 13, -3, -28,
    -- layer=1 filter=23 channel=11
    -30, -16, -6, -11, -8, -23, -14, -24, -19,
    -- layer=1 filter=23 channel=12
    20, 1, -13, -53, -47, -25, -8, -47, 14,
    -- layer=1 filter=23 channel=13
    2, 0, -9, 11, 1, -6, 11, 6, 3,
    -- layer=1 filter=23 channel=14
    -19, 21, -7, -26, -31, -31, 16, -35, -9,
    -- layer=1 filter=23 channel=15
    16, -6, -18, 14, -23, 17, 7, -7, 0,
    -- layer=1 filter=23 channel=16
    2, -13, -25, 7, 0, 7, -4, -11, 16,
    -- layer=1 filter=23 channel=17
    11, 1, 2, 6, 4, 0, -3, -6, -9,
    -- layer=1 filter=23 channel=18
    -23, -15, -16, -6, -22, -13, -42, -40, 1,
    -- layer=1 filter=23 channel=19
    -12, -21, -17, 21, 0, 14, 24, 35, 15,
    -- layer=1 filter=23 channel=20
    5, -12, -14, 12, 8, 12, 11, 15, 19,
    -- layer=1 filter=23 channel=21
    2, -2, 8, -14, 13, 8, -3, 6, 2,
    -- layer=1 filter=23 channel=22
    -18, -6, 0, -6, -3, 4, 0, 8, -2,
    -- layer=1 filter=23 channel=23
    19, -31, -13, -8, -33, 15, 26, -2, 7,
    -- layer=1 filter=23 channel=24
    5, 3, -5, -1, 11, 4, 2, -2, -4,
    -- layer=1 filter=23 channel=25
    -24, -12, -13, -3, -13, -18, 7, -5, -9,
    -- layer=1 filter=23 channel=26
    -2, 0, -12, 10, -5, -2, 8, 1, 1,
    -- layer=1 filter=23 channel=27
    13, 20, 11, 0, 0, -4, -24, -11, -33,
    -- layer=1 filter=23 channel=28
    -13, 9, -8, -22, -3, -4, 5, 10, -7,
    -- layer=1 filter=23 channel=29
    -2, 1, 20, -5, 0, 5, -7, -1, -16,
    -- layer=1 filter=23 channel=30
    -16, -11, -12, 10, -8, -7, -3, -1, 5,
    -- layer=1 filter=23 channel=31
    -15, 2, -4, -20, -19, -25, -20, -20, -3,
    -- layer=1 filter=23 channel=32
    5, 6, 8, -3, 3, -13, 8, 2, 0,
    -- layer=1 filter=23 channel=33
    -6, -14, -11, -8, -5, -5, -13, -14, -9,
    -- layer=1 filter=23 channel=34
    -25, -29, 13, -26, -4, 4, -25, -27, -9,
    -- layer=1 filter=23 channel=35
    18, 17, 7, 18, 15, 16, 16, 15, 7,
    -- layer=1 filter=23 channel=36
    -32, -7, -24, -19, -29, -26, -28, -19, -28,
    -- layer=1 filter=23 channel=37
    -16, -9, -24, 0, -22, -13, 3, -11, -11,
    -- layer=1 filter=23 channel=38
    2, -7, -4, 9, 4, 7, 15, 12, 11,
    -- layer=1 filter=23 channel=39
    0, 4, -4, 2, -18, -6, -19, -8, -17,
    -- layer=1 filter=23 channel=40
    -11, 6, -6, -4, -13, -8, -25, -17, -6,
    -- layer=1 filter=23 channel=41
    4, -6, 43, 2, 6, -42, -7, -9, -6,
    -- layer=1 filter=23 channel=42
    0, 16, 17, -6, 13, 8, -20, 0, -5,
    -- layer=1 filter=23 channel=43
    -16, -18, -8, 8, -18, -7, -5, -1, 6,
    -- layer=1 filter=23 channel=44
    11, 20, 4, 15, 20, -3, 15, 1, 12,
    -- layer=1 filter=23 channel=45
    -7, 0, -6, 4, -5, -2, 12, -7, 0,
    -- layer=1 filter=23 channel=46
    -23, 7, -17, 0, 1, 1, 17, 16, 28,
    -- layer=1 filter=23 channel=47
    2, -15, 18, 0, 2, 0, 2, 22, 25,
    -- layer=1 filter=23 channel=48
    7, -5, 4, -3, 3, -6, 9, 2, 3,
    -- layer=1 filter=23 channel=49
    3, 0, 25, 4, 1, 18, 5, 5, 15,
    -- layer=1 filter=23 channel=50
    0, 1, 0, -8, -6, 15, -8, 0, 5,
    -- layer=1 filter=23 channel=51
    -13, 1, 0, -10, 2, -6, 4, 7, -6,
    -- layer=1 filter=23 channel=52
    12, 6, 6, 3, 1, 5, 15, 4, -4,
    -- layer=1 filter=23 channel=53
    6, 0, -2, 8, 5, 13, -2, 8, 3,
    -- layer=1 filter=23 channel=54
    -9, -6, -17, 6, -34, -2, 11, -5, -14,
    -- layer=1 filter=23 channel=55
    -6, -26, -2, -36, -36, -35, -26, -42, -36,
    -- layer=1 filter=23 channel=56
    3, 4, -1, 2, -1, -9, -8, 0, 5,
    -- layer=1 filter=23 channel=57
    -19, -8, -7, -10, 2, -27, -10, -4, -32,
    -- layer=1 filter=23 channel=58
    -19, -21, -6, 3, -16, 7, 1, 48, -9,
    -- layer=1 filter=23 channel=59
    15, -7, 9, 5, -2, 1, 5, -2, 15,
    -- layer=1 filter=23 channel=60
    -9, -2, -6, -13, -1, -14, -6, -7, -5,
    -- layer=1 filter=23 channel=61
    0, -1, -6, -1, -8, -13, -8, 4, -4,
    -- layer=1 filter=23 channel=62
    -4, -14, -21, 8, -26, 4, 14, 5, 1,
    -- layer=1 filter=23 channel=63
    -19, -5, -10, 4, -9, -8, -7, -16, 5,
    -- layer=1 filter=23 channel=64
    3, 10, 4, -13, 12, 0, 0, 7, 6,
    -- layer=1 filter=23 channel=65
    2, 2, -2, -5, 7, -4, 11, 2, -6,
    -- layer=1 filter=23 channel=66
    -1, -7, 6, -10, -2, 0, 3, -12, 0,
    -- layer=1 filter=23 channel=67
    -15, -22, -14, -45, -44, -27, -65, -70, -60,
    -- layer=1 filter=23 channel=68
    16, 14, 1, -6, 12, -2, 32, 7, 15,
    -- layer=1 filter=23 channel=69
    -7, 14, -24, 5, -13, 22, 0, -17, 10,
    -- layer=1 filter=23 channel=70
    -30, -42, 0, -25, -50, -42, -68, -59, -28,
    -- layer=1 filter=23 channel=71
    -6, 10, -1, 6, -3, -9, 1, -15, -10,
    -- layer=1 filter=23 channel=72
    -16, -17, -6, 0, -22, 1, 1, 4, 13,
    -- layer=1 filter=23 channel=73
    -4, 9, -1, -3, 5, 0, 9, -5, -1,
    -- layer=1 filter=23 channel=74
    2, 14, -3, -4, 14, 0, 5, -13, 15,
    -- layer=1 filter=23 channel=75
    -25, 1, -22, 1, -37, -13, -20, -6, -4,
    -- layer=1 filter=23 channel=76
    16, -4, 5, 12, 26, -10, 5, 2, 2,
    -- layer=1 filter=23 channel=77
    -8, 12, 6, 1, -1, -2, -5, -1, 8,
    -- layer=1 filter=23 channel=78
    -1, 2, -1, 7, 5, -3, -4, -2, 0,
    -- layer=1 filter=23 channel=79
    0, -15, -19, 15, -3, 0, 5, 7, 0,
    -- layer=1 filter=23 channel=80
    -8, 1, -5, 5, 5, -5, 4, 4, -6,
    -- layer=1 filter=23 channel=81
    0, 9, 11, -4, 3, -1, -6, -7, 4,
    -- layer=1 filter=23 channel=82
    4, 9, -9, 8, 15, 2, -7, 2, 1,
    -- layer=1 filter=23 channel=83
    9, 8, -14, 1, -13, 4, 9, -19, 3,
    -- layer=1 filter=23 channel=84
    -11, -11, 13, 18, 2, -25, -18, -13, 17,
    -- layer=1 filter=23 channel=85
    -18, -34, -17, -8, -6, -3, 16, 26, -5,
    -- layer=1 filter=23 channel=86
    -10, -9, -8, -18, -22, 3, -14, -9, -12,
    -- layer=1 filter=23 channel=87
    -7, -10, -12, -9, -12, 7, -11, -7, -5,
    -- layer=1 filter=23 channel=88
    8, 9, 10, 8, -2, -1, -3, -7, -12,
    -- layer=1 filter=23 channel=89
    -6, 11, 8, 5, 0, 0, 8, 10, 10,
    -- layer=1 filter=23 channel=90
    -1, 16, -5, 2, 2, 1, 17, -3, 9,
    -- layer=1 filter=23 channel=91
    0, -6, -3, 8, 5, 9, 8, 10, 8,
    -- layer=1 filter=23 channel=92
    14, -26, -10, 6, -9, -28, -1, 2, -18,
    -- layer=1 filter=23 channel=93
    0, 14, -9, 14, 17, -5, 0, 2, -1,
    -- layer=1 filter=23 channel=94
    10, 3, -1, 2, 7, 0, 14, -9, -7,
    -- layer=1 filter=23 channel=95
    -16, 2, 0, 13, -3, -4, -3, -6, 18,
    -- layer=1 filter=23 channel=96
    -16, -6, 1, -3, -3, 0, 3, -8, 2,
    -- layer=1 filter=23 channel=97
    7, 13, -3, 11, -2, -5, 3, 10, -4,
    -- layer=1 filter=23 channel=98
    -15, -20, -14, -11, -1, 1, 6, 7, -2,
    -- layer=1 filter=23 channel=99
    0, 9, 6, -12, 11, 8, 22, 9, 22,
    -- layer=1 filter=23 channel=100
    -14, -5, -12, -10, -15, -34, 2, -18, 12,
    -- layer=1 filter=23 channel=101
    1, 10, -3, 10, 9, 5, 1, 0, 0,
    -- layer=1 filter=23 channel=102
    3, -1, 13, 23, 10, 5, 19, 12, 4,
    -- layer=1 filter=23 channel=103
    -5, -7, -4, -8, -13, -4, -11, -4, 0,
    -- layer=1 filter=23 channel=104
    6, -26, -4, 3, -24, 0, 18, 8, -6,
    -- layer=1 filter=23 channel=105
    -3, 5, 0, 12, 0, 8, -5, -7, -7,
    -- layer=1 filter=23 channel=106
    7, -4, -5, 7, 8, -6, 8, 11, 7,
    -- layer=1 filter=23 channel=107
    7, 0, -2, -17, 0, -15, -12, 5, 0,
    -- layer=1 filter=23 channel=108
    18, 9, 6, 1, -1, 7, 12, 0, 2,
    -- layer=1 filter=23 channel=109
    -8, -7, 4, 6, -11, 0, -2, 1, -4,
    -- layer=1 filter=23 channel=110
    3, 8, 5, 9, -7, -3, 9, 0, -7,
    -- layer=1 filter=23 channel=111
    -14, 6, 7, 40, 0, 0, 8, -9, 24,
    -- layer=1 filter=23 channel=112
    -7, 2, -2, -4, -1, 9, -12, -14, -16,
    -- layer=1 filter=23 channel=113
    -20, -5, -3, 13, 14, 14, -8, 8, -8,
    -- layer=1 filter=23 channel=114
    -17, -15, -22, -25, -57, -29, -47, -57, -29,
    -- layer=1 filter=23 channel=115
    -18, -7, -11, -2, -17, 0, -2, -6, -26,
    -- layer=1 filter=23 channel=116
    8, 0, 2, -8, -8, 1, -1, -2, 0,
    -- layer=1 filter=23 channel=117
    -8, -9, -8, -9, -10, -2, -18, -14, -17,
    -- layer=1 filter=23 channel=118
    -10, -4, 0, 29, 3, -13, -6, -3, 8,
    -- layer=1 filter=23 channel=119
    0, 11, 14, 12, 3, -1, 14, 1, -5,
    -- layer=1 filter=23 channel=120
    -8, 0, 6, 4, 4, 7, 7, -3, -1,
    -- layer=1 filter=23 channel=121
    -25, -13, -28, -24, -24, -17, 1, -23, 1,
    -- layer=1 filter=23 channel=122
    4, -7, 8, -4, -2, 5, 7, 0, -7,
    -- layer=1 filter=23 channel=123
    -7, -25, -19, -17, -20, -22, -7, -3, -14,
    -- layer=1 filter=23 channel=124
    -11, -3, -5, 0, -5, -11, -4, 7, 4,
    -- layer=1 filter=23 channel=125
    -18, -18, 6, -20, -14, -32, -23, -32, -27,
    -- layer=1 filter=23 channel=126
    1, -13, -6, -7, -9, 14, 28, -8, 3,
    -- layer=1 filter=23 channel=127
    -22, -14, -9, 17, -6, -15, -11, -9, 17,
    -- layer=1 filter=24 channel=0
    19, 17, 12, 13, -13, -10, -9, -15, -14,
    -- layer=1 filter=24 channel=1
    27, -10, -10, -53, -34, 23, -13, 30, 19,
    -- layer=1 filter=24 channel=2
    -68, -62, 7, 9, 4, 18, 20, 27, 9,
    -- layer=1 filter=24 channel=3
    3, -2, 0, -5, -13, 4, 0, -11, -7,
    -- layer=1 filter=24 channel=4
    -2, 3, -6, 0, 0, -1, 3, 2, 0,
    -- layer=1 filter=24 channel=5
    19, -22, -26, -66, -35, 21, -19, 21, -19,
    -- layer=1 filter=24 channel=6
    -4, 31, 30, 4, 19, -6, 21, -8, -25,
    -- layer=1 filter=24 channel=7
    33, -42, -10, -14, -2, 19, 18, 12, 13,
    -- layer=1 filter=24 channel=8
    23, -18, -21, -65, -34, 28, 9, 40, 8,
    -- layer=1 filter=24 channel=9
    -22, -30, 14, 19, 43, 48, -14, 19, -28,
    -- layer=1 filter=24 channel=10
    14, -50, -2, -11, -10, 26, 24, 2, 1,
    -- layer=1 filter=24 channel=11
    9, 7, 26, 0, 8, -2, 0, -13, -30,
    -- layer=1 filter=24 channel=12
    -77, -45, -16, 9, 7, -2, 20, -4, 20,
    -- layer=1 filter=24 channel=13
    -8, 13, 8, 11, 16, -11, 20, 1, -21,
    -- layer=1 filter=24 channel=14
    0, -47, -26, 8, -15, 13, -4, -3, 11,
    -- layer=1 filter=24 channel=15
    -19, 2, -25, -76, -38, 8, 17, 36, 11,
    -- layer=1 filter=24 channel=16
    0, -30, -29, -57, 1, 23, 4, 30, 0,
    -- layer=1 filter=24 channel=17
    15, 20, -3, -2, -3, -17, -1, 8, -25,
    -- layer=1 filter=24 channel=18
    -36, -5, 26, 11, 26, 9, -3, -36, -35,
    -- layer=1 filter=24 channel=19
    33, 3, 13, 29, 77, 76, 59, 38, -40,
    -- layer=1 filter=24 channel=20
    -5, 1, 0, -19, -1, -10, 11, -6, -6,
    -- layer=1 filter=24 channel=21
    6, 0, -10, -8, -28, 1, 0, 21, 14,
    -- layer=1 filter=24 channel=22
    15, 26, -12, -6, -34, -26, -4, 20, 11,
    -- layer=1 filter=24 channel=23
    35, 14, 3, -31, 6, 54, 12, 47, -3,
    -- layer=1 filter=24 channel=24
    -21, -33, -23, -24, -3, -1, 8, -15, -13,
    -- layer=1 filter=24 channel=25
    33, -32, -12, -9, 36, 37, 18, 27, 19,
    -- layer=1 filter=24 channel=26
    -27, -14, 17, 15, 28, 7, 19, 17, 1,
    -- layer=1 filter=24 channel=27
    71, 47, 47, 32, 24, 2, 0, -33, -43,
    -- layer=1 filter=24 channel=28
    25, -27, -29, 4, -36, 14, -10, 24, 6,
    -- layer=1 filter=24 channel=29
    54, 2, 17, 10, -22, -30, -16, -46, -41,
    -- layer=1 filter=24 channel=30
    -46, -45, 41, -13, 45, 16, 14, -7, -51,
    -- layer=1 filter=24 channel=31
    -32, -10, 30, 16, 31, 17, -4, -30, -50,
    -- layer=1 filter=24 channel=32
    -30, -24, 9, 16, 23, 27, 11, 9, -8,
    -- layer=1 filter=24 channel=33
    17, 17, 8, 7, -12, -2, -7, -15, -11,
    -- layer=1 filter=24 channel=34
    0, 3, -5, 7, 12, 0, 11, 13, -14,
    -- layer=1 filter=24 channel=35
    -5, -1, -1, 10, 0, -4, 1, -2, 3,
    -- layer=1 filter=24 channel=36
    6, -1, 15, 7, -6, -7, -25, -30, -30,
    -- layer=1 filter=24 channel=37
    16, -21, -18, -41, 4, 33, 4, 0, -16,
    -- layer=1 filter=24 channel=38
    -3, 12, 19, -2, -1, -3, -1, -14, -7,
    -- layer=1 filter=24 channel=39
    10, 0, -1, -8, -11, -8, -14, -8, -25,
    -- layer=1 filter=24 channel=40
    -22, 13, 17, 7, 0, 3, -8, -26, -32,
    -- layer=1 filter=24 channel=41
    -34, -36, 8, 16, 46, 61, 19, 25, -38,
    -- layer=1 filter=24 channel=42
    -34, -66, -27, -4, -2, 6, 32, 22, 28,
    -- layer=1 filter=24 channel=43
    12, -15, -23, -55, -25, 22, 2, 46, 19,
    -- layer=1 filter=24 channel=44
    -22, 6, 13, 10, 13, 1, 12, -12, -4,
    -- layer=1 filter=24 channel=45
    -9, 7, -21, -9, -3, -15, 0, 12, 13,
    -- layer=1 filter=24 channel=46
    22, -7, -5, 14, 23, 6, 36, -10, -60,
    -- layer=1 filter=24 channel=47
    -7, -20, 17, 31, 39, 58, 45, 28, -33,
    -- layer=1 filter=24 channel=48
    12, -3, 8, -13, -11, 0, 14, -20, -16,
    -- layer=1 filter=24 channel=49
    -13, -3, 9, 15, 4, -4, 3, -11, -9,
    -- layer=1 filter=24 channel=50
    -14, -19, -11, -7, -10, -9, -23, -20, -18,
    -- layer=1 filter=24 channel=51
    23, -5, 20, -3, -15, 8, 4, 11, 16,
    -- layer=1 filter=24 channel=52
    -3, 4, -13, 6, 9, 4, 13, 31, 19,
    -- layer=1 filter=24 channel=53
    0, -3, 3, 4, 0, 4, -8, 1, 4,
    -- layer=1 filter=24 channel=54
    53, -52, 2, -15, 63, 53, 36, 32, 12,
    -- layer=1 filter=24 channel=55
    15, -5, 11, -4, -19, -6, -1, -10, -8,
    -- layer=1 filter=24 channel=56
    -5, 6, -7, 4, 0, 12, 2, -3, -1,
    -- layer=1 filter=24 channel=57
    15, -29, 11, -15, -3, 10, 8, 1, -2,
    -- layer=1 filter=24 channel=58
    26, -6, 37, -4, 42, 63, 37, 41, -3,
    -- layer=1 filter=24 channel=59
    0, -5, -5, 0, 5, 1, 4, 20, -6,
    -- layer=1 filter=24 channel=60
    5, 6, 15, 0, 10, 13, 1, 7, 0,
    -- layer=1 filter=24 channel=61
    8, -2, 8, 16, -2, 1, 8, 8, -12,
    -- layer=1 filter=24 channel=62
    9, -40, -16, -56, 8, 33, 16, 35, 15,
    -- layer=1 filter=24 channel=63
    9, -2, 12, 22, 9, -20, -5, -41, -20,
    -- layer=1 filter=24 channel=64
    7, -2, -1, 4, -2, -1, -8, 12, 1,
    -- layer=1 filter=24 channel=65
    -12, 2, -12, 10, -28, -11, 3, -2, 4,
    -- layer=1 filter=24 channel=66
    27, 1, -2, 11, -22, -7, -25, -27, -5,
    -- layer=1 filter=24 channel=67
    7, 22, 20, 1, -10, -10, 9, -10, -20,
    -- layer=1 filter=24 channel=68
    -22, 13, 25, 28, 24, 6, 10, -8, 17,
    -- layer=1 filter=24 channel=69
    -29, -38, -37, -50, -43, 12, 19, 20, -5,
    -- layer=1 filter=24 channel=70
    13, 12, 21, -1, -3, 0, 0, -10, -49,
    -- layer=1 filter=24 channel=71
    1, -23, -21, -15, -24, -1, -17, -12, 0,
    -- layer=1 filter=24 channel=72
    -15, -17, 9, 31, 55, 65, 34, 10, -31,
    -- layer=1 filter=24 channel=73
    -3, -6, -6, 3, 6, 9, -15, 2, -5,
    -- layer=1 filter=24 channel=74
    -10, -19, 29, 22, 49, 2, -7, -18, 2,
    -- layer=1 filter=24 channel=75
    -88, -44, 2, -12, 10, -20, -5, -65, -29,
    -- layer=1 filter=24 channel=76
    -11, -17, 29, 24, 31, -18, -3, -22, -25,
    -- layer=1 filter=24 channel=77
    -13, -25, -14, -10, -19, -5, -3, 0, 11,
    -- layer=1 filter=24 channel=78
    0, 1, -7, 9, -2, -2, -12, 6, -17,
    -- layer=1 filter=24 channel=79
    1, -29, -23, -55, 0, 23, 22, 25, 9,
    -- layer=1 filter=24 channel=80
    3, 9, -3, 2, -3, -4, -1, -3, 3,
    -- layer=1 filter=24 channel=81
    22, -9, -17, -29, -41, -22, -10, -7, -3,
    -- layer=1 filter=24 channel=82
    -3, -2, 4, -3, -20, -3, -7, -11, 13,
    -- layer=1 filter=24 channel=83
    -10, 10, -7, -20, -23, 16, 8, 17, 20,
    -- layer=1 filter=24 channel=84
    -11, 14, 61, 57, 65, 11, 10, -21, -11,
    -- layer=1 filter=24 channel=85
    32, 1, 28, 11, 31, 53, 18, 40, -24,
    -- layer=1 filter=24 channel=86
    21, 17, 3, -6, -1, -8, -14, -18, -17,
    -- layer=1 filter=24 channel=87
    6, -5, -9, 29, 67, 75, 38, 26, -55,
    -- layer=1 filter=24 channel=88
    -14, 8, 8, 1, -5, -10, 4, -1, 1,
    -- layer=1 filter=24 channel=89
    -11, 15, -1, 26, -17, -31, 2, -28, 0,
    -- layer=1 filter=24 channel=90
    -22, -17, 11, 3, -11, -16, 13, 13, 5,
    -- layer=1 filter=24 channel=91
    -1, 12, 18, 4, 0, -1, 0, -8, -28,
    -- layer=1 filter=24 channel=92
    -32, 9, 20, -13, 8, 38, -3, 16, 21,
    -- layer=1 filter=24 channel=93
    10, -2, -4, -15, -39, -12, -14, -14, 13,
    -- layer=1 filter=24 channel=94
    -1, 15, 13, 1, -14, -3, -15, -16, -12,
    -- layer=1 filter=24 channel=95
    -31, -5, 45, 38, 58, -3, 6, -26, -24,
    -- layer=1 filter=24 channel=96
    9, 18, 14, 2, 5, -8, -10, -4, -15,
    -- layer=1 filter=24 channel=97
    9, 2, -3, -12, -27, -10, -27, -11, -3,
    -- layer=1 filter=24 channel=98
    6, -20, -24, -70, -40, -3, 15, 42, 35,
    -- layer=1 filter=24 channel=99
    15, -18, -32, 2, -40, -20, -26, 23, 0,
    -- layer=1 filter=24 channel=100
    15, 13, 25, 25, 14, -9, -15, -32, -34,
    -- layer=1 filter=24 channel=101
    -2, 22, 14, -8, -1, -26, -6, -14, -1,
    -- layer=1 filter=24 channel=102
    -15, 17, 4, 12, 2, -18, -11, -12, -5,
    -- layer=1 filter=24 channel=103
    33, 24, 25, 29, 7, 7, -4, -2, -32,
    -- layer=1 filter=24 channel=104
    9, -11, 2, 3, 23, 30, 16, 32, 1,
    -- layer=1 filter=24 channel=105
    18, 16, -9, -8, -14, -18, -29, -27, -7,
    -- layer=1 filter=24 channel=106
    -7, 8, 27, 7, 27, -23, 21, -22, -10,
    -- layer=1 filter=24 channel=107
    -3, -7, -24, -11, -21, -19, -19, -8, -6,
    -- layer=1 filter=24 channel=108
    -23, -23, -9, 4, 4, -2, 22, 12, -12,
    -- layer=1 filter=24 channel=109
    6, -10, 2, -5, -4, -6, 7, 3, 5,
    -- layer=1 filter=24 channel=110
    14, -3, 2, -2, -5, -3, -10, -8, -12,
    -- layer=1 filter=24 channel=111
    -57, -29, 32, 6, 34, 6, 6, -45, -61,
    -- layer=1 filter=24 channel=112
    -16, 1, 27, 49, 37, -17, 16, -41, 13,
    -- layer=1 filter=24 channel=113
    19, -1, -8, -23, -27, -17, 9, -19, -26,
    -- layer=1 filter=24 channel=114
    21, -7, -36, -47, -34, -10, -10, 11, -24,
    -- layer=1 filter=24 channel=115
    12, 10, -2, -17, -14, 1, -20, -20, 7,
    -- layer=1 filter=24 channel=116
    4, 7, -2, -8, -12, -2, -10, 8, -2,
    -- layer=1 filter=24 channel=117
    -36, -16, 22, 35, 19, 0, 3, -20, -20,
    -- layer=1 filter=24 channel=118
    -33, -27, 40, 8, 37, 3, -9, -20, -31,
    -- layer=1 filter=24 channel=119
    -24, -11, 21, 22, 31, 28, 25, 13, -7,
    -- layer=1 filter=24 channel=120
    16, -29, 2, -21, -2, 15, 4, 16, 10,
    -- layer=1 filter=24 channel=121
    -16, -20, 9, 0, 11, 10, -1, -20, -64,
    -- layer=1 filter=24 channel=122
    -4, -10, -8, -3, 5, 1, 0, -4, 3,
    -- layer=1 filter=24 channel=123
    -2, 10, 8, 0, 17, 7, -3, -18, -37,
    -- layer=1 filter=24 channel=124
    5, -3, 2, -5, -16, -7, 9, -7, -6,
    -- layer=1 filter=24 channel=125
    12, 15, 14, 0, 3, -1, 8, -17, -38,
    -- layer=1 filter=24 channel=126
    -10, -13, -49, -39, -68, 0, 13, 38, 19,
    -- layer=1 filter=24 channel=127
    -51, -22, 42, 24, 55, 18, 21, -18, -20,
    -- layer=1 filter=25 channel=0
    -8, -13, -21, -15, -24, -15, 0, -4, -3,
    -- layer=1 filter=25 channel=1
    -8, -4, 23, 1, -5, 17, -14, 11, -27,
    -- layer=1 filter=25 channel=2
    35, 29, 11, 10, -30, -22, -11, -35, -45,
    -- layer=1 filter=25 channel=3
    7, -4, -1, 3, -2, -4, -1, -2, 3,
    -- layer=1 filter=25 channel=4
    -7, 13, -5, -12, -10, -12, 4, 2, 0,
    -- layer=1 filter=25 channel=5
    -4, -4, 0, 13, 37, 27, 30, 27, 12,
    -- layer=1 filter=25 channel=6
    19, 17, 13, 12, 30, 0, -4, -11, -27,
    -- layer=1 filter=25 channel=7
    -40, -7, 11, -9, 10, -12, 10, 13, -10,
    -- layer=1 filter=25 channel=8
    9, 20, 9, 9, -8, 0, -17, -12, -42,
    -- layer=1 filter=25 channel=9
    10, 33, 2, -14, -29, -18, -6, -37, 14,
    -- layer=1 filter=25 channel=10
    -26, -15, -5, -14, 21, -20, 18, -6, -16,
    -- layer=1 filter=25 channel=11
    -16, -24, -6, 0, -16, -16, 26, 16, 25,
    -- layer=1 filter=25 channel=12
    16, 41, 20, -17, 17, -29, -42, -40, -62,
    -- layer=1 filter=25 channel=13
    31, 52, 35, 19, 21, 10, -9, -19, -32,
    -- layer=1 filter=25 channel=14
    -19, -25, -7, -30, -19, -26, -9, -13, -18,
    -- layer=1 filter=25 channel=15
    37, 21, 58, 16, 23, -9, 4, -1, -28,
    -- layer=1 filter=25 channel=16
    11, 15, 10, -11, 3, -3, 15, -4, 6,
    -- layer=1 filter=25 channel=17
    40, 68, 35, 39, 38, 14, 3, -1, -15,
    -- layer=1 filter=25 channel=18
    -17, -3, 7, 3, 35, -2, 2, -21, 15,
    -- layer=1 filter=25 channel=19
    40, 23, 26, -32, 11, -8, -3, -9, -11,
    -- layer=1 filter=25 channel=20
    25, 59, 23, 37, 40, 17, -7, -7, -25,
    -- layer=1 filter=25 channel=21
    -49, -60, -24, -31, -36, -26, -5, -6, -31,
    -- layer=1 filter=25 channel=22
    45, 66, 58, 38, 55, 38, -18, -13, -29,
    -- layer=1 filter=25 channel=23
    -34, -28, 3, -54, -53, -53, -7, 8, 1,
    -- layer=1 filter=25 channel=24
    -56, -71, -47, -52, -66, -29, 11, -15, 18,
    -- layer=1 filter=25 channel=25
    -29, 24, 5, -18, 7, 3, -5, 13, -17,
    -- layer=1 filter=25 channel=26
    37, 59, 48, 26, 18, 12, -3, 3, -19,
    -- layer=1 filter=25 channel=27
    25, 24, 35, 48, 41, 40, 65, 65, 65,
    -- layer=1 filter=25 channel=28
    -35, -2, 15, -40, 0, -14, -37, -10, -30,
    -- layer=1 filter=25 channel=29
    -40, -12, 10, -13, -8, 14, -4, 3, 22,
    -- layer=1 filter=25 channel=30
    -10, -54, -3, -23, 10, -20, -26, -35, -14,
    -- layer=1 filter=25 channel=31
    36, 48, 47, 40, 76, 46, 1, 4, -6,
    -- layer=1 filter=25 channel=32
    -48, -27, -8, 1, 4, -22, 13, 4, 13,
    -- layer=1 filter=25 channel=33
    36, 11, 6, 16, 11, -5, 2, -7, -14,
    -- layer=1 filter=25 channel=34
    -19, 1, -23, 21, 14, -20, -21, -11, -27,
    -- layer=1 filter=25 channel=35
    -6, -9, -4, -16, -18, -15, 1, -4, -6,
    -- layer=1 filter=25 channel=36
    0, -21, -16, -2, -32, -28, 24, 5, 22,
    -- layer=1 filter=25 channel=37
    0, 16, 24, 33, 61, 68, 37, 47, 56,
    -- layer=1 filter=25 channel=38
    25, 14, 22, 18, 31, 19, 0, -20, -13,
    -- layer=1 filter=25 channel=39
    -8, -15, -16, -19, -32, -14, 5, -7, 17,
    -- layer=1 filter=25 channel=40
    42, 54, 43, 50, 47, 29, -3, -20, -24,
    -- layer=1 filter=25 channel=41
    -56, -18, -24, -10, -13, -5, 21, 23, 25,
    -- layer=1 filter=25 channel=42
    61, 53, 41, -16, -2, -26, -41, -32, -53,
    -- layer=1 filter=25 channel=43
    -15, -13, -10, -10, -7, -2, -18, -12, -31,
    -- layer=1 filter=25 channel=44
    7, 9, 17, 15, 8, 6, 19, 4, -9,
    -- layer=1 filter=25 channel=45
    -22, -20, -24, 4, -5, -13, 8, -8, -20,
    -- layer=1 filter=25 channel=46
    62, 37, 9, 6, -7, -10, -28, -38, -47,
    -- layer=1 filter=25 channel=47
    -24, 1, 12, 11, 26, 18, 16, 9, 25,
    -- layer=1 filter=25 channel=48
    -22, -21, -21, -39, -34, -44, -10, -30, -39,
    -- layer=1 filter=25 channel=49
    0, -2, -11, 18, 11, -20, -5, -30, -28,
    -- layer=1 filter=25 channel=50
    22, 24, 30, 8, 12, 12, -2, 9, 5,
    -- layer=1 filter=25 channel=51
    -27, -7, -3, -20, -6, -8, -5, -11, -29,
    -- layer=1 filter=25 channel=52
    -15, -10, 14, 19, 15, 15, -7, 26, 22,
    -- layer=1 filter=25 channel=53
    -5, -1, -9, -17, -2, -8, -5, -2, -7,
    -- layer=1 filter=25 channel=54
    -33, -1, -10, -15, 36, 5, 7, 23, 17,
    -- layer=1 filter=25 channel=55
    -33, -30, -13, 6, -23, -19, 39, 31, 58,
    -- layer=1 filter=25 channel=56
    -9, -2, -8, -3, -9, -5, 1, 0, -2,
    -- layer=1 filter=25 channel=57
    40, 47, 42, 30, 67, 28, 30, 17, 4,
    -- layer=1 filter=25 channel=58
    -35, -13, 5, -32, 0, -31, 15, -36, 10,
    -- layer=1 filter=25 channel=59
    0, -16, -9, -8, -15, -9, -5, 5, -18,
    -- layer=1 filter=25 channel=60
    -12, -14, -22, -17, -31, -7, 0, 0, -8,
    -- layer=1 filter=25 channel=61
    4, 5, -6, 15, -5, 6, 10, 4, 12,
    -- layer=1 filter=25 channel=62
    -1, 9, 12, -4, 10, 0, -7, -11, -25,
    -- layer=1 filter=25 channel=63
    -31, -45, -21, -23, -3, -14, 45, 17, 35,
    -- layer=1 filter=25 channel=64
    -13, 5, -4, -7, -2, 0, -13, -12, -9,
    -- layer=1 filter=25 channel=65
    -33, -37, -21, -25, -41, -44, -28, -25, -31,
    -- layer=1 filter=25 channel=66
    -6, -38, -40, 5, -20, -18, 36, 30, 28,
    -- layer=1 filter=25 channel=67
    -35, -44, -55, -55, -76, -60, -18, -54, -73,
    -- layer=1 filter=25 channel=68
    -14, -19, -15, 15, 1, 0, 21, -22, -6,
    -- layer=1 filter=25 channel=69
    6, 3, 26, -29, -2, 1, 0, -14, -20,
    -- layer=1 filter=25 channel=70
    4, 7, -6, 14, 41, 4, -3, 4, -22,
    -- layer=1 filter=25 channel=71
    -38, -79, -33, -33, -71, -38, 18, 9, 8,
    -- layer=1 filter=25 channel=72
    29, 18, 24, 18, 0, 2, -3, -9, -26,
    -- layer=1 filter=25 channel=73
    -2, -11, -9, -2, 0, -12, -3, 8, 4,
    -- layer=1 filter=25 channel=74
    -13, 5, -13, 14, 19, 12, -10, -37, -19,
    -- layer=1 filter=25 channel=75
    -22, -18, -31, -35, -16, -47, -9, -32, -43,
    -- layer=1 filter=25 channel=76
    -45, -41, -9, -14, -17, -31, -5, -41, 8,
    -- layer=1 filter=25 channel=77
    -69, -65, -29, -37, -55, -32, 29, 15, 0,
    -- layer=1 filter=25 channel=78
    -12, 16, 3, 0, 16, 11, -1, 22, 4,
    -- layer=1 filter=25 channel=79
    10, 32, 41, 10, 5, -12, -2, -18, -3,
    -- layer=1 filter=25 channel=80
    -5, -8, -3, 4, 8, -2, 0, 0, 10,
    -- layer=1 filter=25 channel=81
    -32, -39, -26, -49, -58, -52, 17, -9, 44,
    -- layer=1 filter=25 channel=82
    -63, -60, -35, -47, -53, -33, -38, -34, -21,
    -- layer=1 filter=25 channel=83
    -29, -10, 6, -23, 3, -4, 1, -6, -24,
    -- layer=1 filter=25 channel=84
    16, 34, 40, 24, 40, 0, -3, -22, -5,
    -- layer=1 filter=25 channel=85
    -18, -11, 16, -2, 18, 1, -2, -17, 17,
    -- layer=1 filter=25 channel=86
    40, 19, 3, 37, 20, 15, 18, 16, 4,
    -- layer=1 filter=25 channel=87
    36, 32, 13, 5, 21, -17, 20, -9, -18,
    -- layer=1 filter=25 channel=88
    -18, -33, -37, -21, -14, -28, -12, -27, -46,
    -- layer=1 filter=25 channel=89
    -43, -66, -35, -34, -60, -58, -30, -44, -43,
    -- layer=1 filter=25 channel=90
    -21, -7, 25, -13, -8, 3, 10, -18, -22,
    -- layer=1 filter=25 channel=91
    3, 26, 28, 20, 34, 21, 7, 10, -1,
    -- layer=1 filter=25 channel=92
    -63, -56, -3, -42, -9, -57, 22, -33, -3,
    -- layer=1 filter=25 channel=93
    -66, -90, -64, -40, -69, -42, -11, -18, -13,
    -- layer=1 filter=25 channel=94
    17, 2, -1, 10, 13, -16, -9, 11, 0,
    -- layer=1 filter=25 channel=95
    -27, -24, -7, -1, 5, -26, -6, -32, -2,
    -- layer=1 filter=25 channel=96
    -15, -11, -15, 5, -9, -25, -2, 8, 7,
    -- layer=1 filter=25 channel=97
    -7, -17, -13, -38, -44, -21, 1, -5, -15,
    -- layer=1 filter=25 channel=98
    5, 41, 27, 2, 17, 0, -7, -18, -32,
    -- layer=1 filter=25 channel=99
    -30, -42, -34, -50, -29, -23, -30, -6, -42,
    -- layer=1 filter=25 channel=100
    -40, -46, 1, 3, 37, 10, 33, 27, 55,
    -- layer=1 filter=25 channel=101
    -2, 17, 11, 6, 17, 17, 1, -9, -12,
    -- layer=1 filter=25 channel=102
    -2, 3, 0, 0, 19, -4, -4, -20, -20,
    -- layer=1 filter=25 channel=103
    0, -20, -20, 21, 12, 11, 20, 43, 33,
    -- layer=1 filter=25 channel=104
    -31, 18, 3, 1, 3, -5, -11, -7, 0,
    -- layer=1 filter=25 channel=105
    -8, -31, -30, -31, -37, -27, 10, -9, 2,
    -- layer=1 filter=25 channel=106
    20, 32, 5, 27, 22, 14, 1, -13, -17,
    -- layer=1 filter=25 channel=107
    15, -4, -14, -6, -2, -4, 7, 12, -3,
    -- layer=1 filter=25 channel=108
    1, -16, 4, 2, -2, -33, 25, -13, -11,
    -- layer=1 filter=25 channel=109
    -6, -2, -2, -1, 0, -6, -10, -9, -7,
    -- layer=1 filter=25 channel=110
    -5, 8, 2, -1, 0, -7, -8, 0, -17,
    -- layer=1 filter=25 channel=111
    -17, -35, 5, -16, 6, -51, -32, -82, -23,
    -- layer=1 filter=25 channel=112
    -26, -5, -5, 3, -8, -24, 8, -4, -11,
    -- layer=1 filter=25 channel=113
    39, 39, 44, 29, 43, 8, -3, -11, -15,
    -- layer=1 filter=25 channel=114
    -17, -55, -26, -25, 3, -17, 4, 6, 0,
    -- layer=1 filter=25 channel=115
    47, 36, 17, 28, 28, 9, 2, 0, -2,
    -- layer=1 filter=25 channel=116
    -6, -7, -2, 4, -1, 4, -9, 0, -1,
    -- layer=1 filter=25 channel=117
    22, -4, 13, 0, 35, -18, -5, -33, -12,
    -- layer=1 filter=25 channel=118
    -17, -32, -5, -1, 11, -26, -9, -32, -15,
    -- layer=1 filter=25 channel=119
    -46, -38, -31, -10, -22, -37, 17, 0, -12,
    -- layer=1 filter=25 channel=120
    -38, -15, -19, -21, 2, 0, 9, -8, -14,
    -- layer=1 filter=25 channel=121
    16, 1, -21, -3, -3, -7, 0, 11, 10,
    -- layer=1 filter=25 channel=122
    -3, 1, -2, 5, 6, -1, 1, -2, -4,
    -- layer=1 filter=25 channel=123
    -9, -45, -51, 6, -6, -12, 40, 36, 29,
    -- layer=1 filter=25 channel=124
    0, -9, -8, 1, -16, 3, -14, -1, 3,
    -- layer=1 filter=25 channel=125
    -16, 2, -11, 7, 25, 2, -15, -23, -22,
    -- layer=1 filter=25 channel=126
    -31, 14, 41, -6, 12, 16, -6, -1, -28,
    -- layer=1 filter=25 channel=127
    -27, -43, 6, 1, 4, 3, -29, -29, -5,
    -- layer=1 filter=26 channel=0
    0, 15, 4, -14, 12, -13, -36, 18, 3,
    -- layer=1 filter=26 channel=1
    -23, -24, -6, -47, -33, -11, -16, 9, 9,
    -- layer=1 filter=26 channel=2
    -1, 30, 7, -17, 6, -22, 24, -4, 11,
    -- layer=1 filter=26 channel=3
    -2, 0, -8, 5, 6, 7, 4, 3, 9,
    -- layer=1 filter=26 channel=4
    -13, -13, -23, 6, 15, 0, 8, 14, -6,
    -- layer=1 filter=26 channel=5
    -30, -27, 9, -12, -21, -11, 13, 11, 18,
    -- layer=1 filter=26 channel=6
    6, 15, 13, -1, -18, -1, -6, -4, -28,
    -- layer=1 filter=26 channel=7
    -48, 43, -60, -54, 89, -99, -62, 53, -102,
    -- layer=1 filter=26 channel=8
    -39, -17, -18, -51, -16, -14, -1, -2, 13,
    -- layer=1 filter=26 channel=9
    -3, -40, -24, 14, -72, 57, 33, -26, 56,
    -- layer=1 filter=26 channel=10
    -87, 57, -68, -60, 95, -112, -66, 56, -109,
    -- layer=1 filter=26 channel=11
    27, 1, 29, 21, -32, 0, -2, -32, 2,
    -- layer=1 filter=26 channel=12
    -8, 17, 7, -8, -6, 18, 36, 30, 83,
    -- layer=1 filter=26 channel=13
    26, -28, 21, 26, -71, 25, 14, -74, 12,
    -- layer=1 filter=26 channel=14
    -32, -11, -26, -70, 56, -81, 7, 82, -95,
    -- layer=1 filter=26 channel=15
    12, -9, 17, 7, 31, 39, -20, -29, 34,
    -- layer=1 filter=26 channel=16
    -28, 0, -3, -24, 7, 2, 15, 16, 33,
    -- layer=1 filter=26 channel=17
    9, -8, -8, -29, -6, 0, -1, -36, 0,
    -- layer=1 filter=26 channel=18
    11, -1, 14, 12, -5, -30, -1, 19, 36,
    -- layer=1 filter=26 channel=19
    -70, -9, -23, -34, -5, -2, 19, -26, 46,
    -- layer=1 filter=26 channel=20
    13, 13, 22, 3, -29, -8, 14, -33, 9,
    -- layer=1 filter=26 channel=21
    -15, 15, 1, -42, 27, -25, -21, 29, -13,
    -- layer=1 filter=26 channel=22
    9, 1, -11, -11, -7, -4, -17, 0, -19,
    -- layer=1 filter=26 channel=23
    39, 57, 41, 43, 29, 89, 19, 46, 48,
    -- layer=1 filter=26 channel=24
    17, -50, 2, 32, -50, 35, 47, -43, 59,
    -- layer=1 filter=26 channel=25
    -66, 49, -80, -42, 78, -54, -31, 38, -27,
    -- layer=1 filter=26 channel=26
    40, -76, 26, 65, -125, 47, 46, -138, 56,
    -- layer=1 filter=26 channel=27
    30, -9, 4, 2, 0, -2, -12, -29, -27,
    -- layer=1 filter=26 channel=28
    -89, 41, -51, -79, 94, -101, -76, 78, -71,
    -- layer=1 filter=26 channel=29
    17, -4, -6, 28, 18, -19, 6, 1, -30,
    -- layer=1 filter=26 channel=30
    -3, 17, 2, -36, -28, -2, 9, 0, 23,
    -- layer=1 filter=26 channel=31
    10, 17, 12, 0, -30, -36, -14, 23, 8,
    -- layer=1 filter=26 channel=32
    19, -101, 11, 57, -110, 38, 35, -112, 46,
    -- layer=1 filter=26 channel=33
    29, -7, 2, -14, -22, -8, 35, -21, 0,
    -- layer=1 filter=26 channel=34
    30, 0, 1, -5, -7, 10, 9, 4, 16,
    -- layer=1 filter=26 channel=35
    -8, 3, -8, 2, 2, 0, -8, -18, -5,
    -- layer=1 filter=26 channel=36
    26, 0, 8, -2, -23, -3, -5, -40, 4,
    -- layer=1 filter=26 channel=37
    -55, 13, -11, -25, 15, -14, 11, 18, 54,
    -- layer=1 filter=26 channel=38
    5, 12, 30, 2, 9, -1, 12, -3, -1,
    -- layer=1 filter=26 channel=39
    -10, -25, -27, -16, -34, 14, -17, -10, -5,
    -- layer=1 filter=26 channel=40
    -11, 10, 17, -18, -26, -43, 15, 5, -21,
    -- layer=1 filter=26 channel=41
    -5, -57, -9, 36, -71, 54, 27, -74, 60,
    -- layer=1 filter=26 channel=42
    -20, 36, 6, -28, 28, -27, 0, 25, -18,
    -- layer=1 filter=26 channel=43
    -38, 20, -40, -48, 3, -19, -34, 21, 12,
    -- layer=1 filter=26 channel=44
    42, -101, 24, 51, -135, 59, 30, -148, 26,
    -- layer=1 filter=26 channel=45
    28, -35, 16, 39, -41, 32, 24, -17, 31,
    -- layer=1 filter=26 channel=46
    -21, 3, 27, -4, -2, -25, 41, 12, 38,
    -- layer=1 filter=26 channel=47
    44, 16, 15, 47, -18, 64, 35, -52, 24,
    -- layer=1 filter=26 channel=48
    -4, 6, 0, -24, 9, 12, -20, 0, -2,
    -- layer=1 filter=26 channel=49
    34, -3, 4, 25, -22, 49, 7, -52, 28,
    -- layer=1 filter=26 channel=50
    0, 4, -3, -3, 2, -6, -7, 5, 20,
    -- layer=1 filter=26 channel=51
    -43, 37, -12, -40, 53, -57, -44, 26, -31,
    -- layer=1 filter=26 channel=52
    1, 12, 35, 21, 31, 34, 20, 15, 26,
    -- layer=1 filter=26 channel=53
    15, 10, 1, 4, 17, 7, 14, 5, -2,
    -- layer=1 filter=26 channel=54
    -73, 56, -90, -11, 71, -62, -38, 36, 9,
    -- layer=1 filter=26 channel=55
    0, -15, -4, 26, -25, 14, 19, -23, 0,
    -- layer=1 filter=26 channel=56
    -2, -1, 4, -13, -6, -11, 9, 4, -7,
    -- layer=1 filter=26 channel=57
    -68, 38, -72, -62, 84, -100, -56, 44, -116,
    -- layer=1 filter=26 channel=58
    30, 71, 7, 42, 57, 64, 31, 30, 16,
    -- layer=1 filter=26 channel=59
    5, -23, -4, -7, -32, -15, -11, -11, -3,
    -- layer=1 filter=26 channel=60
    0, -30, 33, -18, -40, -1, 27, -49, 39,
    -- layer=1 filter=26 channel=61
    -1, -3, 2, 10, 5, 6, 8, 2, 5,
    -- layer=1 filter=26 channel=62
    -75, 1, -39, -53, -2, -25, -12, 15, 44,
    -- layer=1 filter=26 channel=63
    17, -19, 28, 21, -19, 10, -2, -20, 3,
    -- layer=1 filter=26 channel=64
    -14, 27, 13, -19, 3, -1, -25, 23, 3,
    -- layer=1 filter=26 channel=65
    -15, 4, 17, -30, 0, -19, -19, -4, -3,
    -- layer=1 filter=26 channel=66
    7, -5, -1, -12, 3, -8, -35, -10, -12,
    -- layer=1 filter=26 channel=67
    -13, -4, 37, -11, -19, 19, 12, -21, 29,
    -- layer=1 filter=26 channel=68
    50, -91, 43, 96, -126, 66, 61, -130, 33,
    -- layer=1 filter=26 channel=69
    4, -13, 11, 18, -33, 7, 24, -14, 33,
    -- layer=1 filter=26 channel=70
    -10, -16, 19, 0, 0, 29, 0, 11, 14,
    -- layer=1 filter=26 channel=71
    -27, 19, -2, -25, 31, -33, -23, 26, -2,
    -- layer=1 filter=26 channel=72
    -29, 6, 0, -10, -27, -10, 15, 2, 21,
    -- layer=1 filter=26 channel=73
    0, 12, 20, -12, -15, 5, 11, 0, 31,
    -- layer=1 filter=26 channel=74
    28, -35, 17, 53, 4, 38, 20, 6, 30,
    -- layer=1 filter=26 channel=75
    -13, 23, 10, -28, -6, -15, 20, 31, 30,
    -- layer=1 filter=26 channel=76
    30, -43, 20, 24, -53, 31, 8, -54, 18,
    -- layer=1 filter=26 channel=77
    0, -7, 9, -7, 7, 0, -3, 4, -10,
    -- layer=1 filter=26 channel=78
    -13, 21, -32, -10, 41, -42, -44, 23, -43,
    -- layer=1 filter=26 channel=79
    -30, -8, -35, -24, -12, 2, 16, 15, 54,
    -- layer=1 filter=26 channel=80
    -2, 17, 15, -28, -17, -11, -18, 8, 9,
    -- layer=1 filter=26 channel=81
    -12, -14, -22, -26, -24, 5, -14, 5, 16,
    -- layer=1 filter=26 channel=82
    -2, -7, -2, -11, 2, 2, -21, -16, -3,
    -- layer=1 filter=26 channel=83
    -7, -42, -5, 14, -21, 20, 5, -21, -19,
    -- layer=1 filter=26 channel=84
    14, -27, 23, 63, -44, 31, 9, -3, 64,
    -- layer=1 filter=26 channel=85
    14, 44, 0, 26, 60, 55, 39, 15, 84,
    -- layer=1 filter=26 channel=86
    11, 7, 1, -22, -9, -11, -14, 7, -22,
    -- layer=1 filter=26 channel=87
    -24, 4, -20, -4, -45, 25, 15, -22, 30,
    -- layer=1 filter=26 channel=88
    0, -16, 9, -17, -21, 17, -19, -23, 3,
    -- layer=1 filter=26 channel=89
    11, -29, 34, 14, -55, 21, -9, -37, 18,
    -- layer=1 filter=26 channel=90
    56, -118, 21, 70, -103, 56, 59, -98, 34,
    -- layer=1 filter=26 channel=91
    -12, 15, -8, -17, 20, -13, -29, -2, -24,
    -- layer=1 filter=26 channel=92
    47, -55, 25, 62, -65, 38, 46, -77, 52,
    -- layer=1 filter=26 channel=93
    -5, 0, 3, -9, -4, 3, -9, 0, 12,
    -- layer=1 filter=26 channel=94
    -3, 26, 19, -13, 14, -22, -43, 19, -10,
    -- layer=1 filter=26 channel=95
    9, -16, 14, 35, -37, 1, 8, -3, 24,
    -- layer=1 filter=26 channel=96
    6, -33, -6, -3, -27, -1, -1, -26, 6,
    -- layer=1 filter=26 channel=97
    5, 11, 1, -7, 0, -11, -22, -3, 8,
    -- layer=1 filter=26 channel=98
    -44, 7, -64, -70, 21, 0, -28, 32, 30,
    -- layer=1 filter=26 channel=99
    -7, 34, -5, 65, 121, -29, 49, 101, -43,
    -- layer=1 filter=26 channel=100
    9, -16, 19, 5, -37, 0, -5, -41, -4,
    -- layer=1 filter=26 channel=101
    12, 7, 19, 7, -13, 10, -19, -16, -18,
    -- layer=1 filter=26 channel=102
    7, 34, 29, -19, 20, -24, -17, -10, -8,
    -- layer=1 filter=26 channel=103
    20, 5, 25, 11, -14, -17, -10, 2, 19,
    -- layer=1 filter=26 channel=104
    -20, 12, -4, 15, 8, 14, 24, 0, 35,
    -- layer=1 filter=26 channel=105
    -6, 14, -6, -25, 22, -5, -34, 15, -11,
    -- layer=1 filter=26 channel=106
    48, -61, 20, 62, -83, 40, 25, -107, 25,
    -- layer=1 filter=26 channel=107
    -17, -4, -6, -19, -6, 0, -8, -12, 7,
    -- layer=1 filter=26 channel=108
    55, -76, 16, 68, -112, 56, 41, -96, 50,
    -- layer=1 filter=26 channel=109
    8, 3, -10, -1, -5, 7, 9, 4, 4,
    -- layer=1 filter=26 channel=110
    -28, -17, 1, -14, 0, -27, -16, 0, -25,
    -- layer=1 filter=26 channel=111
    -2, -15, 10, 2, -4, -4, -2, 19, 29,
    -- layer=1 filter=26 channel=112
    10, -24, -10, 27, 15, 16, -20, 18, 67,
    -- layer=1 filter=26 channel=113
    24, 65, 18, -22, 26, -29, -12, 1, -21,
    -- layer=1 filter=26 channel=114
    -16, -32, 22, -15, 8, 12, 6, 3, 12,
    -- layer=1 filter=26 channel=115
    -33, 37, -27, -53, 52, -43, -72, 30, -38,
    -- layer=1 filter=26 channel=116
    -7, -4, -4, 10, -9, 7, 4, 6, 1,
    -- layer=1 filter=26 channel=117
    -14, -40, -12, 9, 40, 11, 13, 51, 64,
    -- layer=1 filter=26 channel=118
    26, -3, 17, 39, -34, 10, 21, 1, 38,
    -- layer=1 filter=26 channel=119
    47, -97, 18, 60, -138, 64, 33, -151, 47,
    -- layer=1 filter=26 channel=120
    -20, 19, -34, -54, 31, -30, -20, 29, -11,
    -- layer=1 filter=26 channel=121
    -3, -3, 6, -2, 12, -20, 19, 22, 0,
    -- layer=1 filter=26 channel=122
    1, 9, 5, -1, 7, 5, 6, -7, -6,
    -- layer=1 filter=26 channel=123
    1, 7, 10, -6, 8, -20, 12, 17, -20,
    -- layer=1 filter=26 channel=124
    9, 0, 1, -2, 1, 2, -13, 2, -17,
    -- layer=1 filter=26 channel=125
    -19, 1, 22, 0, 43, 6, 21, 0, 6,
    -- layer=1 filter=26 channel=126
    -71, -4, -20, -54, -2, -24, -27, 2, -9,
    -- layer=1 filter=26 channel=127
    10, -11, 29, 20, -23, -1, 12, 15, 46,
    -- layer=1 filter=27 channel=0
    -10, 0, -9, 3, 0, -5, -10, 3, -2,
    -- layer=1 filter=27 channel=1
    -9, -8, 0, -5, 2, -8, 4, -10, 2,
    -- layer=1 filter=27 channel=2
    13, 8, -14, -8, -3, 12, 13, -4, 10,
    -- layer=1 filter=27 channel=3
    1, -3, -9, 3, -6, 3, -9, 4, -10,
    -- layer=1 filter=27 channel=4
    -8, -10, -6, -7, -1, -3, -2, -4, 6,
    -- layer=1 filter=27 channel=5
    -5, 12, 8, 3, -12, -8, -11, -15, 8,
    -- layer=1 filter=27 channel=6
    -12, -13, 0, 2, -2, -6, -9, -6, 0,
    -- layer=1 filter=27 channel=7
    -4, 4, -6, -17, -8, -4, -5, -6, -9,
    -- layer=1 filter=27 channel=8
    0, 5, -10, -9, -11, -4, -10, -16, 3,
    -- layer=1 filter=27 channel=9
    5, -8, -12, 10, 5, -5, 1, -4, 1,
    -- layer=1 filter=27 channel=10
    2, 6, -5, -9, 7, 7, 5, -8, 4,
    -- layer=1 filter=27 channel=11
    -7, -3, -12, 4, 0, -4, -2, -7, -17,
    -- layer=1 filter=27 channel=12
    8, -8, 5, -6, -7, 2, -15, 4, 7,
    -- layer=1 filter=27 channel=13
    -7, -4, -8, -15, -1, -17, 0, 0, -4,
    -- layer=1 filter=27 channel=14
    2, 2, -11, 3, -8, -8, -5, -1, 13,
    -- layer=1 filter=27 channel=15
    -13, -10, -10, -1, 0, -20, 8, -6, -10,
    -- layer=1 filter=27 channel=16
    11, 8, 7, 4, 8, 4, -17, 1, -3,
    -- layer=1 filter=27 channel=17
    -4, -10, 2, 1, 1, -6, -15, -10, -6,
    -- layer=1 filter=27 channel=18
    8, -4, -3, 8, 0, -9, 6, -9, -8,
    -- layer=1 filter=27 channel=19
    -4, -3, -10, -5, -2, 0, -6, -11, 4,
    -- layer=1 filter=27 channel=20
    -10, 0, -6, 0, 0, -8, 1, -16, 0,
    -- layer=1 filter=27 channel=21
    0, 2, -1, -12, -10, 4, -10, -4, -17,
    -- layer=1 filter=27 channel=22
    1, -12, -13, -7, -10, 2, 4, 6, 3,
    -- layer=1 filter=27 channel=23
    -14, 0, -7, 3, -6, -8, -5, -20, -7,
    -- layer=1 filter=27 channel=24
    -10, 4, -3, -8, 1, -3, -11, -5, -11,
    -- layer=1 filter=27 channel=25
    -14, -12, 11, 2, 0, 5, 9, -10, 1,
    -- layer=1 filter=27 channel=26
    -8, 11, -1, 3, -2, -1, 3, 5, 1,
    -- layer=1 filter=27 channel=27
    1, -12, -8, 6, -8, -1, -15, 2, 5,
    -- layer=1 filter=27 channel=28
    -4, -6, 4, -1, 6, 0, -3, -3, -18,
    -- layer=1 filter=27 channel=29
    0, -3, -3, -9, 4, -4, -15, -12, -9,
    -- layer=1 filter=27 channel=30
    -10, 6, 0, 3, 13, -7, -3, -14, -16,
    -- layer=1 filter=27 channel=31
    -8, -12, 0, 6, -12, -5, 6, -13, 4,
    -- layer=1 filter=27 channel=32
    -3, 0, -9, -7, -6, -8, 1, -5, -7,
    -- layer=1 filter=27 channel=33
    0, 1, 7, -4, 8, 10, 5, -1, 12,
    -- layer=1 filter=27 channel=34
    4, -4, 2, -9, -8, 2, -6, -8, 1,
    -- layer=1 filter=27 channel=35
    2, 5, 11, 4, -7, -4, -1, -9, -11,
    -- layer=1 filter=27 channel=36
    -11, 0, -14, -11, 0, -14, -13, 5, -5,
    -- layer=1 filter=27 channel=37
    4, 14, -1, 0, 3, -4, -7, -17, 9,
    -- layer=1 filter=27 channel=38
    -10, -2, -5, 0, 0, -9, 4, -4, -15,
    -- layer=1 filter=27 channel=39
    -5, -1, -1, 4, 4, -1, -2, -9, 2,
    -- layer=1 filter=27 channel=40
    -8, 3, -1, 6, -12, -17, 6, -7, 0,
    -- layer=1 filter=27 channel=41
    -10, -17, -9, -3, -11, 7, -11, -5, 3,
    -- layer=1 filter=27 channel=42
    -6, 6, -10, 0, -11, -4, 1, -1, 3,
    -- layer=1 filter=27 channel=43
    -2, 10, -1, 0, -4, 8, -12, 0, 9,
    -- layer=1 filter=27 channel=44
    -17, -7, -11, -2, -12, 2, -14, 1, 1,
    -- layer=1 filter=27 channel=45
    -13, 6, -18, 6, -12, -3, -10, 3, 7,
    -- layer=1 filter=27 channel=46
    -4, 3, -2, -7, -5, -4, -1, 3, -7,
    -- layer=1 filter=27 channel=47
    -2, -15, -9, 4, -2, -1, -3, -10, -11,
    -- layer=1 filter=27 channel=48
    -13, -10, -3, -9, 1, 0, -12, -6, 1,
    -- layer=1 filter=27 channel=49
    -4, -14, -11, -6, 2, 3, -7, -10, -6,
    -- layer=1 filter=27 channel=50
    2, -10, 9, -6, 1, -9, 5, -2, 4,
    -- layer=1 filter=27 channel=51
    -9, -12, 5, -16, -4, -12, -9, 5, -17,
    -- layer=1 filter=27 channel=52
    1, 0, -7, 7, -6, 8, -3, -2, -8,
    -- layer=1 filter=27 channel=53
    -10, -9, 5, 4, -2, -5, 8, -11, -4,
    -- layer=1 filter=27 channel=54
    -1, 7, 7, -3, 12, 4, 4, -9, -7,
    -- layer=1 filter=27 channel=55
    -1, -2, -3, 9, 0, -8, -14, -9, 1,
    -- layer=1 filter=27 channel=56
    -8, 7, -10, -10, -7, -2, 5, 0, -7,
    -- layer=1 filter=27 channel=57
    -3, 5, 8, -14, -6, 0, -8, -10, -15,
    -- layer=1 filter=27 channel=58
    0, -1, 8, 10, -3, 1, 5, -3, 2,
    -- layer=1 filter=27 channel=59
    6, -1, 9, 8, -8, -4, 4, 4, 1,
    -- layer=1 filter=27 channel=60
    3, -1, -5, -5, 0, -7, -1, 0, -4,
    -- layer=1 filter=27 channel=61
    1, 0, -7, 3, -6, 4, -6, -9, 5,
    -- layer=1 filter=27 channel=62
    6, -2, -8, 6, 4, -1, -17, -4, 0,
    -- layer=1 filter=27 channel=63
    -18, -16, 1, -7, -3, -1, -10, -7, 0,
    -- layer=1 filter=27 channel=64
    -1, -2, 2, -6, -13, -9, 8, 3, 1,
    -- layer=1 filter=27 channel=65
    -11, -8, 5, -2, -8, 2, -3, -13, -4,
    -- layer=1 filter=27 channel=66
    -6, 4, 1, -3, -6, -6, -6, 0, 0,
    -- layer=1 filter=27 channel=67
    0, 8, 5, 6, 4, 0, 4, -6, 12,
    -- layer=1 filter=27 channel=68
    -17, 13, 1, -3, 7, 2, -5, 7, -5,
    -- layer=1 filter=27 channel=69
    -12, -1, -4, -8, -4, -18, -10, -4, 6,
    -- layer=1 filter=27 channel=70
    -7, 1, -1, 6, -4, 10, -12, -3, 0,
    -- layer=1 filter=27 channel=71
    1, 4, 2, -9, -5, -10, 0, -13, -11,
    -- layer=1 filter=27 channel=72
    0, 5, 0, 7, -1, 4, -6, -14, 4,
    -- layer=1 filter=27 channel=73
    0, -10, 7, 4, 7, 5, 2, 0, -7,
    -- layer=1 filter=27 channel=74
    5, 3, -7, -6, 0, -10, -12, 3, 0,
    -- layer=1 filter=27 channel=75
    2, 8, 9, 7, 1, -7, 0, -16, -2,
    -- layer=1 filter=27 channel=76
    3, 2, -11, -3, 1, -9, 0, 0, -8,
    -- layer=1 filter=27 channel=77
    -8, 5, 3, 5, 3, 7, 0, 1, -1,
    -- layer=1 filter=27 channel=78
    -6, -7, 1, -11, 7, -16, -9, -4, 0,
    -- layer=1 filter=27 channel=79
    0, -8, 0, -8, 2, 5, -6, -6, -2,
    -- layer=1 filter=27 channel=80
    -7, -2, -1, 0, -11, -1, -2, -6, -1,
    -- layer=1 filter=27 channel=81
    1, -12, 4, -10, 1, 4, -2, -10, -11,
    -- layer=1 filter=27 channel=82
    0, -2, -16, -20, -19, -9, 4, -3, -1,
    -- layer=1 filter=27 channel=83
    -12, -10, -10, 8, -15, 4, 5, 2, 1,
    -- layer=1 filter=27 channel=84
    -12, 3, 13, -1, 0, -6, 5, 0, 0,
    -- layer=1 filter=27 channel=85
    -12, 0, -1, -8, -6, -6, 11, 0, -11,
    -- layer=1 filter=27 channel=86
    -12, 3, -4, -12, 6, -3, -15, -16, -14,
    -- layer=1 filter=27 channel=87
    5, -3, -6, -3, 5, -7, 3, -1, 0,
    -- layer=1 filter=27 channel=88
    -8, 0, -4, -2, -8, -9, -1, 8, -13,
    -- layer=1 filter=27 channel=89
    -12, -3, 1, 1, -1, -18, -16, -13, 1,
    -- layer=1 filter=27 channel=90
    -2, 4, -5, 5, -7, 7, -7, -6, -10,
    -- layer=1 filter=27 channel=91
    -15, -7, -6, 2, -8, -11, 2, -7, -9,
    -- layer=1 filter=27 channel=92
    0, -4, -4, -2, -6, -8, -10, -9, 0,
    -- layer=1 filter=27 channel=93
    -10, 3, -15, -4, -9, 1, -10, 2, -7,
    -- layer=1 filter=27 channel=94
    -9, -12, 0, -10, 1, -8, -7, 3, -14,
    -- layer=1 filter=27 channel=95
    -9, -2, -12, -5, 7, -10, -4, 0, -14,
    -- layer=1 filter=27 channel=96
    -10, 0, 4, 8, 2, 4, -6, 3, 8,
    -- layer=1 filter=27 channel=97
    2, -5, -8, 1, 0, -14, -3, 0, 2,
    -- layer=1 filter=27 channel=98
    -5, 1, 0, 1, 0, 7, -7, -16, -4,
    -- layer=1 filter=27 channel=99
    -15, 2, 3, -15, 9, -16, -8, 5, -16,
    -- layer=1 filter=27 channel=100
    -2, 1, 0, -1, 0, -14, -8, -14, -4,
    -- layer=1 filter=27 channel=101
    1, 1, -2, -3, -8, -6, -10, -9, -10,
    -- layer=1 filter=27 channel=102
    -5, -3, -12, -1, -2, -2, -4, -2, 0,
    -- layer=1 filter=27 channel=103
    1, 1, 2, -8, -11, -16, -7, -10, -12,
    -- layer=1 filter=27 channel=104
    -10, -7, 7, 1, 7, 2, -7, -1, 5,
    -- layer=1 filter=27 channel=105
    -3, -11, -18, 2, -12, 3, -17, -2, -17,
    -- layer=1 filter=27 channel=106
    0, 5, -11, -10, -12, 3, -12, -5, 1,
    -- layer=1 filter=27 channel=107
    -6, 6, -3, -11, -2, 4, 0, -1, 7,
    -- layer=1 filter=27 channel=108
    -7, -6, -10, 4, -16, 3, -6, -14, -3,
    -- layer=1 filter=27 channel=109
    4, 10, 9, -6, -2, 8, -2, 6, 10,
    -- layer=1 filter=27 channel=110
    2, -8, -4, 5, 0, -9, -9, 3, -5,
    -- layer=1 filter=27 channel=111
    7, -6, -3, -9, -8, -8, 7, -7, -15,
    -- layer=1 filter=27 channel=112
    -9, -6, 5, -11, -7, -6, 3, -2, -4,
    -- layer=1 filter=27 channel=113
    -11, -14, 1, -5, 0, 0, -13, 1, 6,
    -- layer=1 filter=27 channel=114
    7, 1, 9, -1, 3, -9, -3, -2, 3,
    -- layer=1 filter=27 channel=115
    -16, -10, 0, -6, -13, -11, -17, -6, -3,
    -- layer=1 filter=27 channel=116
    9, 7, -8, -3, -6, -10, 0, 0, 3,
    -- layer=1 filter=27 channel=117
    -8, 11, -9, 0, 4, -11, 5, 3, 0,
    -- layer=1 filter=27 channel=118
    4, 14, -9, -10, -5, -18, 9, 2, -17,
    -- layer=1 filter=27 channel=119
    1, -6, -3, -6, 3, 7, 4, 2, -7,
    -- layer=1 filter=27 channel=120
    0, 0, 0, -11, -11, -12, -1, -6, -2,
    -- layer=1 filter=27 channel=121
    -11, -14, -15, 3, 9, -6, -8, -6, -13,
    -- layer=1 filter=27 channel=122
    10, -3, 3, 1, -8, -4, 8, 4, -3,
    -- layer=1 filter=27 channel=123
    2, -17, 0, -13, 0, -5, 3, -2, -6,
    -- layer=1 filter=27 channel=124
    -11, 8, -9, -6, 5, 7, 0, -1, -1,
    -- layer=1 filter=27 channel=125
    -1, 1, -6, 8, 4, 14, -5, 8, 6,
    -- layer=1 filter=27 channel=126
    0, -5, 0, 6, -5, 12, -10, -6, 5,
    -- layer=1 filter=27 channel=127
    -4, 5, 12, 4, -9, -12, 8, -2, -2,
    -- layer=1 filter=28 channel=0
    4, 7, -6, -11, 0, -8, 7, -4, -1,
    -- layer=1 filter=28 channel=1
    4, -6, -8, -2, -9, -4, 5, 6, -6,
    -- layer=1 filter=28 channel=2
    -13, -11, -1, -10, -3, -2, -10, 0, 3,
    -- layer=1 filter=28 channel=3
    -3, 0, 4, 8, -4, 6, -10, 0, 2,
    -- layer=1 filter=28 channel=4
    3, -11, 3, 1, -11, -10, 3, -11, -9,
    -- layer=1 filter=28 channel=5
    0, -1, 3, -9, 5, -5, -8, 0, -8,
    -- layer=1 filter=28 channel=6
    1, -11, -10, -14, -10, -16, -19, -8, -17,
    -- layer=1 filter=28 channel=7
    -1, -14, -11, -2, -1, -21, -8, -11, -5,
    -- layer=1 filter=28 channel=8
    3, -1, -8, -5, 0, -1, 7, -10, -3,
    -- layer=1 filter=28 channel=9
    0, 2, -3, -8, -1, 8, -4, -4, 7,
    -- layer=1 filter=28 channel=10
    -12, -3, -9, -14, -2, -20, -14, -1, -16,
    -- layer=1 filter=28 channel=11
    -13, 0, -9, 0, -10, 6, -1, 7, -8,
    -- layer=1 filter=28 channel=12
    5, 7, 19, 0, -2, -4, 2, -9, 0,
    -- layer=1 filter=28 channel=13
    1, -1, -19, -16, 1, -1, -12, -11, -3,
    -- layer=1 filter=28 channel=14
    -12, 10, -3, -9, -10, -7, -16, 0, -6,
    -- layer=1 filter=28 channel=15
    2, 0, 0, -12, -4, -6, -2, -8, 0,
    -- layer=1 filter=28 channel=16
    -12, -8, -14, 4, -6, -12, 6, -9, -5,
    -- layer=1 filter=28 channel=17
    6, 3, -4, -3, 7, -13, 7, 3, 6,
    -- layer=1 filter=28 channel=18
    -14, 7, 5, 2, -9, -3, -10, 6, 5,
    -- layer=1 filter=28 channel=19
    -6, 7, -3, -5, 8, 0, 7, 8, -2,
    -- layer=1 filter=28 channel=20
    -12, -16, -14, -2, -8, -5, 0, -13, -8,
    -- layer=1 filter=28 channel=21
    -2, -14, -1, -5, 1, -10, -5, 0, -14,
    -- layer=1 filter=28 channel=22
    0, -9, -17, -12, -1, -10, -14, -7, -2,
    -- layer=1 filter=28 channel=23
    -5, 8, 4, -8, 7, -5, -5, -1, 6,
    -- layer=1 filter=28 channel=24
    -7, -7, 0, -10, 1, -5, -2, 0, 1,
    -- layer=1 filter=28 channel=25
    -11, -8, 2, -4, 0, -2, -14, -9, -4,
    -- layer=1 filter=28 channel=26
    -11, -7, -7, -10, -5, -12, -16, -19, -6,
    -- layer=1 filter=28 channel=27
    0, -9, 0, 12, -7, -9, -8, -5, 10,
    -- layer=1 filter=28 channel=28
    -9, -10, 3, -10, -2, 5, 2, 1, -8,
    -- layer=1 filter=28 channel=29
    0, -7, 12, -1, 2, -9, 9, -9, 5,
    -- layer=1 filter=28 channel=30
    -5, 0, -5, -1, -4, -15, -7, -10, -4,
    -- layer=1 filter=28 channel=31
    -6, 6, -4, 8, 0, -13, -18, -13, -11,
    -- layer=1 filter=28 channel=32
    -4, 5, -2, 4, -11, -7, 0, 4, 1,
    -- layer=1 filter=28 channel=33
    -1, 8, -3, -2, 9, 4, 1, 4, -1,
    -- layer=1 filter=28 channel=34
    -6, -5, -10, 0, -10, 2, -9, 3, -11,
    -- layer=1 filter=28 channel=35
    -10, -8, -3, 0, 6, 2, 0, 5, -7,
    -- layer=1 filter=28 channel=36
    -1, -9, 7, 5, 7, -6, -8, -12, -11,
    -- layer=1 filter=28 channel=37
    -15, -10, -11, -15, -8, 2, 0, -4, -13,
    -- layer=1 filter=28 channel=38
    -9, -13, -9, -13, -18, -20, 1, -18, -10,
    -- layer=1 filter=28 channel=39
    -7, 4, 3, -11, 8, -4, -2, 0, -10,
    -- layer=1 filter=28 channel=40
    8, -13, -13, -7, 1, -6, -5, -17, -15,
    -- layer=1 filter=28 channel=41
    5, -10, 0, -4, 7, 4, 2, -10, -7,
    -- layer=1 filter=28 channel=42
    -15, -3, -11, -9, -2, -12, -9, -19, -2,
    -- layer=1 filter=28 channel=43
    -5, -9, -9, 2, -8, -10, 0, -3, 8,
    -- layer=1 filter=28 channel=44
    0, 4, -6, 7, -7, 1, 3, 3, 0,
    -- layer=1 filter=28 channel=45
    2, 3, 4, -7, 5, 3, 3, 6, 1,
    -- layer=1 filter=28 channel=46
    -20, -2, 2, -9, -7, -1, -8, -1, 1,
    -- layer=1 filter=28 channel=47
    3, -15, -7, -8, 1, 3, -6, -6, -14,
    -- layer=1 filter=28 channel=48
    -3, -3, 3, 6, -6, 6, -6, 6, 7,
    -- layer=1 filter=28 channel=49
    0, -6, 0, -7, -16, 0, -8, -16, -15,
    -- layer=1 filter=28 channel=50
    -1, -8, -2, 5, -7, 4, 4, 7, -5,
    -- layer=1 filter=28 channel=51
    -1, -13, -11, -7, -10, 0, 0, -2, -3,
    -- layer=1 filter=28 channel=52
    11, 10, -5, -9, 0, 7, -1, 11, -8,
    -- layer=1 filter=28 channel=53
    -10, 6, 5, -11, -10, -9, 1, 6, 8,
    -- layer=1 filter=28 channel=54
    4, -3, -6, -12, -12, -5, -10, 0, -13,
    -- layer=1 filter=28 channel=55
    -7, -9, 6, -8, -10, -4, -15, -11, 0,
    -- layer=1 filter=28 channel=56
    4, 9, 2, -4, 2, 3, 0, -6, -8,
    -- layer=1 filter=28 channel=57
    4, -14, -17, -13, -15, -9, -5, -6, 1,
    -- layer=1 filter=28 channel=58
    -1, -6, -8, 3, 0, -16, -16, -12, 3,
    -- layer=1 filter=28 channel=59
    6, 1, 4, 2, -11, -3, -9, -4, -4,
    -- layer=1 filter=28 channel=60
    5, 3, -5, 5, 11, -1, 6, 3, -8,
    -- layer=1 filter=28 channel=61
    0, 1, -1, 8, 2, -9, -9, 0, 7,
    -- layer=1 filter=28 channel=62
    -16, -15, -15, 1, -4, -18, -7, -2, -7,
    -- layer=1 filter=28 channel=63
    -2, 0, 0, 7, -7, 3, -12, -5, 4,
    -- layer=1 filter=28 channel=64
    -12, 0, -3, -12, -5, -1, -10, -8, -3,
    -- layer=1 filter=28 channel=65
    6, -10, 3, -5, 4, -1, -4, -2, 7,
    -- layer=1 filter=28 channel=66
    -4, 0, 0, 3, -6, -1, -8, -3, -4,
    -- layer=1 filter=28 channel=67
    0, 5, 0, -13, -7, -7, 2, -5, 5,
    -- layer=1 filter=28 channel=68
    -5, 3, -5, -12, 4, 1, 5, -8, 3,
    -- layer=1 filter=28 channel=69
    -7, -12, -16, -9, -12, -2, -2, -8, -1,
    -- layer=1 filter=28 channel=70
    8, 2, -10, 9, -11, -7, -4, -1, -1,
    -- layer=1 filter=28 channel=71
    4, 5, -9, -1, -3, -4, -4, 6, 0,
    -- layer=1 filter=28 channel=72
    -9, 7, -5, 1, -8, -6, 9, 8, 8,
    -- layer=1 filter=28 channel=73
    8, 4, -1, -2, 1, -2, -3, 1, -8,
    -- layer=1 filter=28 channel=74
    4, 2, 0, 4, -3, -6, -2, -12, -2,
    -- layer=1 filter=28 channel=75
    -10, 4, 26, -6, -7, -9, -8, -6, -5,
    -- layer=1 filter=28 channel=76
    0, -5, -6, 2, -7, -7, -2, 3, -11,
    -- layer=1 filter=28 channel=77
    5, 2, 5, 4, -9, -5, 4, -11, 5,
    -- layer=1 filter=28 channel=78
    7, 3, -8, -11, -4, 5, -10, 5, -9,
    -- layer=1 filter=28 channel=79
    -4, 6, -7, 0, 6, -1, 3, -9, -8,
    -- layer=1 filter=28 channel=80
    -2, 1, 8, -1, 8, -7, 5, 5, -11,
    -- layer=1 filter=28 channel=81
    5, -6, -7, -10, 0, -2, 5, -7, -11,
    -- layer=1 filter=28 channel=82
    5, 3, 0, -5, -6, -11, -8, 5, -7,
    -- layer=1 filter=28 channel=83
    -4, 5, 3, -1, -6, -12, 7, 0, 2,
    -- layer=1 filter=28 channel=84
    -2, 4, -10, -1, -7, 2, -4, 0, -7,
    -- layer=1 filter=28 channel=85
    0, 4, -5, 7, -2, -3, -7, 5, 8,
    -- layer=1 filter=28 channel=86
    4, -8, -9, 2, -9, -3, -2, -5, -8,
    -- layer=1 filter=28 channel=87
    -3, -12, -9, 0, 4, 8, -11, -5, -4,
    -- layer=1 filter=28 channel=88
    -16, -14, -8, 3, 2, -12, -14, -10, -5,
    -- layer=1 filter=28 channel=89
    -8, -6, 4, -4, 1, -14, -10, -4, -3,
    -- layer=1 filter=28 channel=90
    7, -4, 0, -7, 4, 5, -9, -1, 1,
    -- layer=1 filter=28 channel=91
    2, -7, -13, 0, -7, 0, -8, -17, -3,
    -- layer=1 filter=28 channel=92
    0, -8, -2, -7, -5, -6, -11, 5, -2,
    -- layer=1 filter=28 channel=93
    0, 3, -4, -13, -1, -5, 5, -10, 1,
    -- layer=1 filter=28 channel=94
    -2, 2, -8, -8, -11, -7, 3, -5, -3,
    -- layer=1 filter=28 channel=95
    5, 3, 1, -12, 5, 0, 3, -6, 1,
    -- layer=1 filter=28 channel=96
    7, 1, -11, -3, 1, -7, 2, 0, 0,
    -- layer=1 filter=28 channel=97
    -12, 0, 5, -3, -6, -2, 3, 4, -1,
    -- layer=1 filter=28 channel=98
    -9, 0, 1, -7, -13, 1, -2, -13, -4,
    -- layer=1 filter=28 channel=99
    0, 3, 5, -10, -5, -2, -2, 7, -7,
    -- layer=1 filter=28 channel=100
    2, -7, -11, -3, 7, -10, 0, -2, -3,
    -- layer=1 filter=28 channel=101
    -1, 0, -4, -5, -11, 0, -4, 1, 1,
    -- layer=1 filter=28 channel=102
    0, -2, -12, -9, -1, -4, 7, 5, -10,
    -- layer=1 filter=28 channel=103
    -5, 3, -4, -13, -9, -9, -8, 0, 1,
    -- layer=1 filter=28 channel=104
    1, 2, 0, 6, -9, 2, -11, 3, 8,
    -- layer=1 filter=28 channel=105
    -5, 5, 0, 0, 3, 0, 5, 6, 2,
    -- layer=1 filter=28 channel=106
    -2, -18, -18, -16, -1, -6, -4, -12, -3,
    -- layer=1 filter=28 channel=107
    1, -9, -2, -2, -4, 0, 8, -7, -1,
    -- layer=1 filter=28 channel=108
    -2, -8, -19, -2, -13, -21, 12, -4, -4,
    -- layer=1 filter=28 channel=109
    -1, -4, -2, 2, 9, -3, 7, -7, 1,
    -- layer=1 filter=28 channel=110
    -1, 1, -9, -2, -5, -3, 2, -10, -10,
    -- layer=1 filter=28 channel=111
    -2, -8, 5, 2, -13, -12, 5, -6, -8,
    -- layer=1 filter=28 channel=112
    8, -11, 4, -5, 3, -10, 0, 0, 5,
    -- layer=1 filter=28 channel=113
    -12, 0, -1, -5, -14, -8, -6, -5, -8,
    -- layer=1 filter=28 channel=114
    -1, 0, 6, 1, -2, -4, -10, -11, 1,
    -- layer=1 filter=28 channel=115
    0, 6, 7, -1, -12, 4, -7, -7, 1,
    -- layer=1 filter=28 channel=116
    -5, 1, -8, -9, -4, -2, 2, -7, 3,
    -- layer=1 filter=28 channel=117
    4, 0, -9, -8, -7, 5, -13, -8, 0,
    -- layer=1 filter=28 channel=118
    -8, -4, 2, -9, 2, -2, -8, -9, -9,
    -- layer=1 filter=28 channel=119
    -15, -4, -9, -2, -11, 4, -1, 3, -15,
    -- layer=1 filter=28 channel=120
    0, -13, -14, -13, -9, 2, -3, -16, -10,
    -- layer=1 filter=28 channel=121
    6, 2, 3, -14, 3, -4, -2, 1, -8,
    -- layer=1 filter=28 channel=122
    -2, 0, -4, 7, -9, -6, 6, -10, 10,
    -- layer=1 filter=28 channel=123
    -7, -4, 7, -4, -8, -8, 2, -10, -2,
    -- layer=1 filter=28 channel=124
    6, 1, 4, -8, 2, 7, 9, 4, -5,
    -- layer=1 filter=28 channel=125
    3, 0, -7, 7, 3, 0, 0, -1, 4,
    -- layer=1 filter=28 channel=126
    6, 2, 5, -6, 6, 1, 6, -2, -3,
    -- layer=1 filter=28 channel=127
    -17, 0, 9, 0, -6, -8, -12, -5, 0,
    -- layer=1 filter=29 channel=0
    8, 1, 1, 6, 3, 8, 2, -11, 0,
    -- layer=1 filter=29 channel=1
    -6, -9, 3, 23, 12, 18, 0, -4, -16,
    -- layer=1 filter=29 channel=2
    -14, -24, -7, -1, -3, -1, 20, -17, -13,
    -- layer=1 filter=29 channel=3
    -2, 7, 3, 2, -11, -1, 2, -10, 12,
    -- layer=1 filter=29 channel=4
    -2, 3, 0, 2, 7, 4, 4, 12, 16,
    -- layer=1 filter=29 channel=5
    -4, 1, -13, 32, 15, 11, -3, -16, -28,
    -- layer=1 filter=29 channel=6
    15, 23, 11, -10, 0, 0, 5, 1, 14,
    -- layer=1 filter=29 channel=7
    11, -13, 13, 8, 7, -5, 7, 22, 22,
    -- layer=1 filter=29 channel=8
    -10, -28, -15, 8, -6, 3, -3, -27, -29,
    -- layer=1 filter=29 channel=9
    29, 36, 32, 31, -17, 20, 12, 8, 23,
    -- layer=1 filter=29 channel=10
    14, -4, 13, 5, 14, -2, -2, 26, 27,
    -- layer=1 filter=29 channel=11
    7, 10, -11, -13, -7, -10, -4, -1, 0,
    -- layer=1 filter=29 channel=12
    28, 35, 9, 20, 4, -41, 46, 25, 48,
    -- layer=1 filter=29 channel=13
    5, 6, 5, -12, 9, -8, -3, -5, -11,
    -- layer=1 filter=29 channel=14
    -11, -39, 8, 0, 13, -1, 9, 5, 16,
    -- layer=1 filter=29 channel=15
    0, -6, -11, 17, 14, 1, 31, 5, -3,
    -- layer=1 filter=29 channel=16
    4, -3, -6, 16, 0, 3, -2, -29, -6,
    -- layer=1 filter=29 channel=17
    -12, 14, -6, -17, -1, -8, -19, -13, -22,
    -- layer=1 filter=29 channel=18
    17, 13, 2, 15, 9, -9, 0, 9, 22,
    -- layer=1 filter=29 channel=19
    48, 59, 34, 59, 39, 17, 31, 53, 44,
    -- layer=1 filter=29 channel=20
    -9, 3, 6, -4, -9, -10, -9, -14, -18,
    -- layer=1 filter=29 channel=21
    6, 10, 8, 1, 2, 19, -10, -15, -6,
    -- layer=1 filter=29 channel=22
    1, 12, -14, -7, 5, 3, -12, -13, -36,
    -- layer=1 filter=29 channel=23
    25, 21, 13, 18, -29, 24, 2, 14, 7,
    -- layer=1 filter=29 channel=24
    1, 11, 4, -1, -2, -8, -10, -21, -20,
    -- layer=1 filter=29 channel=25
    3, -7, 13, 6, 9, 8, -4, 12, 8,
    -- layer=1 filter=29 channel=26
    -8, 2, -2, -2, 4, 9, -8, -7, -13,
    -- layer=1 filter=29 channel=27
    43, 41, 36, 12, 33, 29, 7, 1, 7,
    -- layer=1 filter=29 channel=28
    -1, -6, 2, -1, 20, -1, -3, 9, 18,
    -- layer=1 filter=29 channel=29
    21, 21, 34, 3, 2, 20, 8, 1, 12,
    -- layer=1 filter=29 channel=30
    4, 7, 5, 29, 4, -4, 16, 29, 27,
    -- layer=1 filter=29 channel=31
    29, 29, 19, 16, 3, -16, 9, 25, 19,
    -- layer=1 filter=29 channel=32
    6, 17, 3, 7, -12, 25, 0, 25, 15,
    -- layer=1 filter=29 channel=33
    27, 23, 18, 13, 3, 2, 18, 2, -16,
    -- layer=1 filter=29 channel=34
    10, 19, 16, -4, 25, -10, 5, 12, -9,
    -- layer=1 filter=29 channel=35
    -12, 0, -10, 2, -1, -8, 1, 4, -8,
    -- layer=1 filter=29 channel=36
    1, 8, 0, -9, 3, 0, -22, -21, -2,
    -- layer=1 filter=29 channel=37
    21, 24, 0, 21, 22, 0, 10, -16, -6,
    -- layer=1 filter=29 channel=38
    4, -3, -4, 0, 14, 9, -2, -8, -2,
    -- layer=1 filter=29 channel=39
    3, 1, 6, 14, 9, 9, -5, -25, -20,
    -- layer=1 filter=29 channel=40
    22, 15, 4, 7, 21, -7, 16, 16, -2,
    -- layer=1 filter=29 channel=41
    -9, 16, -6, 22, -5, 20, -1, 12, 15,
    -- layer=1 filter=29 channel=42
    -35, -14, -28, -2, -8, -6, 25, 9, 9,
    -- layer=1 filter=29 channel=43
    9, -7, -19, 13, 0, 15, 5, -1, -17,
    -- layer=1 filter=29 channel=44
    -5, 12, -13, -10, -15, 16, -2, 16, 2,
    -- layer=1 filter=29 channel=45
    -8, 7, -6, 4, 13, 14, 5, -6, -11,
    -- layer=1 filter=29 channel=46
    20, 50, 36, 27, 32, 8, 42, 72, 32,
    -- layer=1 filter=29 channel=47
    14, 15, 13, 34, 7, 40, 0, 3, 36,
    -- layer=1 filter=29 channel=48
    1, 7, 9, -9, 9, 2, -16, -16, -4,
    -- layer=1 filter=29 channel=49
    7, 10, 9, 0, 8, 12, 6, -7, -8,
    -- layer=1 filter=29 channel=50
    -4, 8, 11, -7, -13, -6, -5, 0, -15,
    -- layer=1 filter=29 channel=51
    6, 0, 6, 8, -2, 4, -6, 6, -4,
    -- layer=1 filter=29 channel=52
    -6, -7, 8, -4, -3, -7, 17, 17, 9,
    -- layer=1 filter=29 channel=53
    -26, -13, -16, -16, 2, -13, -18, -1, -8,
    -- layer=1 filter=29 channel=54
    0, 9, 0, 14, -7, 5, 8, 3, 26,
    -- layer=1 filter=29 channel=55
    4, -1, 1, -2, -19, -12, -18, -15, 3,
    -- layer=1 filter=29 channel=56
    -3, -4, -10, 8, 10, 11, 10, 1, 4,
    -- layer=1 filter=29 channel=57
    5, -16, 21, -7, -1, -5, 2, 8, 19,
    -- layer=1 filter=29 channel=58
    32, 11, 37, 39, 8, 20, 13, 27, 34,
    -- layer=1 filter=29 channel=59
    -6, 13, 0, 3, 5, 6, -4, 4, 1,
    -- layer=1 filter=29 channel=60
    17, 1, 3, 20, 13, 0, 20, 2, 9,
    -- layer=1 filter=29 channel=61
    4, 5, -8, -5, 4, 4, 3, 8, -2,
    -- layer=1 filter=29 channel=62
    12, -12, -25, 11, 18, 3, 11, -29, -6,
    -- layer=1 filter=29 channel=63
    0, -6, -12, -6, -2, -2, -18, -9, -6,
    -- layer=1 filter=29 channel=64
    -1, -6, 4, -3, 7, -3, -1, -11, -17,
    -- layer=1 filter=29 channel=65
    7, 9, 21, 2, 11, 4, -17, -23, -10,
    -- layer=1 filter=29 channel=66
    11, 5, 10, -1, -12, -3, -14, -7, -9,
    -- layer=1 filter=29 channel=67
    37, 36, 21, 44, 31, 18, 17, 13, 31,
    -- layer=1 filter=29 channel=68
    11, 18, 3, 0, -5, 16, 21, 12, 18,
    -- layer=1 filter=29 channel=69
    -6, -9, -19, 9, 17, 8, 2, -10, -19,
    -- layer=1 filter=29 channel=70
    48, 34, 16, 26, 25, 8, 32, 40, 30,
    -- layer=1 filter=29 channel=71
    10, 5, 20, -10, 2, 18, -15, -27, -3,
    -- layer=1 filter=29 channel=72
    9, 23, 7, 41, 5, 18, 29, 33, 12,
    -- layer=1 filter=29 channel=73
    0, -2, -4, 4, -8, 13, 5, -1, 0,
    -- layer=1 filter=29 channel=74
    12, 11, 1, -3, 0, 22, -4, 23, 24,
    -- layer=1 filter=29 channel=75
    1, 15, 15, 15, 18, 4, 19, 26, 38,
    -- layer=1 filter=29 channel=76
    2, 12, 5, 6, -2, 17, -2, 0, 7,
    -- layer=1 filter=29 channel=77
    -2, 22, 21, -9, 12, 15, -24, -10, -3,
    -- layer=1 filter=29 channel=78
    10, 15, 18, 5, 14, 4, 0, -3, 13,
    -- layer=1 filter=29 channel=79
    -7, 4, 0, 0, 6, -14, -7, -22, -11,
    -- layer=1 filter=29 channel=80
    9, 9, 2, 1, 11, 11, -1, 6, 11,
    -- layer=1 filter=29 channel=81
    17, 25, 18, 2, 13, 17, -21, -31, -12,
    -- layer=1 filter=29 channel=82
    -1, 16, 1, -8, -10, 6, -12, -10, -16,
    -- layer=1 filter=29 channel=83
    -11, -6, -15, -17, 10, -8, -9, -20, -3,
    -- layer=1 filter=29 channel=84
    43, 36, 6, 29, 24, 5, 17, 22, 35,
    -- layer=1 filter=29 channel=85
    -3, 15, 4, 35, 0, 17, -19, 11, 18,
    -- layer=1 filter=29 channel=86
    7, 4, 7, -11, 2, -5, -9, -21, -27,
    -- layer=1 filter=29 channel=87
    14, 27, 24, 41, 21, 4, 1, 52, 30,
    -- layer=1 filter=29 channel=88
    16, 14, 9, 19, 2, 1, -7, -9, 1,
    -- layer=1 filter=29 channel=89
    12, 18, 14, 6, 0, 16, -10, -9, -12,
    -- layer=1 filter=29 channel=90
    -15, 13, -4, -5, 11, 22, 12, 13, 9,
    -- layer=1 filter=29 channel=91
    -1, 1, -4, -2, 2, -10, -16, 3, -9,
    -- layer=1 filter=29 channel=92
    -31, 27, -1, -17, -6, 25, -8, -3, 24,
    -- layer=1 filter=29 channel=93
    -8, -3, -4, -14, 1, -4, -18, -22, -15,
    -- layer=1 filter=29 channel=94
    -1, -6, -2, 4, -7, 4, -17, -8, -15,
    -- layer=1 filter=29 channel=95
    32, 17, 4, 34, 14, 8, 31, 45, 39,
    -- layer=1 filter=29 channel=96
    2, 0, 1, -11, -9, -9, -5, -8, -10,
    -- layer=1 filter=29 channel=97
    0, 6, 7, -6, -3, -9, -22, -29, -25,
    -- layer=1 filter=29 channel=98
    -3, -11, -28, 3, 15, 2, -7, -18, -15,
    -- layer=1 filter=29 channel=99
    20, 11, 10, 7, 16, 22, 8, 24, 29,
    -- layer=1 filter=29 channel=100
    3, 5, 3, 1, -15, 16, -25, -7, 11,
    -- layer=1 filter=29 channel=101
    -6, 2, 5, 2, 0, -1, -9, -13, -9,
    -- layer=1 filter=29 channel=102
    -3, 0, -8, -16, -1, 0, -12, -10, -7,
    -- layer=1 filter=29 channel=103
    19, 14, 11, 6, 10, 6, 2, 6, 18,
    -- layer=1 filter=29 channel=104
    3, 4, 10, 17, 6, 12, 8, 3, 34,
    -- layer=1 filter=29 channel=105
    14, 11, 12, -10, -3, -9, -15, -7, -7,
    -- layer=1 filter=29 channel=106
    2, 13, -4, -4, -8, -6, 4, -12, -16,
    -- layer=1 filter=29 channel=107
    -15, -12, 3, -9, -18, -7, -1, 10, -15,
    -- layer=1 filter=29 channel=108
    -11, 3, -4, -5, 0, 4, 20, 3, 4,
    -- layer=1 filter=29 channel=109
    2, -1, -3, -5, -5, 11, 7, 5, 7,
    -- layer=1 filter=29 channel=110
    0, 0, 5, 11, 0, -2, -8, -10, 7,
    -- layer=1 filter=29 channel=111
    11, 13, 8, 18, 7, 4, 18, 33, 31,
    -- layer=1 filter=29 channel=112
    35, 9, -9, 1, 22, -21, 32, 16, 42,
    -- layer=1 filter=29 channel=113
    12, 21, 3, 11, 19, 5, -14, 11, -27,
    -- layer=1 filter=29 channel=114
    -13, -19, -14, 2, 15, -11, -3, -28, -17,
    -- layer=1 filter=29 channel=115
    7, 3, 8, -14, -4, -11, -27, -11, -8,
    -- layer=1 filter=29 channel=116
    1, -2, 7, 6, -7, -7, -9, -3, -1,
    -- layer=1 filter=29 channel=117
    52, 7, 39, 63, 63, 18, 40, 56, 72,
    -- layer=1 filter=29 channel=118
    12, 24, -2, 12, -1, -8, -3, 13, 13,
    -- layer=1 filter=29 channel=119
    0, 21, 0, 0, -1, 16, 12, 21, 25,
    -- layer=1 filter=29 channel=120
    -4, 5, 0, -4, 6, 7, -6, -13, 0,
    -- layer=1 filter=29 channel=121
    -9, 3, 10, -10, -13, -2, 5, 20, 28,
    -- layer=1 filter=29 channel=122
    8, 0, -6, 3, -8, -2, 3, -10, 6,
    -- layer=1 filter=29 channel=123
    -6, 8, -5, 0, -2, -6, -25, 4, -1,
    -- layer=1 filter=29 channel=124
    0, 6, 14, 4, 11, 15, 7, 6, 9,
    -- layer=1 filter=29 channel=125
    10, 21, 28, 11, 41, 11, 0, 25, 18,
    -- layer=1 filter=29 channel=126
    16, 20, -22, 5, 10, 18, 31, 20, 8,
    -- layer=1 filter=29 channel=127
    12, 15, -9, 3, 11, -6, 10, 31, 36,
    -- layer=1 filter=30 channel=0
    -12, -3, -5, 0, -11, -6, -7, 2, 6,
    -- layer=1 filter=30 channel=1
    -6, -4, -2, -1, -4, 0, -5, -11, -4,
    -- layer=1 filter=30 channel=2
    -5, 4, -11, -10, -13, -7, -14, -12, -2,
    -- layer=1 filter=30 channel=3
    -1, 9, -6, -1, 8, 2, 7, -7, 0,
    -- layer=1 filter=30 channel=4
    7, -11, 6, 2, -8, 1, 6, -10, 3,
    -- layer=1 filter=30 channel=5
    -7, 10, -1, 0, -10, 0, -3, 4, -2,
    -- layer=1 filter=30 channel=6
    5, -2, 2, -2, 2, -2, -3, 4, -1,
    -- layer=1 filter=30 channel=7
    -1, 14, 8, -1, 17, -7, -1, 10, 0,
    -- layer=1 filter=30 channel=8
    -10, 1, 5, 5, -9, 0, -2, 2, 5,
    -- layer=1 filter=30 channel=9
    0, -5, -3, -6, 9, -8, -5, -6, -11,
    -- layer=1 filter=30 channel=10
    7, 2, 3, 11, -4, -18, 4, 4, -3,
    -- layer=1 filter=30 channel=11
    -1, -9, 0, 4, -1, -7, -8, 1, -3,
    -- layer=1 filter=30 channel=12
    -10, 3, 8, 0, 0, 4, -12, -6, 6,
    -- layer=1 filter=30 channel=13
    4, -13, -10, -2, -3, 1, -6, -12, -7,
    -- layer=1 filter=30 channel=14
    -11, -2, 3, 6, 6, -6, 2, 0, -5,
    -- layer=1 filter=30 channel=15
    -8, 9, -3, 6, -9, 2, -6, 8, 9,
    -- layer=1 filter=30 channel=16
    -8, 0, -11, -12, -11, -14, -6, 5, -1,
    -- layer=1 filter=30 channel=17
    -8, -6, 4, -8, -4, -6, 3, -13, -10,
    -- layer=1 filter=30 channel=18
    4, -2, -4, 2, -1, -6, -2, -5, -8,
    -- layer=1 filter=30 channel=19
    5, 7, 6, -10, -2, -3, -1, 8, -11,
    -- layer=1 filter=30 channel=20
    -11, 5, -12, 2, 0, 4, -8, -7, -12,
    -- layer=1 filter=30 channel=21
    4, -7, 3, 4, 7, 3, -13, -6, 1,
    -- layer=1 filter=30 channel=22
    5, -6, -10, 8, -9, -1, 4, 3, -13,
    -- layer=1 filter=30 channel=23
    0, -4, -12, -2, 0, 0, -11, -11, 7,
    -- layer=1 filter=30 channel=24
    7, -6, -6, -14, -13, 6, -5, 3, -5,
    -- layer=1 filter=30 channel=25
    7, 0, -5, -6, 7, -1, 3, 13, -1,
    -- layer=1 filter=30 channel=26
    0, 4, -4, -3, 4, -7, 0, 3, 3,
    -- layer=1 filter=30 channel=27
    3, -10, -1, -10, 2, -14, 0, 0, -7,
    -- layer=1 filter=30 channel=28
    -4, 5, -1, -1, 1, -10, -10, -12, -5,
    -- layer=1 filter=30 channel=29
    0, 0, 1, -4, -2, 0, 1, 6, 7,
    -- layer=1 filter=30 channel=30
    1, 7, -6, 8, -10, 9, 4, 5, -7,
    -- layer=1 filter=30 channel=31
    -3, 3, 8, 0, -4, 4, 13, 6, -14,
    -- layer=1 filter=30 channel=32
    -4, -10, -13, 2, -12, 3, -7, -14, -2,
    -- layer=1 filter=30 channel=33
    -2, 6, -4, 5, -6, -8, -4, 2, -4,
    -- layer=1 filter=30 channel=34
    1, -9, -6, -11, -5, -10, 5, 1, 7,
    -- layer=1 filter=30 channel=35
    0, 6, -6, -4, -2, -1, 5, -3, 0,
    -- layer=1 filter=30 channel=36
    5, -6, -1, 4, -7, -5, 0, -5, 2,
    -- layer=1 filter=30 channel=37
    -6, 9, -6, -5, -14, 0, -2, -11, -8,
    -- layer=1 filter=30 channel=38
    -5, -2, 0, -8, 3, -14, -3, 0, -11,
    -- layer=1 filter=30 channel=39
    -6, 1, 0, -5, 3, -12, 6, -10, -8,
    -- layer=1 filter=30 channel=40
    -1, -9, -7, 6, -7, -14, 4, 1, -1,
    -- layer=1 filter=30 channel=41
    4, -9, -10, -5, -6, 7, 0, -6, -4,
    -- layer=1 filter=30 channel=42
    9, 0, -1, -2, -1, 0, -5, -15, -9,
    -- layer=1 filter=30 channel=43
    5, -8, 2, -11, -9, -10, 1, -2, -10,
    -- layer=1 filter=30 channel=44
    5, 2, 6, 7, -8, -7, 8, 5, -11,
    -- layer=1 filter=30 channel=45
    -2, -5, 0, -11, -8, -2, -6, -6, 6,
    -- layer=1 filter=30 channel=46
    8, 2, 0, -4, 0, -11, -2, 2, -8,
    -- layer=1 filter=30 channel=47
    7, -11, -6, -6, -12, -8, -9, -13, 6,
    -- layer=1 filter=30 channel=48
    3, -5, -14, 0, -3, -7, 2, 5, 4,
    -- layer=1 filter=30 channel=49
    -1, -5, -13, -5, -11, -13, -4, 1, -9,
    -- layer=1 filter=30 channel=50
    -12, -6, -4, 6, 1, 10, 0, 6, 3,
    -- layer=1 filter=30 channel=51
    -13, -12, 5, -7, 4, -2, -1, -13, 4,
    -- layer=1 filter=30 channel=52
    12, 0, -4, 14, 2, 0, 5, -13, -2,
    -- layer=1 filter=30 channel=53
    5, 8, 0, -5, 3, -5, -8, 7, -8,
    -- layer=1 filter=30 channel=54
    4, -2, 4, -4, 10, -2, 3, -9, 7,
    -- layer=1 filter=30 channel=55
    -7, 2, -11, -3, -5, 0, -7, -6, 7,
    -- layer=1 filter=30 channel=56
    -7, 0, -2, 7, -8, -4, -5, 6, -4,
    -- layer=1 filter=30 channel=57
    -1, 2, -12, 8, 4, -10, 1, 5, -5,
    -- layer=1 filter=30 channel=58
    -2, -5, 4, -6, -1, -3, -4, 5, -7,
    -- layer=1 filter=30 channel=59
    2, 8, -6, 6, -7, -9, 1, -7, 0,
    -- layer=1 filter=30 channel=60
    -7, 9, 8, 0, 7, 10, -4, 6, -3,
    -- layer=1 filter=30 channel=61
    4, 8, -3, -1, 10, -8, 2, 4, 5,
    -- layer=1 filter=30 channel=62
    5, 6, -2, 8, -11, -4, 8, -5, 8,
    -- layer=1 filter=30 channel=63
    2, -8, 3, -4, 0, -10, 2, 0, 2,
    -- layer=1 filter=30 channel=64
    1, -10, 0, -6, -12, -13, -14, -1, -1,
    -- layer=1 filter=30 channel=65
    -13, 2, -12, -6, 5, 4, -2, -13, 4,
    -- layer=1 filter=30 channel=66
    0, 0, 1, -11, -8, 5, -12, 3, -2,
    -- layer=1 filter=30 channel=67
    3, 3, -14, -4, -11, 6, -5, -7, -14,
    -- layer=1 filter=30 channel=68
    3, -13, 6, -2, -2, 0, -13, -4, 7,
    -- layer=1 filter=30 channel=69
    7, 2, -13, -10, -8, 6, -9, -16, 1,
    -- layer=1 filter=30 channel=70
    -9, -5, -9, 2, 0, -6, -2, 6, 4,
    -- layer=1 filter=30 channel=71
    -15, -7, 2, -9, 0, -9, -5, 1, -13,
    -- layer=1 filter=30 channel=72
    -2, 2, -3, -13, 2, -9, -7, -4, -2,
    -- layer=1 filter=30 channel=73
    -6, -1, -5, 11, -2, -4, -11, 7, -3,
    -- layer=1 filter=30 channel=74
    -5, 8, -8, 2, -8, -7, 0, -11, 3,
    -- layer=1 filter=30 channel=75
    -1, 5, -3, 0, 9, 2, 8, -2, -12,
    -- layer=1 filter=30 channel=76
    -11, -12, -1, -11, -8, -3, -12, 2, -12,
    -- layer=1 filter=30 channel=77
    -11, 5, -4, -11, 4, 3, -10, 2, -8,
    -- layer=1 filter=30 channel=78
    -1, 6, -5, -12, -2, 4, 2, -10, -2,
    -- layer=1 filter=30 channel=79
    -4, 8, 4, -7, 5, -14, -3, -6, -6,
    -- layer=1 filter=30 channel=80
    10, -4, 0, 6, -7, 2, 2, 4, -9,
    -- layer=1 filter=30 channel=81
    -4, -8, 2, -13, -3, 3, 5, -1, -8,
    -- layer=1 filter=30 channel=82
    0, -1, 3, -15, 2, 1, -2, 0, 1,
    -- layer=1 filter=30 channel=83
    -6, -11, 3, 1, 1, -2, 4, -11, -3,
    -- layer=1 filter=30 channel=84
    -9, -6, -7, -9, -8, 8, -1, 12, 5,
    -- layer=1 filter=30 channel=85
    -3, -7, -3, -6, 0, -11, 3, -9, -3,
    -- layer=1 filter=30 channel=86
    6, 8, -5, 7, 1, 4, 7, 3, -13,
    -- layer=1 filter=30 channel=87
    0, -6, 7, 6, -6, 7, 6, -2, 1,
    -- layer=1 filter=30 channel=88
    0, 2, 0, 3, -6, 4, -9, -7, 5,
    -- layer=1 filter=30 channel=89
    -9, -4, -7, -14, 0, -3, -8, 0, 3,
    -- layer=1 filter=30 channel=90
    -1, -4, -1, -11, -5, 6, -2, 5, -2,
    -- layer=1 filter=30 channel=91
    -3, -5, -12, -6, -9, 0, -8, -14, -10,
    -- layer=1 filter=30 channel=92
    5, -4, 3, 4, 8, -5, 2, -5, -10,
    -- layer=1 filter=30 channel=93
    -16, -11, 1, -6, -5, 2, -2, -8, -1,
    -- layer=1 filter=30 channel=94
    -6, -9, -6, -14, -7, 0, -1, -4, -12,
    -- layer=1 filter=30 channel=95
    2, 3, -7, 0, -8, -5, -2, 0, 1,
    -- layer=1 filter=30 channel=96
    -1, -12, 5, 1, -10, 5, -9, 2, -9,
    -- layer=1 filter=30 channel=97
    0, -7, 3, 2, 5, -4, -13, -9, -5,
    -- layer=1 filter=30 channel=98
    -9, 2, 5, -6, -5, 0, 3, -1, 7,
    -- layer=1 filter=30 channel=99
    -7, 0, 0, -7, -9, 3, 3, 0, 1,
    -- layer=1 filter=30 channel=100
    -11, 4, 2, -11, -3, -12, -8, 0, -10,
    -- layer=1 filter=30 channel=101
    -4, 4, -4, -8, -6, -1, -8, 0, -5,
    -- layer=1 filter=30 channel=102
    -12, -6, 0, -4, 4, 4, -3, 0, 2,
    -- layer=1 filter=30 channel=103
    1, 6, -6, 10, 7, 6, 3, -8, 8,
    -- layer=1 filter=30 channel=104
    -2, -11, 3, 8, 0, 0, 0, -2, -9,
    -- layer=1 filter=30 channel=105
    -4, -2, 0, -9, 3, -11, 4, 4, -2,
    -- layer=1 filter=30 channel=106
    -5, -15, 0, -7, -10, 1, -4, -5, -14,
    -- layer=1 filter=30 channel=107
    -2, 1, -5, 8, 0, -10, -7, 2, 0,
    -- layer=1 filter=30 channel=108
    -3, 5, -9, -10, -11, 5, -13, -6, 3,
    -- layer=1 filter=30 channel=109
    8, -3, -3, -7, 6, -3, -6, 5, 9,
    -- layer=1 filter=30 channel=110
    1, -9, -12, -10, -5, -4, 2, -10, -1,
    -- layer=1 filter=30 channel=111
    2, -11, -9, -2, 0, 9, -3, -1, 7,
    -- layer=1 filter=30 channel=112
    -3, 2, -3, -10, -3, 1, -5, 8, -6,
    -- layer=1 filter=30 channel=113
    8, -1, 7, 1, 4, -15, -1, 4, -10,
    -- layer=1 filter=30 channel=114
    -9, -8, -10, -6, 0, 7, -9, -7, -2,
    -- layer=1 filter=30 channel=115
    -2, -2, -13, -13, 6, -7, 5, 5, -6,
    -- layer=1 filter=30 channel=116
    10, -3, 5, 1, -8, -2, -3, -8, 7,
    -- layer=1 filter=30 channel=117
    -4, -11, -1, -10, 4, 4, 8, -8, -5,
    -- layer=1 filter=30 channel=118
    -10, -10, -7, -1, -2, -2, -7, 7, -10,
    -- layer=1 filter=30 channel=119
    -7, -4, 3, -3, -7, -8, -2, -3, -7,
    -- layer=1 filter=30 channel=120
    -2, 7, 3, -6, 6, -14, -10, 4, -11,
    -- layer=1 filter=30 channel=121
    -4, 7, -10, 6, -1, -8, 8, -7, -14,
    -- layer=1 filter=30 channel=122
    -9, -7, -3, -4, -5, 9, 9, -4, -5,
    -- layer=1 filter=30 channel=123
    -12, -11, 1, 7, -9, -4, 3, -11, 0,
    -- layer=1 filter=30 channel=124
    5, 4, -2, -6, -3, -10, 0, -3, 6,
    -- layer=1 filter=30 channel=125
    -10, -3, -10, -1, 0, -8, -6, -5, -11,
    -- layer=1 filter=30 channel=126
    3, 6, 2, -1, 3, 1, 0, -1, -11,
    -- layer=1 filter=30 channel=127
    -7, -8, -14, -5, -7, -4, 0, 13, 7,
    -- layer=1 filter=31 channel=0
    -22, -36, -30, 13, -26, -40, 22, -10, -9,
    -- layer=1 filter=31 channel=1
    5, 11, -38, 22, 5, -3, 9, 11, 19,
    -- layer=1 filter=31 channel=2
    -2, 38, 50, -2, 37, 62, -14, 36, 58,
    -- layer=1 filter=31 channel=3
    7, -3, -9, -12, 6, 1, 0, -3, 21,
    -- layer=1 filter=31 channel=4
    10, 0, 13, -4, -17, -32, 5, -14, 15,
    -- layer=1 filter=31 channel=5
    24, 20, -26, 30, 43, 17, 14, 13, 29,
    -- layer=1 filter=31 channel=6
    -38, -39, 18, -61, -68, -8, 3, -25, -20,
    -- layer=1 filter=31 channel=7
    -61, -45, -17, -87, -124, -37, -35, -127, -94,
    -- layer=1 filter=31 channel=8
    4, 21, -15, 30, 12, 2, -2, 17, 19,
    -- layer=1 filter=31 channel=9
    -15, -44, 13, -35, -5, -22, -9, -8, -30,
    -- layer=1 filter=31 channel=10
    -89, -83, -17, -64, -143, -51, -37, -127, -102,
    -- layer=1 filter=31 channel=11
    27, 7, 8, 28, -8, -22, 38, 13, -27,
    -- layer=1 filter=31 channel=12
    3, -46, 40, -67, -5, 71, -11, 21, -7,
    -- layer=1 filter=31 channel=13
    39, -9, -1, 29, 28, -4, 27, 9, 10,
    -- layer=1 filter=31 channel=14
    -2, 10, 4, -34, -8, 64, -24, -44, -43,
    -- layer=1 filter=31 channel=15
    37, 58, 0, 37, 54, 89, 36, 34, 29,
    -- layer=1 filter=31 channel=16
    12, 11, -7, 0, 20, 13, 21, 17, 13,
    -- layer=1 filter=31 channel=17
    23, -57, -53, 42, -14, -49, 25, 0, -20,
    -- layer=1 filter=31 channel=18
    18, 31, 19, -2, -26, 8, 8, 0, -24,
    -- layer=1 filter=31 channel=19
    -4, -49, -31, -64, -34, -19, -35, -56, -68,
    -- layer=1 filter=31 channel=20
    27, 11, -10, 20, 13, -9, 17, 0, -3,
    -- layer=1 filter=31 channel=21
    -13, -1, 11, 3, -6, 3, -2, 0, -4,
    -- layer=1 filter=31 channel=22
    9, 1, 3, 25, 23, -7, 5, -16, 8,
    -- layer=1 filter=31 channel=23
    -32, 20, -46, -56, 10, -23, -24, -50, -15,
    -- layer=1 filter=31 channel=24
    33, -5, 9, 35, 40, 21, 0, 22, 22,
    -- layer=1 filter=31 channel=25
    -76, -52, -29, -100, -88, -57, -68, -78, -34,
    -- layer=1 filter=31 channel=26
    58, -7, 4, 53, 43, -12, 34, 24, 24,
    -- layer=1 filter=31 channel=27
    5, 0, -7, -7, -7, 5, -3, -6, 8,
    -- layer=1 filter=31 channel=28
    -60, -96, -27, -99, -131, -53, -45, -107, -107,
    -- layer=1 filter=31 channel=29
    2, -20, -23, -12, -25, -36, -27, -40, -20,
    -- layer=1 filter=31 channel=30
    -4, -2, -11, -8, -35, 17, 27, 2, -42,
    -- layer=1 filter=31 channel=31
    7, 11, 21, -54, -4, 47, -5, -28, -32,
    -- layer=1 filter=31 channel=32
    51, 7, -1, 16, 27, -7, 19, 10, -7,
    -- layer=1 filter=31 channel=33
    13, 6, 36, -3, 6, 7, -27, -21, -7,
    -- layer=1 filter=31 channel=34
    -3, 26, 61, -5, -24, 8, -3, -16, -30,
    -- layer=1 filter=31 channel=35
    -5, 25, -56, -7, 6, 21, 20, 9, -4,
    -- layer=1 filter=31 channel=36
    28, -9, 4, 29, -16, -24, 41, 0, -22,
    -- layer=1 filter=31 channel=37
    1, 7, -24, 10, 15, 10, -11, -4, 35,
    -- layer=1 filter=31 channel=38
    16, -10, -1, -9, -6, 3, 0, 4, -1,
    -- layer=1 filter=31 channel=39
    -4, -32, -45, 32, -9, -18, 5, 0, -16,
    -- layer=1 filter=31 channel=40
    -5, -9, 25, -57, -54, -5, -15, -35, -33,
    -- layer=1 filter=31 channel=41
    19, -29, 24, -24, -9, -34, -14, -30, -52,
    -- layer=1 filter=31 channel=42
    3, 38, 50, -10, 43, 69, -10, 36, 67,
    -- layer=1 filter=31 channel=43
    -28, -4, -30, -18, -5, -21, 0, -18, 21,
    -- layer=1 filter=31 channel=44
    53, 2, -7, 39, 55, 0, 37, 12, 20,
    -- layer=1 filter=31 channel=45
    19, -3, -2, 24, 31, -5, 0, 0, 26,
    -- layer=1 filter=31 channel=46
    53, 17, 41, -31, 45, 83, -14, 25, 13,
    -- layer=1 filter=31 channel=47
    6, 33, -24, -27, -3, 25, -5, -36, -14,
    -- layer=1 filter=31 channel=48
    -25, -17, -8, -13, -9, -2, -10, -13, -24,
    -- layer=1 filter=31 channel=49
    0, 11, 21, -26, -20, 15, -27, -11, -4,
    -- layer=1 filter=31 channel=50
    10, -20, -5, -17, -24, -22, 6, 4, 28,
    -- layer=1 filter=31 channel=51
    -41, -17, 18, -25, -50, -23, -4, -31, -45,
    -- layer=1 filter=31 channel=52
    -20, -13, 3, 15, 42, 25, 4, -29, -9,
    -- layer=1 filter=31 channel=53
    -13, -5, -5, -20, 4, -5, -15, -3, -1,
    -- layer=1 filter=31 channel=54
    -65, -58, -42, -79, -75, -66, -74, -99, -20,
    -- layer=1 filter=31 channel=55
    33, 28, 31, 38, 14, 12, 43, 38, 32,
    -- layer=1 filter=31 channel=56
    1, 0, 5, 5, 0, -9, 0, 1, -4,
    -- layer=1 filter=31 channel=57
    -52, -28, -4, -61, -114, -31, -30, -97, -90,
    -- layer=1 filter=31 channel=58
    -133, -53, -64, -114, -130, -70, -106, -140, -71,
    -- layer=1 filter=31 channel=59
    -5, -4, -17, -16, -8, -15, -1, 10, 8,
    -- layer=1 filter=31 channel=60
    -36, -10, -55, 11, 7, 10, 2, 18, 0,
    -- layer=1 filter=31 channel=61
    5, 2, 0, -10, -4, -8, -5, 2, 0,
    -- layer=1 filter=31 channel=62
    11, 8, -8, 21, 28, 2, 4, 15, 37,
    -- layer=1 filter=31 channel=63
    19, 9, -2, -5, -16, -1, 36, 0, -10,
    -- layer=1 filter=31 channel=64
    -6, 21, 14, 1, 7, -9, -11, -16, -8,
    -- layer=1 filter=31 channel=65
    -13, -25, -11, -7, -15, -2, 0, -17, -24,
    -- layer=1 filter=31 channel=66
    -2, -14, -36, 16, -10, -38, 22, -4, -13,
    -- layer=1 filter=31 channel=67
    6, 53, 68, -12, 28, 70, 26, 63, 67,
    -- layer=1 filter=31 channel=68
    34, -29, -13, 24, 37, -31, 39, -2, -5,
    -- layer=1 filter=31 channel=69
    54, 59, -1, 63, 80, 42, 19, 6, 52,
    -- layer=1 filter=31 channel=70
    5, 28, 55, -10, -32, 43, -26, 17, -17,
    -- layer=1 filter=31 channel=71
    -6, -2, -7, -16, 0, 8, 15, -1, 17,
    -- layer=1 filter=31 channel=72
    -4, -9, 11, -37, -11, -18, -12, -33, -41,
    -- layer=1 filter=31 channel=73
    0, 12, -7, 16, 27, 4, 21, 28, -9,
    -- layer=1 filter=31 channel=74
    -17, -6, 10, -51, -61, -20, -6, -55, -36,
    -- layer=1 filter=31 channel=75
    19, 35, 14, -64, -5, 86, 25, 20, 40,
    -- layer=1 filter=31 channel=76
    19, -40, -26, -1, -20, -74, 33, -21, -58,
    -- layer=1 filter=31 channel=77
    -4, -33, -7, 0, -15, -21, 4, -19, -1,
    -- layer=1 filter=31 channel=78
    -18, -27, 1, 9, -52, -33, 23, -27, -40,
    -- layer=1 filter=31 channel=79
    40, 42, -10, 32, 29, 13, -2, 4, 31,
    -- layer=1 filter=31 channel=80
    -1, 17, -39, 19, -18, -27, -27, -1, -11,
    -- layer=1 filter=31 channel=81
    -11, -25, -1, 11, 1, 4, -6, -1, 19,
    -- layer=1 filter=31 channel=82
    -18, -4, -8, -7, -5, 1, -9, -5, 6,
    -- layer=1 filter=31 channel=83
    12, -30, -24, 38, 37, 0, 10, -15, 9,
    -- layer=1 filter=31 channel=84
    0, -1, 16, -19, -21, -24, 12, 7, -31,
    -- layer=1 filter=31 channel=85
    -44, -33, -15, -43, -42, -35, -69, -64, -6,
    -- layer=1 filter=31 channel=86
    15, -10, -23, 22, 1, -17, 36, -4, -32,
    -- layer=1 filter=31 channel=87
    -4, -6, -27, -63, -39, -18, -34, -10, -4,
    -- layer=1 filter=31 channel=88
    -10, -8, 2, -24, -3, 10, -25, -17, 10,
    -- layer=1 filter=31 channel=89
    -33, 0, 7, -18, 3, 4, 4, -21, 0,
    -- layer=1 filter=31 channel=90
    57, -9, 0, 49, 49, 10, 39, 11, 22,
    -- layer=1 filter=31 channel=91
    -10, 7, 9, -1, -25, 5, -6, -18, -22,
    -- layer=1 filter=31 channel=92
    4, -16, -11, 0, -13, 11, 25, -33, -18,
    -- layer=1 filter=31 channel=93
    7, 2, 0, 2, 14, -14, 9, -1, -1,
    -- layer=1 filter=31 channel=94
    -35, -47, -50, -22, -75, -63, 21, -15, -37,
    -- layer=1 filter=31 channel=95
    12, 13, 0, -35, -38, 21, 39, 4, -39,
    -- layer=1 filter=31 channel=96
    -21, -28, -23, -18, -28, -20, -28, -9, -21,
    -- layer=1 filter=31 channel=97
    -4, -13, -29, 11, 0, -34, 22, 9, -3,
    -- layer=1 filter=31 channel=98
    -22, -16, -25, 13, 7, -18, -11, -2, 28,
    -- layer=1 filter=31 channel=99
    -40, -78, -32, -52, -125, -120, -8, -73, -161,
    -- layer=1 filter=31 channel=100
    13, 5, -15, 0, -27, -25, 32, -9, -30,
    -- layer=1 filter=31 channel=101
    -13, -1, 2, 11, 4, 6, 3, 0, -6,
    -- layer=1 filter=31 channel=102
    -37, -56, -25, -6, -34, -28, 22, -1, -26,
    -- layer=1 filter=31 channel=103
    35, 24, 25, 16, -6, -21, 13, 13, -14,
    -- layer=1 filter=31 channel=104
    3, 21, 14, -6, -2, 23, 12, -43, -8,
    -- layer=1 filter=31 channel=105
    -18, -36, -20, -1, -52, -52, 15, -4, -37,
    -- layer=1 filter=31 channel=106
    24, 7, -6, 10, 17, 1, 24, 14, 5,
    -- layer=1 filter=31 channel=107
    0, -1, 13, 1, 12, 12, 10, 11, 0,
    -- layer=1 filter=31 channel=108
    62, 26, 22, 39, 56, 30, 20, 34, 37,
    -- layer=1 filter=31 channel=109
    1, 2, 1, 5, 0, -3, 8, -11, 3,
    -- layer=1 filter=31 channel=110
    -28, -25, -36, -18, -20, -25, -19, -13, -39,
    -- layer=1 filter=31 channel=111
    5, 7, 11, -2, -39, 12, 22, 5, -40,
    -- layer=1 filter=31 channel=112
    10, 5, -2, 16, -24, 2, 3, -17, -25,
    -- layer=1 filter=31 channel=113
    23, 36, 31, -36, -24, 8, -18, -28, -12,
    -- layer=1 filter=31 channel=114
    25, 39, -3, 50, 35, 33, 35, 17, 22,
    -- layer=1 filter=31 channel=115
    -42, -24, -38, -27, -75, -68, -8, -46, -61,
    -- layer=1 filter=31 channel=116
    -9, 8, -7, 0, -6, -2, 9, 8, 0,
    -- layer=1 filter=31 channel=117
    -1, 26, 35, 33, 0, 46, -25, -32, 6,
    -- layer=1 filter=31 channel=118
    -2, -6, 4, -42, -37, -27, 25, -6, -19,
    -- layer=1 filter=31 channel=119
    56, -20, -7, 33, 35, -12, 40, 12, 6,
    -- layer=1 filter=31 channel=120
    -13, 7, 21, -30, -36, 0, -17, -28, 7,
    -- layer=1 filter=31 channel=121
    23, 3, -4, -27, 19, 73, 23, 36, 15,
    -- layer=1 filter=31 channel=122
    10, 4, 5, -1, 2, 9, 0, 2, 8,
    -- layer=1 filter=31 channel=123
    21, 6, 4, -14, 10, 29, 21, 0, -5,
    -- layer=1 filter=31 channel=124
    -13, -11, -13, 12, 17, 15, -10, -10, 7,
    -- layer=1 filter=31 channel=125
    -3, 15, 30, -17, -46, 9, -20, -19, -43,
    -- layer=1 filter=31 channel=126
    -12, -18, 0, 33, 38, -7, 5, 0, 57,
    -- layer=1 filter=31 channel=127
    12, 6, 8, -27, -16, 6, 22, 13, -17,
    -- layer=1 filter=32 channel=0
    -5, -22, -12, 3, -4, 12, 9, 20, 4,
    -- layer=1 filter=32 channel=1
    10, -14, 16, 27, 19, 3, 15, -2, -5,
    -- layer=1 filter=32 channel=2
    8, 11, 17, -14, -2, 2, -42, -37, -50,
    -- layer=1 filter=32 channel=3
    14, 1, 5, -3, 9, -9, -1, 6, 4,
    -- layer=1 filter=32 channel=4
    -15, 2, -13, -14, -4, -8, 3, 9, 7,
    -- layer=1 filter=32 channel=5
    37, 35, 42, 13, 26, 8, 0, 0, 13,
    -- layer=1 filter=32 channel=6
    -21, -17, 0, -36, -23, 0, -5, 21, 8,
    -- layer=1 filter=32 channel=7
    -21, 3, 10, -42, -14, -6, -5, -26, -31,
    -- layer=1 filter=32 channel=8
    42, 44, 46, 51, 62, 17, 23, 30, 20,
    -- layer=1 filter=32 channel=9
    -5, 0, -31, -24, -58, 14, -21, -18, 12,
    -- layer=1 filter=32 channel=10
    -34, -1, 16, -26, 0, -27, 12, -20, -30,
    -- layer=1 filter=32 channel=11
    -14, -17, -11, -16, -17, 0, 9, 18, 17,
    -- layer=1 filter=32 channel=12
    12, -17, -27, -48, -54, -47, -19, 20, -9,
    -- layer=1 filter=32 channel=13
    -2, 7, 2, 4, -5, 12, 5, 5, 10,
    -- layer=1 filter=32 channel=14
    0, 33, 12, -54, -12, -8, 8, -2, -34,
    -- layer=1 filter=32 channel=15
    24, 6, 19, 18, 22, -9, -8, -12, 8,
    -- layer=1 filter=32 channel=16
    49, 53, 55, 27, 40, 15, 34, 17, 13,
    -- layer=1 filter=32 channel=17
    -20, -1, -11, 28, 28, 10, 7, -1, 8,
    -- layer=1 filter=32 channel=18
    -13, -33, 1, -23, -24, -36, -21, 30, 0,
    -- layer=1 filter=32 channel=19
    46, 77, 53, 95, 94, 58, 54, 25, 49,
    -- layer=1 filter=32 channel=20
    -4, -6, -12, 11, 7, 15, 13, 4, 9,
    -- layer=1 filter=32 channel=21
    -33, -22, -6, -13, 22, -6, 19, 23, 5,
    -- layer=1 filter=32 channel=22
    -9, -24, 2, 17, 24, 32, 14, 10, -3,
    -- layer=1 filter=32 channel=23
    -1, 4, -38, -18, -34, -21, -28, -57, -1,
    -- layer=1 filter=32 channel=24
    1, 8, 17, 27, 13, 10, 9, 0, 24,
    -- layer=1 filter=32 channel=25
    -9, 29, 28, 17, 14, 22, 21, -16, 0,
    -- layer=1 filter=32 channel=26
    13, 24, 0, 12, -21, 19, -22, -10, 3,
    -- layer=1 filter=32 channel=27
    -23, -10, -20, -35, -22, -28, -9, 9, -9,
    -- layer=1 filter=32 channel=28
    -24, -10, -2, -14, 4, 0, 12, -9, -10,
    -- layer=1 filter=32 channel=29
    -32, -35, -37, -15, -33, -22, 6, -5, -7,
    -- layer=1 filter=32 channel=30
    -3, 14, 6, 20, 12, 18, 19, 64, 39,
    -- layer=1 filter=32 channel=31
    -26, -15, -13, -56, -35, -13, -19, 0, -23,
    -- layer=1 filter=32 channel=32
    18, -8, -31, -31, -73, 0, -10, 0, -9,
    -- layer=1 filter=32 channel=33
    -17, -16, -6, 9, 17, 31, 10, 4, -3,
    -- layer=1 filter=32 channel=34
    -7, -3, 23, 4, 5, 32, -19, -2, -4,
    -- layer=1 filter=32 channel=35
    32, 27, 20, 2, 20, 10, -2, 6, 21,
    -- layer=1 filter=32 channel=36
    -15, -21, -21, -4, -15, -15, 10, 11, 9,
    -- layer=1 filter=32 channel=37
    30, 49, 38, 40, 42, 8, 6, -7, 10,
    -- layer=1 filter=32 channel=38
    -19, -19, -7, -1, 2, 5, 13, 11, 7,
    -- layer=1 filter=32 channel=39
    -25, -2, -7, -9, 5, 8, -3, -3, -17,
    -- layer=1 filter=32 channel=40
    -5, 0, 14, -38, -18, -8, -11, 13, -24,
    -- layer=1 filter=32 channel=41
    -1, 20, -42, -18, -50, 39, -10, 38, 22,
    -- layer=1 filter=32 channel=42
    -27, 11, 1, 12, 21, 26, -35, -37, -47,
    -- layer=1 filter=32 channel=43
    18, 39, 24, 33, 46, -10, 4, 25, -6,
    -- layer=1 filter=32 channel=44
    0, -10, -8, -3, -35, 19, 1, -2, -13,
    -- layer=1 filter=32 channel=45
    -5, 0, 19, 15, 4, 1, -8, 10, 13,
    -- layer=1 filter=32 channel=46
    46, 58, 62, 53, 63, 17, 26, -12, -23,
    -- layer=1 filter=32 channel=47
    12, -31, -52, -27, -31, 6, -53, -9, 17,
    -- layer=1 filter=32 channel=48
    -31, -18, -32, -5, -1, 2, 7, 26, 12,
    -- layer=1 filter=32 channel=49
    -14, -5, -20, -24, -7, 5, 2, 25, 0,
    -- layer=1 filter=32 channel=50
    -15, -25, 3, -9, -19, -11, -8, -9, -3,
    -- layer=1 filter=32 channel=51
    -45, -29, -8, -14, -10, -3, 21, 14, 14,
    -- layer=1 filter=32 channel=52
    0, -3, 2, 2, -8, 3, -3, -9, -1,
    -- layer=1 filter=32 channel=53
    1, 5, 4, -2, 7, -8, 8, 17, 4,
    -- layer=1 filter=32 channel=54
    -15, 25, 20, 11, 14, 0, 30, -20, 5,
    -- layer=1 filter=32 channel=55
    2, -1, -11, -9, -6, 0, -4, -1, -9,
    -- layer=1 filter=32 channel=56
    0, -9, 0, 8, -8, 9, -10, 11, 1,
    -- layer=1 filter=32 channel=57
    -40, -4, 7, -15, 4, -19, 6, -20, -9,
    -- layer=1 filter=32 channel=58
    -23, -26, -27, -42, -57, -39, -33, -59, -10,
    -- layer=1 filter=32 channel=59
    10, 0, 11, 0, 23, 15, 22, 17, -3,
    -- layer=1 filter=32 channel=60
    -7, -7, -11, -12, -17, -6, -5, -21, -10,
    -- layer=1 filter=32 channel=61
    5, -5, -2, -4, 3, 14, 0, 0, 3,
    -- layer=1 filter=32 channel=62
    51, 68, 42, 62, 62, 31, 23, 8, 29,
    -- layer=1 filter=32 channel=63
    -23, -18, -17, -12, -16, -13, 7, 26, 27,
    -- layer=1 filter=32 channel=64
    -17, -12, -12, 6, 10, 11, 19, 19, 0,
    -- layer=1 filter=32 channel=65
    -31, -19, -5, -4, 16, -8, 30, 23, 15,
    -- layer=1 filter=32 channel=66
    -11, -6, -15, -3, 9, 9, 20, 12, 20,
    -- layer=1 filter=32 channel=67
    -41, -42, -31, -6, -10, -6, 0, 25, 3,
    -- layer=1 filter=32 channel=68
    19, -18, 2, -29, -64, 4, -16, 7, -5,
    -- layer=1 filter=32 channel=69
    36, 32, 32, 19, 2, -2, -18, -3, 7,
    -- layer=1 filter=32 channel=70
    9, 26, 27, -11, -14, 5, 0, 11, 12,
    -- layer=1 filter=32 channel=71
    -26, -7, -9, -4, 8, 0, 19, 0, 0,
    -- layer=1 filter=32 channel=72
    0, -6, -2, 32, 18, 21, 5, 43, -1,
    -- layer=1 filter=32 channel=73
    -2, -13, -14, -8, -5, 1, -5, 1, 0,
    -- layer=1 filter=32 channel=74
    2, -28, 1, -30, -75, -8, 9, 1, -17,
    -- layer=1 filter=32 channel=75
    -20, -40, -13, -6, -48, -6, -25, 15, -1,
    -- layer=1 filter=32 channel=76
    -22, -26, -35, -3, -39, 14, 11, 23, 28,
    -- layer=1 filter=32 channel=77
    -30, -42, -28, -8, -10, -5, 18, 21, 18,
    -- layer=1 filter=32 channel=78
    -17, -13, 8, -1, -14, 0, 31, 7, 13,
    -- layer=1 filter=32 channel=79
    44, 35, 40, 33, 44, 12, 12, 4, 22,
    -- layer=1 filter=32 channel=80
    12, 2, 17, 19, 0, 17, 9, 2, 6,
    -- layer=1 filter=32 channel=81
    -9, -11, -19, 0, 22, -1, 4, -4, 11,
    -- layer=1 filter=32 channel=82
    -26, -20, -14, -4, 10, 0, 22, 40, 17,
    -- layer=1 filter=32 channel=83
    20, -3, 22, 10, 3, 23, -4, 9, 17,
    -- layer=1 filter=32 channel=84
    30, 1, 1, -13, -23, 0, -17, 32, -2,
    -- layer=1 filter=32 channel=85
    6, -28, -29, -32, -49, -42, -58, -36, 17,
    -- layer=1 filter=32 channel=86
    -13, -3, 0, -11, -13, -7, 0, -3, 12,
    -- layer=1 filter=32 channel=87
    4, 29, 17, 19, 0, 25, 18, 12, 21,
    -- layer=1 filter=32 channel=88
    -11, -4, -28, -13, 3, 0, 2, 14, 0,
    -- layer=1 filter=32 channel=89
    -18, -23, -13, -10, -7, 0, 12, 34, 10,
    -- layer=1 filter=32 channel=90
    18, 9, 14, 12, -13, 22, -16, -26, 2,
    -- layer=1 filter=32 channel=91
    -28, -38, -8, -17, -14, -2, 17, 18, 2,
    -- layer=1 filter=32 channel=92
    -3, -5, 0, 3, -62, 17, -3, 3, 19,
    -- layer=1 filter=32 channel=93
    -17, -18, -20, 8, 4, 13, 22, 3, 11,
    -- layer=1 filter=32 channel=94
    -18, -21, -3, -2, -3, 1, 19, 11, 22,
    -- layer=1 filter=32 channel=95
    11, 17, 17, -17, -8, 0, 13, 33, 26,
    -- layer=1 filter=32 channel=96
    2, 0, 0, 0, -5, -7, -1, -7, -2,
    -- layer=1 filter=32 channel=97
    -17, -19, -17, 8, 0, 12, 15, 15, 12,
    -- layer=1 filter=32 channel=98
    8, 24, 12, 34, 51, 2, 16, 0, 3,
    -- layer=1 filter=32 channel=99
    -31, -11, -17, -28, -31, -64, 20, -20, -14,
    -- layer=1 filter=32 channel=100
    -18, -29, -12, -18, -24, 3, 21, 31, 21,
    -- layer=1 filter=32 channel=101
    -19, -26, -9, -8, 2, -11, 20, 29, 8,
    -- layer=1 filter=32 channel=102
    -16, -35, -11, -2, -12, 2, 18, 38, 29,
    -- layer=1 filter=32 channel=103
    -25, -21, -20, -6, -14, -6, 2, 25, 17,
    -- layer=1 filter=32 channel=104
    25, -9, -3, -29, -35, -21, -21, 0, 18,
    -- layer=1 filter=32 channel=105
    -10, -12, -13, 0, 2, -6, 25, 1, 11,
    -- layer=1 filter=32 channel=106
    1, -21, -30, -21, -28, 0, 3, 12, 13,
    -- layer=1 filter=32 channel=107
    -10, -11, -28, -3, -22, -7, -14, 0, -5,
    -- layer=1 filter=32 channel=108
    16, 9, 2, -9, -28, 16, -7, -4, 13,
    -- layer=1 filter=32 channel=109
    0, -5, 0, 8, 7, -5, 0, -2, 10,
    -- layer=1 filter=32 channel=110
    -23, -23, -3, 2, 10, -5, 17, 3, 0,
    -- layer=1 filter=32 channel=111
    17, 6, 7, 4, -2, -6, 4, 38, 28,
    -- layer=1 filter=32 channel=112
    20, 23, 49, 17, 7, 42, 11, 24, -4,
    -- layer=1 filter=32 channel=113
    -31, 25, 20, 10, 16, 41, 0, -4, -5,
    -- layer=1 filter=32 channel=114
    30, 21, 43, 12, 14, -9, -23, -7, -4,
    -- layer=1 filter=32 channel=115
    -21, -19, -14, 1, -3, -17, 0, -6, 7,
    -- layer=1 filter=32 channel=116
    -1, -3, -3, 4, -4, 8, 7, 8, -5,
    -- layer=1 filter=32 channel=117
    39, 52, 59, 38, 48, 20, 33, 17, 11,
    -- layer=1 filter=32 channel=118
    2, -1, -3, -5, -33, -10, 9, 34, 21,
    -- layer=1 filter=32 channel=119
    9, 10, -20, -13, -49, 15, -29, -6, -3,
    -- layer=1 filter=32 channel=120
    -25, -6, -3, -9, 10, 15, 13, 17, 12,
    -- layer=1 filter=32 channel=121
    -4, 5, 0, -8, 22, 29, 27, 16, 23,
    -- layer=1 filter=32 channel=122
    9, -7, -3, 1, -6, -4, 5, 8, -2,
    -- layer=1 filter=32 channel=123
    -14, -12, -12, -23, -13, 7, 5, 11, 4,
    -- layer=1 filter=32 channel=124
    -5, 6, 4, 17, 0, -6, -3, 0, 3,
    -- layer=1 filter=32 channel=125
    -3, 17, 15, -26, 0, 20, -12, 8, 2,
    -- layer=1 filter=32 channel=126
    35, 23, 29, 74, 75, 47, 36, 33, 11,
    -- layer=1 filter=32 channel=127
    10, 1, 3, -2, -3, 2, 22, 53, 14,
    -- layer=1 filter=33 channel=0
    9, 11, 15, -4, -6, -7, 4, -15, -2,
    -- layer=1 filter=33 channel=1
    -13, -4, -13, -4, 14, 0, -15, 1, -19,
    -- layer=1 filter=33 channel=2
    -37, -34, -2, -23, -38, -31, 0, -9, 6,
    -- layer=1 filter=33 channel=3
    -2, -7, 0, -7, -5, 0, -2, 1, 7,
    -- layer=1 filter=33 channel=4
    8, 8, 7, 6, 4, -7, 0, -7, -2,
    -- layer=1 filter=33 channel=5
    -24, -32, -11, 0, 24, -17, 2, -9, -16,
    -- layer=1 filter=33 channel=6
    20, 21, 10, -21, 0, 8, -17, 10, 6,
    -- layer=1 filter=33 channel=7
    14, -11, 5, 24, 1, 23, 8, -16, -6,
    -- layer=1 filter=33 channel=8
    -35, -35, -19, 4, 15, 11, 10, 16, -22,
    -- layer=1 filter=33 channel=9
    -11, 49, 7, 8, -52, 11, -24, -8, 11,
    -- layer=1 filter=33 channel=10
    0, 2, 22, 8, 0, 29, -11, 2, -3,
    -- layer=1 filter=33 channel=11
    0, -2, 8, -29, -10, -24, -10, -2, -9,
    -- layer=1 filter=33 channel=12
    19, 2, -28, 22, -8, 7, 40, 29, 23,
    -- layer=1 filter=33 channel=13
    -9, 7, 7, 9, 19, 8, -6, 13, -13,
    -- layer=1 filter=33 channel=14
    -4, -28, 11, 22, 20, 37, 23, 9, 21,
    -- layer=1 filter=33 channel=15
    -37, 3, -2, -18, 9, -24, 37, 12, 20,
    -- layer=1 filter=33 channel=16
    -12, -26, -19, 5, 34, 0, 6, 0, -23,
    -- layer=1 filter=33 channel=17
    -7, 6, 9, 9, 2, -1, 2, -9, -20,
    -- layer=1 filter=33 channel=18
    16, 29, 5, -8, -25, -22, 19, 27, 15,
    -- layer=1 filter=33 channel=19
    28, 68, 36, 79, 27, 4, 11, 47, 4,
    -- layer=1 filter=33 channel=20
    -4, 5, -1, -11, 2, 11, 1, -10, -15,
    -- layer=1 filter=33 channel=21
    -8, -32, -4, -24, -12, 8, -34, -11, -11,
    -- layer=1 filter=33 channel=22
    -8, -6, -11, -9, 18, 15, -5, -5, -8,
    -- layer=1 filter=33 channel=23
    22, 36, -11, 7, -17, 8, 21, 16, -15,
    -- layer=1 filter=33 channel=24
    -19, -18, -10, 4, -9, -34, -29, -17, -14,
    -- layer=1 filter=33 channel=25
    13, -5, 3, 10, 15, 14, 4, -8, -14,
    -- layer=1 filter=33 channel=26
    -16, 25, 13, 15, 0, -6, 2, 8, -6,
    -- layer=1 filter=33 channel=27
    21, 29, 20, -26, -30, -5, -41, -29, -39,
    -- layer=1 filter=33 channel=28
    6, -5, 19, 4, 1, 27, -28, -13, -12,
    -- layer=1 filter=33 channel=29
    6, 4, -1, -20, -29, -33, -17, -17, -22,
    -- layer=1 filter=33 channel=30
    18, 29, 34, 0, -3, 0, 20, 35, 22,
    -- layer=1 filter=33 channel=31
    34, 1, -4, 22, -2, 3, 19, 13, 3,
    -- layer=1 filter=33 channel=32
    3, 26, 2, 29, 1, 13, -6, 17, 12,
    -- layer=1 filter=33 channel=33
    21, 28, 24, 6, -1, -2, -2, 5, -14,
    -- layer=1 filter=33 channel=34
    29, 22, 10, 15, 20, 11, 18, 12, 0,
    -- layer=1 filter=33 channel=35
    -8, -6, -5, -7, -17, -20, -9, 4, 0,
    -- layer=1 filter=33 channel=36
    2, 5, 0, -27, -15, -20, -20, -21, -18,
    -- layer=1 filter=33 channel=37
    -5, -13, -24, 8, 28, -20, -19, -5, -19,
    -- layer=1 filter=33 channel=38
    0, 8, 15, -7, 8, 9, -15, -16, 1,
    -- layer=1 filter=33 channel=39
    0, 13, 0, -8, -7, -15, -13, -16, -19,
    -- layer=1 filter=33 channel=40
    11, 9, 21, -11, -21, 6, 11, 17, 0,
    -- layer=1 filter=33 channel=41
    -22, 26, -10, 38, 10, 29, -7, 19, 20,
    -- layer=1 filter=33 channel=42
    -38, -41, -27, -28, -41, -28, 6, 0, -4,
    -- layer=1 filter=33 channel=43
    -2, -23, -15, -5, 12, 0, -1, 13, -22,
    -- layer=1 filter=33 channel=44
    -10, 16, 6, 8, 2, 7, -5, 14, 5,
    -- layer=1 filter=33 channel=45
    -25, -10, -2, 8, 6, -3, -3, -11, 4,
    -- layer=1 filter=33 channel=46
    31, 19, 23, 22, 33, 3, 2, 10, 30,
    -- layer=1 filter=33 channel=47
    -4, 22, -21, 46, -15, 13, -7, 1, -20,
    -- layer=1 filter=33 channel=48
    -6, -5, 16, -20, -13, 0, -24, -12, -2,
    -- layer=1 filter=33 channel=49
    6, 15, -9, 2, -5, -3, -16, -13, -12,
    -- layer=1 filter=33 channel=50
    4, 2, -6, 2, -16, -4, 0, -16, -14,
    -- layer=1 filter=33 channel=51
    12, 2, 4, -19, -10, 8, -7, -19, 0,
    -- layer=1 filter=33 channel=52
    12, -1, 5, -8, -10, -8, 6, 27, 22,
    -- layer=1 filter=33 channel=53
    -13, 3, 1, 1, -12, -1, 0, -5, -5,
    -- layer=1 filter=33 channel=54
    22, 0, 4, 9, 34, -4, 11, -13, -23,
    -- layer=1 filter=33 channel=55
    -18, -24, -15, -15, -24, -28, -11, -18, -23,
    -- layer=1 filter=33 channel=56
    -2, -6, 3, 3, -3, 10, 7, -1, 14,
    -- layer=1 filter=33 channel=57
    11, -3, 15, 6, 12, 10, -13, -15, -5,
    -- layer=1 filter=33 channel=58
    23, 23, 14, 38, 5, 18, 17, 12, -20,
    -- layer=1 filter=33 channel=59
    -8, -11, 2, -14, 2, -9, -5, 5, -5,
    -- layer=1 filter=33 channel=60
    0, -12, 12, 0, 7, 7, 0, 1, 7,
    -- layer=1 filter=33 channel=61
    -5, 6, 4, 12, 4, 8, 2, -2, 4,
    -- layer=1 filter=33 channel=62
    -2, -13, -22, 14, 39, -9, 13, 1, -11,
    -- layer=1 filter=33 channel=63
    4, 2, 14, -11, -16, -18, -18, -17, -26,
    -- layer=1 filter=33 channel=64
    -3, 5, -7, -14, -2, -6, -3, -7, -6,
    -- layer=1 filter=33 channel=65
    7, -2, 8, -13, -17, 2, -15, -21, 10,
    -- layer=1 filter=33 channel=66
    15, 0, 11, 2, 0, -4, -4, -17, -4,
    -- layer=1 filter=33 channel=67
    7, 3, -16, -24, -42, -29, -39, -36, -20,
    -- layer=1 filter=33 channel=68
    4, 22, 10, 13, 7, 9, 3, 8, 15,
    -- layer=1 filter=33 channel=69
    -47, -37, -31, 25, 27, -19, 22, 0, 2,
    -- layer=1 filter=33 channel=70
    27, 14, 0, 1, 13, 10, -6, 13, 0,
    -- layer=1 filter=33 channel=71
    -4, -2, -5, -38, -9, -27, -32, -36, -27,
    -- layer=1 filter=33 channel=72
    11, 39, 27, 33, -11, 28, 20, 42, 15,
    -- layer=1 filter=33 channel=73
    -2, -9, 3, -1, -4, -6, -7, -5, -15,
    -- layer=1 filter=33 channel=74
    25, 22, 2, -17, -17, 13, 0, 16, 15,
    -- layer=1 filter=33 channel=75
    24, 22, -13, 12, -14, 19, 34, 14, 18,
    -- layer=1 filter=33 channel=76
    15, 33, 19, 1, -1, -12, 4, 7, 0,
    -- layer=1 filter=33 channel=77
    -5, -9, -10, -16, -21, -3, -32, -30, -2,
    -- layer=1 filter=33 channel=78
    9, -1, 4, -6, 7, 6, 2, 2, -8,
    -- layer=1 filter=33 channel=79
    -7, -19, -3, 16, 21, -20, 6, 3, -19,
    -- layer=1 filter=33 channel=80
    16, 0, 4, 4, 0, 3, 15, 13, 0,
    -- layer=1 filter=33 channel=81
    -11, 0, -17, -11, -26, -35, -24, -32, -38,
    -- layer=1 filter=33 channel=82
    -16, 0, -4, -30, -17, -5, -14, -15, -5,
    -- layer=1 filter=33 channel=83
    -22, 16, -5, 9, 12, -7, 15, 17, 3,
    -- layer=1 filter=33 channel=84
    23, 40, 32, 0, -1, 2, 14, 47, 22,
    -- layer=1 filter=33 channel=85
    -5, 22, 0, 34, -2, 5, 0, 20, -20,
    -- layer=1 filter=33 channel=86
    -10, -12, 4, -9, -7, 0, -4, -17, -28,
    -- layer=1 filter=33 channel=87
    -3, 22, -4, 78, -1, 18, -27, 51, 27,
    -- layer=1 filter=33 channel=88
    -2, 6, -11, -16, -3, 0, -20, -3, -18,
    -- layer=1 filter=33 channel=89
    0, -1, 0, -29, -24, -16, -29, -8, -20,
    -- layer=1 filter=33 channel=90
    -37, 1, 2, 12, 15, 0, 8, 20, -4,
    -- layer=1 filter=33 channel=91
    -4, 3, 9, 1, -11, 0, -5, 6, 5,
    -- layer=1 filter=33 channel=92
    -63, 31, 13, 0, -34, 24, -18, -14, 39,
    -- layer=1 filter=33 channel=93
    5, -10, -16, -22, -11, -3, -22, -18, -17,
    -- layer=1 filter=33 channel=94
    18, 1, 5, -9, -16, 0, 0, -7, -7,
    -- layer=1 filter=33 channel=95
    50, 31, 11, 6, 1, 4, 37, 49, 16,
    -- layer=1 filter=33 channel=96
    2, 17, 11, -4, 0, 6, 0, -6, -16,
    -- layer=1 filter=33 channel=97
    -1, 2, 1, 0, -7, -14, -14, -20, -7,
    -- layer=1 filter=33 channel=98
    -15, -15, -20, -2, 7, 7, 19, 20, 10,
    -- layer=1 filter=33 channel=99
    19, -4, 40, -2, 2, 23, -24, -4, 11,
    -- layer=1 filter=33 channel=100
    8, 4, 12, -19, -7, -12, -3, -11, 3,
    -- layer=1 filter=33 channel=101
    12, 8, 16, -17, -16, 3, -9, 3, -11,
    -- layer=1 filter=33 channel=102
    24, 9, 15, -5, -8, -4, 9, -15, -10,
    -- layer=1 filter=33 channel=103
    -8, 3, 1, -21, -5, -16, -2, -6, 2,
    -- layer=1 filter=33 channel=104
    3, 28, -15, 18, -8, 22, 9, 17, 27,
    -- layer=1 filter=33 channel=105
    17, -4, 16, -3, -12, -7, 0, -26, -12,
    -- layer=1 filter=33 channel=106
    4, 21, 0, 4, 3, 1, -15, -2, -4,
    -- layer=1 filter=33 channel=107
    -18, -13, -17, -29, -29, -22, -13, -10, -1,
    -- layer=1 filter=33 channel=108
    -18, 6, 0, 15, 2, -3, -5, 16, 7,
    -- layer=1 filter=33 channel=109
    -7, -2, 4, -3, -7, -6, -1, -6, 8,
    -- layer=1 filter=33 channel=110
    11, 14, 0, 4, -4, 1, 5, 0, -2,
    -- layer=1 filter=33 channel=111
    26, 26, 32, 2, -11, -6, 6, 47, 13,
    -- layer=1 filter=33 channel=112
    30, 9, -14, -6, -8, -20, 17, 19, 0,
    -- layer=1 filter=33 channel=113
    7, -9, -6, -1, 9, -5, -17, -14, -28,
    -- layer=1 filter=33 channel=114
    -33, -52, -41, -3, 20, -27, 9, 7, -6,
    -- layer=1 filter=33 channel=115
    -1, -4, 15, -3, -8, 13, -19, -31, -7,
    -- layer=1 filter=33 channel=116
    6, -5, -6, 6, 3, -2, 2, 10, -7,
    -- layer=1 filter=33 channel=117
    30, 20, 26, 22, 29, 3, 37, 47, 19,
    -- layer=1 filter=33 channel=118
    27, 39, 23, -10, -8, -2, 16, 27, 10,
    -- layer=1 filter=33 channel=119
    -6, 28, 6, 25, -1, 6, 0, 15, 8,
    -- layer=1 filter=33 channel=120
    -10, -6, 5, -17, -7, 0, -1, -31, -3,
    -- layer=1 filter=33 channel=121
    5, 0, 9, 14, -1, 0, -2, 20, 8,
    -- layer=1 filter=33 channel=122
    4, -1, 0, 0, -10, 8, -7, 0, 10,
    -- layer=1 filter=33 channel=123
    0, 4, 3, -14, -9, -8, -21, -12, -16,
    -- layer=1 filter=33 channel=124
    0, 5, -17, -1, -3, -6, -4, -5, 5,
    -- layer=1 filter=33 channel=125
    8, 17, 11, 16, 4, 14, -29, -1, -4,
    -- layer=1 filter=33 channel=126
    -24, 14, -14, 14, -4, 7, 22, 19, 1,
    -- layer=1 filter=33 channel=127
    19, 36, 12, 0, -7, 4, 32, 55, 23,
    -- layer=1 filter=34 channel=0
    -1, 12, 24, -7, 0, 19, 10, 7, 14,
    -- layer=1 filter=34 channel=1
    16, 31, 26, 40, 28, 10, 13, 15, 5,
    -- layer=1 filter=34 channel=2
    43, 47, 35, 19, 26, -11, 1, 1, -16,
    -- layer=1 filter=34 channel=3
    0, 5, 5, -7, 0, -5, 6, 7, 8,
    -- layer=1 filter=34 channel=4
    -5, 4, 10, 3, 12, 9, -5, 7, -5,
    -- layer=1 filter=34 channel=5
    11, 34, 16, 64, 26, 18, 7, 21, 23,
    -- layer=1 filter=34 channel=6
    42, 23, 9, 25, 10, 17, 31, 22, -6,
    -- layer=1 filter=34 channel=7
    17, 34, 20, 5, 17, -7, 16, 9, -21,
    -- layer=1 filter=34 channel=8
    13, 28, 22, 55, 35, 21, 18, 28, 11,
    -- layer=1 filter=34 channel=9
    11, 32, 44, -8, -35, 0, -2, -19, -6,
    -- layer=1 filter=34 channel=10
    30, 34, 6, -11, 13, 0, 7, 9, -23,
    -- layer=1 filter=34 channel=11
    -6, -3, 14, -11, 2, 11, -4, -4, -6,
    -- layer=1 filter=34 channel=12
    71, 61, 54, 7, 75, 8, -2, 14, 4,
    -- layer=1 filter=34 channel=13
    -3, -17, -23, 19, -12, -5, 13, 0, -11,
    -- layer=1 filter=34 channel=14
    17, 48, -2, -5, 29, 6, -55, -6, -6,
    -- layer=1 filter=34 channel=15
    2, -10, -24, 73, -21, 3, -29, -10, 10,
    -- layer=1 filter=34 channel=16
    0, 26, 0, 54, 40, -7, 23, 16, -3,
    -- layer=1 filter=34 channel=17
    3, 8, 33, -2, 22, 33, 15, 24, 16,
    -- layer=1 filter=34 channel=18
    7, 19, -2, 8, 12, 27, -4, -1, 9,
    -- layer=1 filter=34 channel=19
    27, -9, -1, 3, 0, -15, -8, -37, -35,
    -- layer=1 filter=34 channel=20
    9, 2, 10, 10, 19, 0, 10, 11, 14,
    -- layer=1 filter=34 channel=21
    0, -9, -20, 26, -15, -10, -6, 20, -9,
    -- layer=1 filter=34 channel=22
    10, 22, 12, 25, 15, 2, 19, 11, 13,
    -- layer=1 filter=34 channel=23
    -19, -43, -49, -50, -22, -47, -40, -85, -28,
    -- layer=1 filter=34 channel=24
    -34, -44, -50, -49, -41, -55, -28, -35, -25,
    -- layer=1 filter=34 channel=25
    28, 31, 17, 24, 28, 2, 42, 19, 5,
    -- layer=1 filter=34 channel=26
    -31, -63, -40, -21, -59, -20, -34, -27, 6,
    -- layer=1 filter=34 channel=27
    21, 11, -14, 4, 13, 3, 0, -5, -22,
    -- layer=1 filter=34 channel=28
    3, 41, 8, 9, 19, 6, 0, 13, -21,
    -- layer=1 filter=34 channel=29
    6, -1, -9, 4, -2, -10, 9, -3, -18,
    -- layer=1 filter=34 channel=30
    22, 10, -10, -9, 0, 28, -27, -45, -28,
    -- layer=1 filter=34 channel=31
    24, 31, 7, 3, 9, 0, -4, -11, 1,
    -- layer=1 filter=34 channel=32
    -50, -91, -72, -75, -152, -77, -66, -100, -29,
    -- layer=1 filter=34 channel=33
    -13, -4, -24, -7, -8, 2, -13, -6, -21,
    -- layer=1 filter=34 channel=34
    28, 13, 10, 11, -7, 0, -5, -12, -5,
    -- layer=1 filter=34 channel=35
    -11, -14, -14, -11, -6, -4, -2, 0, -15,
    -- layer=1 filter=34 channel=36
    -3, 6, 22, 1, 0, 20, 0, -1, 12,
    -- layer=1 filter=34 channel=37
    35, 34, 7, 39, 39, -12, 22, 34, 17,
    -- layer=1 filter=34 channel=38
    4, -12, -8, 2, 5, 4, 18, 1, -4,
    -- layer=1 filter=34 channel=39
    4, 2, 5, 11, 17, 8, 0, -10, -2,
    -- layer=1 filter=34 channel=40
    24, 21, -12, 27, 8, 25, 11, 2, 8,
    -- layer=1 filter=34 channel=41
    5, -37, -5, -7, -58, -8, -32, -69, -40,
    -- layer=1 filter=34 channel=42
    52, 24, 29, 18, 43, 1, 30, -4, -1,
    -- layer=1 filter=34 channel=43
    0, 23, 16, 56, 29, 15, 26, 28, 17,
    -- layer=1 filter=34 channel=44
    -62, -117, -55, -56, -106, -50, -63, -41, -17,
    -- layer=1 filter=34 channel=45
    -16, -1, -7, 20, 3, -9, -6, 15, 23,
    -- layer=1 filter=34 channel=46
    44, 4, 20, 20, 34, -4, 30, -21, -8,
    -- layer=1 filter=34 channel=47
    -4, -41, -36, -24, -42, -57, -1, -73, -39,
    -- layer=1 filter=34 channel=48
    13, -5, -10, 10, -3, -4, 1, 1, 10,
    -- layer=1 filter=34 channel=49
    2, -8, -15, 0, -12, -21, 11, 0, -8,
    -- layer=1 filter=34 channel=50
    2, 3, -4, 0, 0, -14, 21, 17, 7,
    -- layer=1 filter=34 channel=51
    8, -3, -13, 5, 7, -11, 26, 16, -6,
    -- layer=1 filter=34 channel=52
    7, -16, -39, 18, 12, -5, -2, -16, -19,
    -- layer=1 filter=34 channel=53
    7, 4, 16, 19, 8, 19, 17, 8, 19,
    -- layer=1 filter=34 channel=54
    30, -1, 15, -11, 29, -17, 38, 22, 3,
    -- layer=1 filter=34 channel=55
    -10, -25, -12, 3, -17, -7, -15, -30, -29,
    -- layer=1 filter=34 channel=56
    -8, 0, 7, 1, 10, 4, -7, 8, -8,
    -- layer=1 filter=34 channel=57
    30, 36, 11, 7, 25, 6, 29, 31, 0,
    -- layer=1 filter=34 channel=58
    -10, -21, -79, -41, -32, -108, -2, -41, -65,
    -- layer=1 filter=34 channel=59
    -2, -9, 11, 15, 0, 0, -5, 0, 0,
    -- layer=1 filter=34 channel=60
    -11, -11, 5, 16, 8, 18, -1, -1, 7,
    -- layer=1 filter=34 channel=61
    6, 9, 3, 0, -2, 1, 9, 0, 0,
    -- layer=1 filter=34 channel=62
    16, 31, 18, 31, 33, -1, 14, 9, 2,
    -- layer=1 filter=34 channel=63
    1, 3, 2, 6, -3, 23, -12, 3, 14,
    -- layer=1 filter=34 channel=64
    6, 0, 20, 12, 21, 6, 10, 19, 3,
    -- layer=1 filter=34 channel=65
    3, 6, 0, 0, 11, -9, 2, 12, 13,
    -- layer=1 filter=34 channel=66
    -1, 6, 11, -1, -2, 11, 4, -1, -1,
    -- layer=1 filter=34 channel=67
    -14, -14, -33, 9, -23, -30, 1, 1, -14,
    -- layer=1 filter=34 channel=68
    -94, -139, -71, -112, -165, -40, -99, -62, -21,
    -- layer=1 filter=34 channel=69
    0, 5, -36, 27, -18, -19, -4, -8, -20,
    -- layer=1 filter=34 channel=70
    34, 15, 4, 12, 11, 5, 34, 9, -6,
    -- layer=1 filter=34 channel=71
    -12, -20, -31, -10, -9, -35, -7, 2, -33,
    -- layer=1 filter=34 channel=72
    26, -9, 36, -13, -20, 23, -12, -64, -6,
    -- layer=1 filter=34 channel=73
    -2, -5, -10, 8, 6, 6, -3, -1, -7,
    -- layer=1 filter=34 channel=74
    -22, -18, -15, -16, -20, 29, -10, -1, 5,
    -- layer=1 filter=34 channel=75
    62, 57, 15, 12, 55, 7, -20, -20, -5,
    -- layer=1 filter=34 channel=76
    -13, -26, 12, -20, -5, 23, -12, 7, -3,
    -- layer=1 filter=34 channel=77
    0, -5, -2, -9, -17, -12, -6, 9, -4,
    -- layer=1 filter=34 channel=78
    -19, 11, 11, -5, 7, 5, -4, 19, 0,
    -- layer=1 filter=34 channel=79
    7, 27, 4, 39, 33, -14, 28, 2, -8,
    -- layer=1 filter=34 channel=80
    -7, 8, 2, -5, 5, 0, -7, 4, 5,
    -- layer=1 filter=34 channel=81
    -5, -23, -31, 0, -17, -14, -1, -15, -26,
    -- layer=1 filter=34 channel=82
    1, -23, -11, 1, -15, -12, 13, 14, -5,
    -- layer=1 filter=34 channel=83
    -9, -6, 2, 40, -1, 1, -22, 11, -11,
    -- layer=1 filter=34 channel=84
    -11, -25, -13, -34, -34, 4, -42, -24, -3,
    -- layer=1 filter=34 channel=85
    41, -30, -31, -12, -23, -41, 5, -17, -32,
    -- layer=1 filter=34 channel=86
    -13, 5, 23, -7, 16, 10, -4, 1, 10,
    -- layer=1 filter=34 channel=87
    31, 15, 44, 1, -40, -28, 27, -53, -18,
    -- layer=1 filter=34 channel=88
    2, -9, 10, 12, -7, 9, 20, 0, 18,
    -- layer=1 filter=34 channel=89
    -1, -16, -26, -10, -15, -6, 3, -7, -11,
    -- layer=1 filter=34 channel=90
    -65, -96, -72, -55, -101, -61, -82, -64, -37,
    -- layer=1 filter=34 channel=91
    8, 6, 12, 24, 20, 6, 21, 3, 16,
    -- layer=1 filter=34 channel=92
    -2, -19, 1, 21, -23, -51, 3, -32, -52,
    -- layer=1 filter=34 channel=93
    -4, -7, -12, -14, -13, -14, 4, -3, -8,
    -- layer=1 filter=34 channel=94
    -10, 27, 35, 5, 16, 37, 19, 23, 18,
    -- layer=1 filter=34 channel=95
    -4, 7, -27, -33, -18, 2, -41, -35, -16,
    -- layer=1 filter=34 channel=96
    21, -1, 9, 4, 5, 0, 0, 1, -5,
    -- layer=1 filter=34 channel=97
    -11, -2, 26, 5, 1, 3, 8, 0, 16,
    -- layer=1 filter=34 channel=98
    14, 33, 28, 34, 23, 1, 25, 16, -5,
    -- layer=1 filter=34 channel=99
    -84, -32, -24, -103, -71, 7, -85, -10, -42,
    -- layer=1 filter=34 channel=100
    10, -2, 16, 4, -8, -6, -11, -14, -13,
    -- layer=1 filter=34 channel=101
    -13, 1, -15, 16, 11, 2, -1, 15, 7,
    -- layer=1 filter=34 channel=102
    8, 26, 28, 23, 34, 46, 18, 38, 33,
    -- layer=1 filter=34 channel=103
    11, 19, 3, -2, -1, -5, -21, -23, -10,
    -- layer=1 filter=34 channel=104
    17, 0, -6, -22, 6, -21, -15, -34, -6,
    -- layer=1 filter=34 channel=105
    5, 7, 21, -6, 8, 19, -9, 12, 0,
    -- layer=1 filter=34 channel=106
    -22, -32, -25, -11, -28, -10, -11, 4, -5,
    -- layer=1 filter=34 channel=107
    7, 7, 9, 19, 15, 1, 2, 4, 6,
    -- layer=1 filter=34 channel=108
    -71, -143, -102, -72, -133, -72, -87, -72, -40,
    -- layer=1 filter=34 channel=109
    0, 5, 5, 0, -6, 4, 7, -3, 9,
    -- layer=1 filter=34 channel=110
    -2, 7, 14, -7, 6, 4, -5, 10, 9,
    -- layer=1 filter=34 channel=111
    25, 23, 10, 1, 19, 24, -20, -23, -8,
    -- layer=1 filter=34 channel=112
    4, 3, -16, 20, 2, -11, -6, 5, -1,
    -- layer=1 filter=34 channel=113
    21, 11, 18, 33, -7, 10, 25, -3, -4,
    -- layer=1 filter=34 channel=114
    -3, 7, -20, 56, 11, 8, -13, 12, 11,
    -- layer=1 filter=34 channel=115
    -1, 34, 32, -6, 27, 26, 8, 16, 9,
    -- layer=1 filter=34 channel=116
    4, -9, 2, 2, -3, 9, -3, -5, 1,
    -- layer=1 filter=34 channel=117
    -2, 40, 3, 13, -9, -28, -29, -27, -32,
    -- layer=1 filter=34 channel=118
    -4, -13, -5, -35, -24, 14, -38, -29, -24,
    -- layer=1 filter=34 channel=119
    -60, -119, -82, -85, -161, -88, -75, -106, -41,
    -- layer=1 filter=34 channel=120
    15, 0, -11, 21, 1, -21, 28, 12, 9,
    -- layer=1 filter=34 channel=121
    33, 12, 3, -14, 5, -8, -40, -46, -30,
    -- layer=1 filter=34 channel=122
    -2, 8, -7, -10, -2, -8, 2, 4, 5,
    -- layer=1 filter=34 channel=123
    28, -7, -15, -3, 4, -9, -28, -29, -25,
    -- layer=1 filter=34 channel=124
    -5, -16, -4, 2, 10, -9, -11, 0, 0,
    -- layer=1 filter=34 channel=125
    42, 19, 2, 12, -7, -14, 35, 1, -1,
    -- layer=1 filter=34 channel=126
    0, 15, 29, 36, 5, -4, -4, 10, -3,
    -- layer=1 filter=34 channel=127
    1, 3, -5, -28, -4, 6, -13, -18, 0,
    -- layer=1 filter=35 channel=0
    -4, -8, -15, -14, -13, -13, 9, 1, 6,
    -- layer=1 filter=35 channel=1
    -27, -24, -31, -4, 14, 5, 34, 0, 14,
    -- layer=1 filter=35 channel=2
    4, 30, 11, 5, 22, 22, 2, 3, 10,
    -- layer=1 filter=35 channel=3
    -3, 1, 1, 2, 4, 5, -10, 5, 4,
    -- layer=1 filter=35 channel=4
    -8, -2, -6, -7, -6, -5, 9, 3, 5,
    -- layer=1 filter=35 channel=5
    -12, 6, -13, 7, 21, 22, 35, 17, 17,
    -- layer=1 filter=35 channel=6
    11, 18, 42, 10, -32, -37, 13, 11, 4,
    -- layer=1 filter=35 channel=7
    -120, -83, -9, -68, -120, -41, -77, -70, 15,
    -- layer=1 filter=35 channel=8
    -21, 6, -17, 24, 19, 14, 31, 24, 37,
    -- layer=1 filter=35 channel=9
    14, -4, 7, -19, 17, -19, 34, 14, 31,
    -- layer=1 filter=35 channel=10
    -111, -88, 3, -66, -97, -35, -67, -54, 27,
    -- layer=1 filter=35 channel=11
    8, 6, 8, 28, 20, 27, 13, 20, 9,
    -- layer=1 filter=35 channel=12
    48, 24, 47, 48, 24, -9, 37, 46, 41,
    -- layer=1 filter=35 channel=13
    -23, -28, -37, -35, -36, -22, -5, -29, -23,
    -- layer=1 filter=35 channel=14
    -51, -17, 35, -42, -61, -41, -46, -26, 31,
    -- layer=1 filter=35 channel=15
    -9, -4, 5, 10, 28, 36, 16, -14, -32,
    -- layer=1 filter=35 channel=16
    -20, -8, -20, 15, 25, 21, 48, 49, 48,
    -- layer=1 filter=35 channel=17
    -23, -6, -8, -4, 0, -13, 23, 9, 6,
    -- layer=1 filter=35 channel=18
    -18, 0, 0, -10, -6, -23, -19, -11, 30,
    -- layer=1 filter=35 channel=19
    -9, -11, 13, -13, -20, -13, 14, 18, 20,
    -- layer=1 filter=35 channel=20
    -40, -24, -20, -24, -15, -33, -12, -7, -14,
    -- layer=1 filter=35 channel=21
    -27, -27, -33, -27, -19, 2, -1, -14, -12,
    -- layer=1 filter=35 channel=22
    -57, -39, -56, 4, -8, -14, 7, -16, -4,
    -- layer=1 filter=35 channel=23
    -21, -10, -7, -34, -23, 7, 3, -2, 11,
    -- layer=1 filter=35 channel=24
    6, -30, -27, -11, -2, 11, 12, -3, 14,
    -- layer=1 filter=35 channel=25
    -95, -73, -22, -20, -17, -5, -7, 4, 23,
    -- layer=1 filter=35 channel=26
    -7, -47, -62, 7, -8, -30, 22, 9, 36,
    -- layer=1 filter=35 channel=27
    -3, 3, -19, 8, 10, -11, -31, -20, -26,
    -- layer=1 filter=35 channel=28
    -116, -100, -37, -38, -78, -31, -23, -39, 10,
    -- layer=1 filter=35 channel=29
    -57, -30, -39, -52, -22, -19, -44, -35, -34,
    -- layer=1 filter=35 channel=30
    -24, -9, 5, -67, -60, -69, -48, -41, 6,
    -- layer=1 filter=35 channel=31
    -4, 16, 38, -13, -8, -14, -8, -8, 10,
    -- layer=1 filter=35 channel=32
    -9, -73, -56, -10, -63, -50, -4, -30, 34,
    -- layer=1 filter=35 channel=33
    -2, 16, -3, 2, 9, 2, 0, 5, -1,
    -- layer=1 filter=35 channel=34
    18, 8, 32, 4, -1, -9, -5, 9, -2,
    -- layer=1 filter=35 channel=35
    8, -1, -7, -5, -1, -1, 1, 7, 9,
    -- layer=1 filter=35 channel=36
    22, 16, 2, 34, 32, 14, 26, 34, 17,
    -- layer=1 filter=35 channel=37
    -9, 3, -15, 23, 37, 7, 27, 26, 19,
    -- layer=1 filter=35 channel=38
    -18, -24, 0, -25, -31, -26, -10, -25, -21,
    -- layer=1 filter=35 channel=39
    2, 0, -8, 26, 21, 13, 9, 10, -2,
    -- layer=1 filter=35 channel=40
    -32, -24, 0, -24, -52, -57, -1, 12, 3,
    -- layer=1 filter=35 channel=41
    12, -26, -34, 2, -9, -16, -12, 0, 53,
    -- layer=1 filter=35 channel=42
    13, 25, 14, -13, 0, 9, 1, 2, -1,
    -- layer=1 filter=35 channel=43
    -48, -34, -29, 27, 24, 33, 37, 19, 45,
    -- layer=1 filter=35 channel=44
    -41, -110, -74, -27, -53, -32, -2, -16, 40,
    -- layer=1 filter=35 channel=45
    -15, -37, -36, -5, 4, 12, 26, -3, -16,
    -- layer=1 filter=35 channel=46
    0, 27, 52, -25, 20, 18, 23, 39, 40,
    -- layer=1 filter=35 channel=47
    3, -12, -3, -20, -44, -15, -7, -24, 4,
    -- layer=1 filter=35 channel=48
    -33, -33, -25, -14, -13, -14, -19, -24, -18,
    -- layer=1 filter=35 channel=49
    6, -2, 12, 0, -1, -11, -12, -2, -8,
    -- layer=1 filter=35 channel=50
    3, -15, -27, -7, -13, -17, -28, -12, -3,
    -- layer=1 filter=35 channel=51
    -45, -19, 2, -25, -34, -35, -15, -37, 26,
    -- layer=1 filter=35 channel=52
    -20, -33, -15, 16, 1, 12, 13, -3, 4,
    -- layer=1 filter=35 channel=53
    10, 13, 10, 9, -2, 4, 4, 5, 9,
    -- layer=1 filter=35 channel=54
    -35, -37, -8, -9, -1, 13, -25, 21, 48,
    -- layer=1 filter=35 channel=55
    18, 27, 0, 25, 31, 25, 21, 29, 20,
    -- layer=1 filter=35 channel=56
    -2, -3, 2, -10, 3, 6, -4, -2, -9,
    -- layer=1 filter=35 channel=57
    -74, -78, -11, -47, -102, -35, -60, -62, 11,
    -- layer=1 filter=35 channel=58
    -113, -73, -19, -75, -114, -21, -37, -40, 21,
    -- layer=1 filter=35 channel=59
    -11, -1, -14, 11, -2, 3, -10, -11, -1,
    -- layer=1 filter=35 channel=60
    0, -11, -1, -13, -15, -6, -21, -7, -2,
    -- layer=1 filter=35 channel=61
    -3, 5, -4, 11, 6, -9, -3, 3, -3,
    -- layer=1 filter=35 channel=62
    -31, -22, -25, 0, 21, 14, 45, 37, 36,
    -- layer=1 filter=35 channel=63
    7, 7, 0, 19, 11, 6, 10, 21, 15,
    -- layer=1 filter=35 channel=64
    5, -12, -3, 3, -6, 10, 4, -5, 13,
    -- layer=1 filter=35 channel=65
    -29, -30, -34, -19, -19, -15, -5, -12, -16,
    -- layer=1 filter=35 channel=66
    4, -9, 8, 2, 0, -3, 15, 11, 3,
    -- layer=1 filter=35 channel=67
    -20, -10, -11, 25, -1, 24, -4, 4, 44,
    -- layer=1 filter=35 channel=68
    -60, -108, -95, -50, -94, -76, -4, -21, 29,
    -- layer=1 filter=35 channel=69
    -9, -3, -27, 29, 33, 36, 56, 32, 16,
    -- layer=1 filter=35 channel=70
    46, 65, 79, 11, -13, 0, 13, -10, 15,
    -- layer=1 filter=35 channel=71
    -12, 9, 7, -3, 5, 25, 7, 26, 21,
    -- layer=1 filter=35 channel=72
    -12, 4, 3, -32, -31, -41, -17, 0, 21,
    -- layer=1 filter=35 channel=73
    10, -2, -1, 9, -2, 5, 2, 11, 5,
    -- layer=1 filter=35 channel=74
    -27, -30, -30, -62, -61, -43, -48, 6, 25,
    -- layer=1 filter=35 channel=75
    -19, -5, 36, -51, -69, -52, -21, 19, 48,
    -- layer=1 filter=35 channel=76
    -14, -33, -18, -27, -15, -22, -13, 5, 12,
    -- layer=1 filter=35 channel=77
    -17, -16, -15, -15, -9, 2, -6, -29, -9,
    -- layer=1 filter=35 channel=78
    6, -4, -9, 0, -12, -16, -12, 7, -4,
    -- layer=1 filter=35 channel=79
    -21, -18, -21, 28, 20, 30, 48, 29, 42,
    -- layer=1 filter=35 channel=80
    1, 2, -9, 6, 5, 5, 10, -5, -10,
    -- layer=1 filter=35 channel=81
    -8, -18, -23, 9, 1, 12, 11, -1, 7,
    -- layer=1 filter=35 channel=82
    -36, -28, -26, -49, -42, -23, -12, -42, -12,
    -- layer=1 filter=35 channel=83
    -3, -27, -8, 2, 10, -20, 34, -14, 0,
    -- layer=1 filter=35 channel=84
    -48, -47, -20, -30, -49, -54, -41, 11, 51,
    -- layer=1 filter=35 channel=85
    -24, -44, -9, -46, -62, -12, -1, -37, 5,
    -- layer=1 filter=35 channel=86
    11, 18, 17, 8, 22, 22, 17, 24, 1,
    -- layer=1 filter=35 channel=87
    14, 20, 36, -36, 21, -32, 38, 48, 38,
    -- layer=1 filter=35 channel=88
    1, 2, 20, 3, 16, -1, 10, -11, 15,
    -- layer=1 filter=35 channel=89
    -31, -17, -14, -20, -29, -23, -13, -4, -4,
    -- layer=1 filter=35 channel=90
    -54, -104, -110, -19, -31, -26, 23, -27, 1,
    -- layer=1 filter=35 channel=91
    -29, -11, 0, -30, -42, -47, -10, -19, -21,
    -- layer=1 filter=35 channel=92
    22, -16, -15, -23, -3, -27, 1, -9, -5,
    -- layer=1 filter=35 channel=93
    -19, -18, -13, -14, -10, -3, 9, -14, -7,
    -- layer=1 filter=35 channel=94
    -7, -11, -5, 0, -13, -13, -8, 11, 0,
    -- layer=1 filter=35 channel=95
    -45, -33, -2, -54, -78, -65, -59, -6, 38,
    -- layer=1 filter=35 channel=96
    12, 22, 11, 22, 11, 2, 6, 25, 7,
    -- layer=1 filter=35 channel=97
    -8, -10, -15, 5, -6, 1, 14, -1, -8,
    -- layer=1 filter=35 channel=98
    -74, -46, -53, 28, 1, 1, 19, -7, 27,
    -- layer=1 filter=35 channel=99
    -112, -137, -63, -94, -100, -68, -30, -75, -54,
    -- layer=1 filter=35 channel=100
    25, 27, 6, 8, 12, 1, -12, 12, 1,
    -- layer=1 filter=35 channel=101
    -34, -24, 0, -51, -49, -42, -43, -43, -36,
    -- layer=1 filter=35 channel=102
    -12, -12, -23, -25, -11, -12, -7, -17, -11,
    -- layer=1 filter=35 channel=103
    2, 7, -2, -1, 9, -3, -17, -11, -5,
    -- layer=1 filter=35 channel=104
    12, 5, 10, -20, -46, 0, 3, -6, 22,
    -- layer=1 filter=35 channel=105
    -10, -18, -5, -10, 7, -10, 2, 3, 0,
    -- layer=1 filter=35 channel=106
    -13, -24, -3, -30, -56, -63, -26, -30, -7,
    -- layer=1 filter=35 channel=107
    1, 6, 8, 13, 9, 16, 11, -7, 11,
    -- layer=1 filter=35 channel=108
    -16, -92, -87, -17, -54, -26, 5, -5, 15,
    -- layer=1 filter=35 channel=109
    0, -2, -6, -4, -4, 11, 11, 1, -7,
    -- layer=1 filter=35 channel=110
    -8, -5, 1, -5, -6, 1, 6, 1, 11,
    -- layer=1 filter=35 channel=111
    -22, -19, -15, -20, -30, -46, -36, -3, 38,
    -- layer=1 filter=35 channel=112
    -26, -42, -19, -16, -29, -22, -33, -9, 31,
    -- layer=1 filter=35 channel=113
    15, 21, 26, 6, 8, 8, 0, 0, 9,
    -- layer=1 filter=35 channel=114
    -6, 17, -21, 28, 43, 35, 62, 53, 25,
    -- layer=1 filter=35 channel=115
    -4, 1, 4, -1, 5, -2, -3, 7, 8,
    -- layer=1 filter=35 channel=116
    7, 1, -11, -7, 0, 7, -11, 0, -2,
    -- layer=1 filter=35 channel=117
    -41, -47, 4, 43, 0, -28, 1, 17, 57,
    -- layer=1 filter=35 channel=118
    -8, -29, -4, -56, -55, -55, -25, -15, 9,
    -- layer=1 filter=35 channel=119
    -23, -76, -83, -37, -71, -55, -5, -30, -1,
    -- layer=1 filter=35 channel=120
    -46, -27, -23, -21, -15, -17, -29, -24, -5,
    -- layer=1 filter=35 channel=121
    20, 15, 9, -25, -1, -3, -13, 3, -1,
    -- layer=1 filter=35 channel=122
    -6, 2, 10, -6, -10, 8, 10, -7, -2,
    -- layer=1 filter=35 channel=123
    22, 27, 21, 7, 14, 15, -13, 12, -2,
    -- layer=1 filter=35 channel=124
    1, 7, 9, 12, 14, 2, 13, 14, 16,
    -- layer=1 filter=35 channel=125
    53, 54, 65, 24, 19, 13, 11, -4, 12,
    -- layer=1 filter=35 channel=126
    -41, -35, -20, -4, -18, -24, 29, -6, 9,
    -- layer=1 filter=35 channel=127
    -22, -19, 4, -55, -41, -50, -38, -5, 34,
    -- layer=1 filter=36 channel=0
    4, -3, 0, 1, 1, 3, -4, -1, -1,
    -- layer=1 filter=36 channel=1
    -31, 10, -11, 13, -2, -16, 9, -8, 31,
    -- layer=1 filter=36 channel=2
    -41, -22, -17, -34, -15, -14, -39, -24, -52,
    -- layer=1 filter=36 channel=3
    -4, -4, -17, -3, 4, -3, 0, -3, -15,
    -- layer=1 filter=36 channel=4
    3, -1, 3, 2, -8, -9, 5, 8, 3,
    -- layer=1 filter=36 channel=5
    -30, -8, -32, 7, -23, -23, -8, -22, 16,
    -- layer=1 filter=36 channel=6
    -6, -2, -5, -12, -5, -1, -16, -3, -7,
    -- layer=1 filter=36 channel=7
    5, 16, 29, 10, -2, 47, 23, -9, 18,
    -- layer=1 filter=36 channel=8
    -22, -6, -26, 0, -25, -14, -11, -16, 40,
    -- layer=1 filter=36 channel=9
    2, -46, 19, -15, -15, -19, 21, -9, -10,
    -- layer=1 filter=36 channel=10
    2, -2, 24, 17, -14, 18, -4, -12, 13,
    -- layer=1 filter=36 channel=11
    -9, -20, -22, -3, 15, -9, -4, 5, 1,
    -- layer=1 filter=36 channel=12
    -36, -58, -28, -12, -32, -58, -28, -85, -25,
    -- layer=1 filter=36 channel=13
    10, -19, -4, -10, 9, 15, 11, 10, 13,
    -- layer=1 filter=36 channel=14
    -17, -11, -17, -9, -50, 28, 3, -44, 17,
    -- layer=1 filter=36 channel=15
    2, -33, 0, 2, -16, -1, -7, -21, 23,
    -- layer=1 filter=36 channel=16
    -16, 0, -8, 9, -12, 1, -2, 1, 32,
    -- layer=1 filter=36 channel=17
    -14, 0, -12, -5, -2, 8, -7, -5, -3,
    -- layer=1 filter=36 channel=18
    -41, -29, -54, 3, -22, -14, 4, -14, 5,
    -- layer=1 filter=36 channel=19
    11, -54, 0, 16, -13, 30, 25, 44, 27,
    -- layer=1 filter=36 channel=20
    4, 2, -9, 0, 9, 9, 6, 11, 12,
    -- layer=1 filter=36 channel=21
    -1, 1, -2, 4, -11, -12, 3, -17, 24,
    -- layer=1 filter=36 channel=22
    -4, -7, 0, 4, -8, 0, -1, 4, 16,
    -- layer=1 filter=36 channel=23
    13, 22, 67, 29, 25, 28, 23, 43, 1,
    -- layer=1 filter=36 channel=24
    15, -24, -13, -11, -6, 1, -6, 12, -3,
    -- layer=1 filter=36 channel=25
    -1, 16, 10, 20, 4, 16, 16, 6, 22,
    -- layer=1 filter=36 channel=26
    5, -29, 13, -18, 6, 27, 5, 0, 6,
    -- layer=1 filter=36 channel=27
    -46, -35, -31, -48, -27, -39, -74, -31, -38,
    -- layer=1 filter=36 channel=28
    3, 13, 13, 18, -3, 12, 0, -35, 28,
    -- layer=1 filter=36 channel=29
    6, 0, 6, 3, -6, -10, -11, -7, -11,
    -- layer=1 filter=36 channel=30
    -42, -50, -40, -12, -25, -9, 0, 7, 5,
    -- layer=1 filter=36 channel=31
    -38, -17, -19, -17, -29, -36, -22, -12, -10,
    -- layer=1 filter=36 channel=32
    8, -6, 40, 10, 21, 25, 16, -11, 5,
    -- layer=1 filter=36 channel=33
    0, 0, -11, -3, 7, 1, 12, 18, 8,
    -- layer=1 filter=36 channel=34
    0, 6, 30, -17, 5, 33, 4, 15, 36,
    -- layer=1 filter=36 channel=35
    6, 17, 11, 17, 3, 3, 4, 4, 14,
    -- layer=1 filter=36 channel=36
    -7, -22, -15, -1, -11, 0, -11, -9, -15,
    -- layer=1 filter=36 channel=37
    -23, -19, -2, 1, -24, -19, -14, 2, 12,
    -- layer=1 filter=36 channel=38
    -4, -5, -6, 0, -8, -3, 9, 12, 3,
    -- layer=1 filter=36 channel=39
    -4, -3, 6, 3, -6, 6, -9, 3, -7,
    -- layer=1 filter=36 channel=40
    -18, -21, -19, -8, 2, -5, -13, 4, 4,
    -- layer=1 filter=36 channel=41
    25, -13, 53, -10, 6, 19, 1, 0, -6,
    -- layer=1 filter=36 channel=42
    -37, -1, -3, -16, -27, -13, -39, -28, -48,
    -- layer=1 filter=36 channel=43
    -18, -5, 5, 24, -19, 9, 5, -8, 26,
    -- layer=1 filter=36 channel=44
    9, -10, 31, -2, 5, 13, 18, -3, 19,
    -- layer=1 filter=36 channel=45
    -4, -2, 2, 6, 9, 3, 8, 9, 23,
    -- layer=1 filter=36 channel=46
    -15, -47, -19, 11, -11, -10, 9, 21, 27,
    -- layer=1 filter=36 channel=47
    12, 4, 65, -2, 9, -6, 0, 35, -12,
    -- layer=1 filter=36 channel=48
    -3, 5, 5, -1, -8, -3, 7, -1, 7,
    -- layer=1 filter=36 channel=49
    -12, -1, 10, -1, 2, 12, -4, 8, 17,
    -- layer=1 filter=36 channel=50
    -14, -9, -15, -11, -12, -2, -10, 1, -12,
    -- layer=1 filter=36 channel=51
    8, 7, -12, 12, -7, 0, 8, -16, 13,
    -- layer=1 filter=36 channel=52
    19, 15, -1, -1, -3, 2, 14, 4, 9,
    -- layer=1 filter=36 channel=53
    6, 8, 9, -11, -2, 12, -6, -7, 2,
    -- layer=1 filter=36 channel=54
    12, 12, 32, 23, -16, 24, 3, 5, 35,
    -- layer=1 filter=36 channel=55
    -6, -6, 3, -16, -13, -11, -32, -5, -21,
    -- layer=1 filter=36 channel=56
    5, 15, 12, 4, 0, 7, 0, -5, 9,
    -- layer=1 filter=36 channel=57
    -4, -1, 7, 2, -18, 14, 7, -20, 3,
    -- layer=1 filter=36 channel=58
    28, 57, 64, 44, 23, 46, -1, 50, 7,
    -- layer=1 filter=36 channel=59
    5, -4, 16, 6, 7, 16, -4, 13, 13,
    -- layer=1 filter=36 channel=60
    16, 16, 0, 3, -4, 4, -3, 0, 4,
    -- layer=1 filter=36 channel=61
    11, -7, 0, -17, -2, -9, -2, -6, -6,
    -- layer=1 filter=36 channel=62
    -8, -13, -16, 12, -37, 7, -7, 0, 32,
    -- layer=1 filter=36 channel=63
    -15, -19, -17, 3, 2, -18, 4, -1, -9,
    -- layer=1 filter=36 channel=64
    0, -3, -1, -12, 5, -1, 0, -4, 3,
    -- layer=1 filter=36 channel=65
    7, 3, -6, 3, -2, -10, 10, -2, -2,
    -- layer=1 filter=36 channel=66
    6, -11, -5, -9, 0, 8, -5, -13, 6,
    -- layer=1 filter=36 channel=67
    8, 14, 13, 0, -5, 9, -26, -22, 3,
    -- layer=1 filter=36 channel=68
    31, -5, 25, -5, 18, 17, 29, 4, 24,
    -- layer=1 filter=36 channel=69
    10, -3, -10, -6, -28, 6, 2, -5, 11,
    -- layer=1 filter=36 channel=70
    -22, -43, 0, -21, -17, -14, -44, -22, -18,
    -- layer=1 filter=36 channel=71
    3, 5, -17, 6, -11, 1, -9, -4, 8,
    -- layer=1 filter=36 channel=72
    -28, -52, -40, -24, -43, -27, 24, 0, -5,
    -- layer=1 filter=36 channel=73
    8, 0, 1, 1, 12, -8, 5, 9, -4,
    -- layer=1 filter=36 channel=74
    15, -8, 1, 5, 6, -10, 9, -7, 3,
    -- layer=1 filter=36 channel=75
    -57, -66, -41, -10, -16, -33, -9, -21, -19,
    -- layer=1 filter=36 channel=76
    -4, -12, 1, 30, 2, -19, 22, 6, 2,
    -- layer=1 filter=36 channel=77
    7, -2, -6, -3, -10, -11, 2, -5, 8,
    -- layer=1 filter=36 channel=78
    -7, 3, 7, -4, 0, 11, -5, 12, 3,
    -- layer=1 filter=36 channel=79
    -14, -12, -8, 6, -22, -6, -6, 10, 25,
    -- layer=1 filter=36 channel=80
    3, 2, -2, 0, -10, 8, 0, -12, -1,
    -- layer=1 filter=36 channel=81
    12, 3, -1, -5, -7, -15, 1, 8, 5,
    -- layer=1 filter=36 channel=82
    -11, 1, -1, -3, -4, 8, -5, -3, -1,
    -- layer=1 filter=36 channel=83
    0, -25, -13, -13, -21, -8, -8, -13, 5,
    -- layer=1 filter=36 channel=84
    -20, -29, -7, 25, -2, 7, 16, 3, 18,
    -- layer=1 filter=36 channel=85
    14, 7, 73, 39, 24, 30, 17, 17, -30,
    -- layer=1 filter=36 channel=86
    1, -5, -14, -3, -1, -3, -17, -10, 1,
    -- layer=1 filter=36 channel=87
    11, -38, 20, -28, -25, -14, 23, 4, -47,
    -- layer=1 filter=36 channel=88
    -2, 5, -6, -6, 5, 16, -8, 3, 13,
    -- layer=1 filter=36 channel=89
    -8, -16, 11, -9, -1, 8, 4, 10, 3,
    -- layer=1 filter=36 channel=90
    16, -27, 23, -3, 13, 28, 26, -15, 11,
    -- layer=1 filter=36 channel=91
    5, 2, -8, -6, 9, 0, -3, -7, 12,
    -- layer=1 filter=36 channel=92
    12, -68, 8, 3, -40, -49, 8, -33, -8,
    -- layer=1 filter=36 channel=93
    8, 8, -6, -7, -8, 8, 6, -5, 8,
    -- layer=1 filter=36 channel=94
    -11, -11, -12, 12, 12, 2, 13, -4, 0,
    -- layer=1 filter=36 channel=95
    -45, -23, -24, 10, 7, -3, 9, -10, 14,
    -- layer=1 filter=36 channel=96
    7, -6, -12, 0, 5, -7, 3, -12, -9,
    -- layer=1 filter=36 channel=97
    7, -3, -9, -10, 2, -1, 2, 0, 4,
    -- layer=1 filter=36 channel=98
    -31, 2, 7, -2, -19, -6, -7, 7, 31,
    -- layer=1 filter=36 channel=99
    35, 7, 5, 25, -21, 31, 17, -9, 30,
    -- layer=1 filter=36 channel=100
    -3, -19, -5, -11, -4, -1, 10, 0, 23,
    -- layer=1 filter=36 channel=101
    2, -9, 0, -2, 1, -14, 8, 8, -3,
    -- layer=1 filter=36 channel=102
    -14, -15, -12, 4, -12, 3, -11, -11, -8,
    -- layer=1 filter=36 channel=103
    -21, -11, -23, -21, -19, -8, -22, 2, -6,
    -- layer=1 filter=36 channel=104
    19, 12, 29, 22, 3, 22, 29, 1, -19,
    -- layer=1 filter=36 channel=105
    -1, -5, -12, 12, -2, 0, -5, -14, 7,
    -- layer=1 filter=36 channel=106
    -9, -4, 3, 0, 14, 13, 3, 0, 3,
    -- layer=1 filter=36 channel=107
    -13, -3, 0, -13, -5, -2, -7, -1, -2,
    -- layer=1 filter=36 channel=108
    17, -15, 50, 1, 9, 31, 7, -15, 5,
    -- layer=1 filter=36 channel=109
    10, -1, 8, -3, 1, 0, -6, 2, 4,
    -- layer=1 filter=36 channel=110
    3, -4, -9, -6, 2, -9, 4, 7, -6,
    -- layer=1 filter=36 channel=111
    -46, -29, -35, 16, 0, 3, 11, 0, 0,
    -- layer=1 filter=36 channel=112
    -15, 0, -16, 38, 10, -4, 4, -3, 18,
    -- layer=1 filter=36 channel=113
    -4, -9, 21, -1, 6, 15, -5, -2, 29,
    -- layer=1 filter=36 channel=114
    -26, -50, -62, -21, -58, -55, -42, -39, -3,
    -- layer=1 filter=36 channel=115
    -13, -7, 2, 1, -21, 0, -12, -17, 3,
    -- layer=1 filter=36 channel=116
    -3, 0, -7, 6, -9, -8, 6, -4, -9,
    -- layer=1 filter=36 channel=117
    -49, -19, -38, 11, -13, 9, 9, -1, 18,
    -- layer=1 filter=36 channel=118
    -36, -32, -24, 12, 0, -9, 10, -2, 10,
    -- layer=1 filter=36 channel=119
    26, -8, 38, -2, 23, 37, 17, 6, 6,
    -- layer=1 filter=36 channel=120
    -3, 11, -4, 13, -6, 8, -5, -13, 7,
    -- layer=1 filter=36 channel=121
    -34, -56, -39, -30, -47, -46, -18, -10, -22,
    -- layer=1 filter=36 channel=122
    -7, 2, 9, 8, 9, -5, 3, -3, 1,
    -- layer=1 filter=36 channel=123
    -52, -51, -48, -33, -27, -43, -41, -14, -34,
    -- layer=1 filter=36 channel=124
    -6, 4, 1, -5, 3, -3, 1, -10, 5,
    -- layer=1 filter=36 channel=125
    -12, -25, 6, 7, -22, 0, -27, -22, 6,
    -- layer=1 filter=36 channel=126
    -37, -31, 0, -45, -34, -9, -11, -6, 13,
    -- layer=1 filter=36 channel=127
    -48, -30, -37, 8, -5, -16, 8, 1, 3,
    -- layer=1 filter=37 channel=0
    1, -7, -9, 15, 5, -25, 8, 4, 23,
    -- layer=1 filter=37 channel=1
    -28, -39, -39, 66, 54, 46, -15, -42, -26,
    -- layer=1 filter=37 channel=2
    8, 6, 24, -54, -41, -6, 50, 39, 17,
    -- layer=1 filter=37 channel=3
    9, 9, -1, 2, -8, 1, 2, 1, -11,
    -- layer=1 filter=37 channel=4
    10, -12, 1, -4, 2, -5, 0, 16, 3,
    -- layer=1 filter=37 channel=5
    -4, -18, -23, 45, 69, 68, -57, -88, -53,
    -- layer=1 filter=37 channel=6
    -37, -24, -47, -8, -50, 15, 64, 47, 44,
    -- layer=1 filter=37 channel=7
    -4, -39, -66, -28, -70, -70, -18, 7, -1,
    -- layer=1 filter=37 channel=8
    -9, -34, -41, 68, 74, 66, -66, -47, -24,
    -- layer=1 filter=37 channel=9
    -21, 14, 44, -6, -71, -13, 37, -35, -28,
    -- layer=1 filter=37 channel=10
    3, -36, -47, -1, -51, -58, -14, 4, -31,
    -- layer=1 filter=37 channel=11
    -10, 13, -4, -13, 18, 14, 0, 11, 36,
    -- layer=1 filter=37 channel=12
    17, -36, -42, -2, -22, -24, 0, 13, 0,
    -- layer=1 filter=37 channel=13
    -38, -44, -46, 30, 16, 20, 30, 16, 28,
    -- layer=1 filter=37 channel=14
    1, -19, -48, -22, -45, -48, -9, 17, 40,
    -- layer=1 filter=37 channel=15
    -42, -63, -32, 18, 38, 61, 23, -35, 39,
    -- layer=1 filter=37 channel=16
    14, -18, -37, 75, 76, 85, -82, -68, -53,
    -- layer=1 filter=37 channel=17
    -6, -24, -21, 31, 32, 17, 0, 25, 43,
    -- layer=1 filter=37 channel=18
    -23, -53, -13, -95, -49, -50, 36, 34, 7,
    -- layer=1 filter=37 channel=19
    -10, -14, 4, 40, 100, 72, 15, -33, -48,
    -- layer=1 filter=37 channel=20
    -48, -56, -71, 22, 8, 12, 20, 11, 6,
    -- layer=1 filter=37 channel=21
    -4, -12, -14, 44, 2, 5, 15, 17, 19,
    -- layer=1 filter=37 channel=22
    -70, -71, -65, 39, 27, 16, -3, 3, 3,
    -- layer=1 filter=37 channel=23
    -32, -8, -13, -1, 0, 35, 4, -11, 35,
    -- layer=1 filter=37 channel=24
    -8, -28, -23, 4, 27, 28, -15, -22, 1,
    -- layer=1 filter=37 channel=25
    3, -22, -53, 63, 43, 31, -31, -12, -54,
    -- layer=1 filter=37 channel=26
    -38, -47, -34, -4, 30, 31, 10, -4, 11,
    -- layer=1 filter=37 channel=27
    -15, -18, -4, -21, 2, 28, -21, -25, -5,
    -- layer=1 filter=37 channel=28
    6, -34, -58, 44, 0, -38, -5, 11, -26,
    -- layer=1 filter=37 channel=29
    -45, -28, -24, -26, -14, 6, -6, 30, 32,
    -- layer=1 filter=37 channel=30
    -35, -60, -22, -81, -62, -45, 37, 35, -7,
    -- layer=1 filter=37 channel=31
    -3, -21, -39, -10, -41, -12, 28, 22, 33,
    -- layer=1 filter=37 channel=32
    -11, -20, 2, -16, -40, -10, 37, -21, 12,
    -- layer=1 filter=37 channel=33
    -9, -9, -2, 14, 21, 1, 9, 4, -12,
    -- layer=1 filter=37 channel=34
    3, 8, 4, 30, 15, 20, 30, 34, 24,
    -- layer=1 filter=37 channel=35
    5, 11, 11, 19, 30, 19, -10, 3, 6,
    -- layer=1 filter=37 channel=36
    -6, 11, 6, -23, 15, 10, -3, 5, 15,
    -- layer=1 filter=37 channel=37
    25, -25, -26, 48, 61, 64, -61, -65, -60,
    -- layer=1 filter=37 channel=38
    -26, -36, -54, 0, -3, -10, 41, 35, 12,
    -- layer=1 filter=37 channel=39
    30, 21, 6, 26, 44, 68, -14, -24, 3,
    -- layer=1 filter=37 channel=40
    -22, -63, -67, -25, -10, -6, 23, 30, 22,
    -- layer=1 filter=37 channel=41
    -6, -11, 28, 10, -67, 13, 38, -44, -8,
    -- layer=1 filter=37 channel=42
    8, 14, 7, -35, -12, -11, 47, 50, 25,
    -- layer=1 filter=37 channel=43
    -9, -41, -57, 78, 75, 62, -34, -47, -43,
    -- layer=1 filter=37 channel=44
    -35, -42, -27, -1, -3, 32, 8, 0, 29,
    -- layer=1 filter=37 channel=45
    -14, -42, -18, 18, 43, 53, -6, 7, 23,
    -- layer=1 filter=37 channel=46
    3, -21, -4, 67, 119, 93, 40, 47, 14,
    -- layer=1 filter=37 channel=47
    -12, 6, 14, 27, -22, 17, 46, -24, 59,
    -- layer=1 filter=37 channel=48
    -34, -29, -28, -19, -12, -14, 43, 12, 17,
    -- layer=1 filter=37 channel=49
    -4, 18, 22, 0, -36, 26, 66, 29, 36,
    -- layer=1 filter=37 channel=50
    9, 2, 38, 29, 2, 5, 0, -9, 5,
    -- layer=1 filter=37 channel=51
    -13, -18, -42, -24, -49, -55, 34, 13, 20,
    -- layer=1 filter=37 channel=52
    8, 6, -5, 4, -5, -5, 19, 7, 18,
    -- layer=1 filter=37 channel=53
    -1, 9, 9, 17, 18, 15, 10, 5, 16,
    -- layer=1 filter=37 channel=54
    32, -22, -36, 52, 38, 35, -28, -40, -92,
    -- layer=1 filter=37 channel=55
    -5, 22, 12, 2, 15, 29, -37, -28, 12,
    -- layer=1 filter=37 channel=56
    -9, 4, 5, -1, -2, 0, 1, 3, -5,
    -- layer=1 filter=37 channel=57
    0, -41, -68, -3, -42, -43, 1, 32, -12,
    -- layer=1 filter=37 channel=58
    -35, -29, -31, -30, -60, -26, 8, -16, 20,
    -- layer=1 filter=37 channel=59
    -2, -7, -1, -4, 7, 1, -3, -19, 3,
    -- layer=1 filter=37 channel=60
    -8, -26, -11, -5, 1, -19, -22, -20, -11,
    -- layer=1 filter=37 channel=61
    -11, 1, 0, -1, 6, -3, -4, 0, 5,
    -- layer=1 filter=37 channel=62
    9, -31, -40, 72, 69, 71, -70, -66, -40,
    -- layer=1 filter=37 channel=63
    -21, -4, -8, -32, -10, 5, 18, 21, 23,
    -- layer=1 filter=37 channel=64
    -66, -27, -55, 21, -7, -24, 29, 11, 19,
    -- layer=1 filter=37 channel=65
    -19, -40, -45, 16, 13, 5, 31, 24, 4,
    -- layer=1 filter=37 channel=66
    -10, 12, -2, -11, 6, 6, -9, 5, 3,
    -- layer=1 filter=37 channel=67
    -29, -20, -33, -24, -41, 9, 38, 41, 24,
    -- layer=1 filter=37 channel=68
    -49, -41, -37, -21, -4, -6, 11, 13, 14,
    -- layer=1 filter=37 channel=69
    2, -24, -27, 54, 69, 76, -68, -51, -22,
    -- layer=1 filter=37 channel=70
    39, 28, -16, -54, -83, 31, 69, 52, 49,
    -- layer=1 filter=37 channel=71
    10, 11, -7, 24, 31, 42, -9, -21, -37,
    -- layer=1 filter=37 channel=72
    -51, -70, -20, 32, 12, 7, 48, -6, -7,
    -- layer=1 filter=37 channel=73
    -6, -8, 4, -9, 0, -5, -10, 5, 2,
    -- layer=1 filter=37 channel=74
    -19, 9, -16, -35, 1, -15, 28, 17, -10,
    -- layer=1 filter=37 channel=75
    -31, -55, -43, -38, -37, -2, -19, 13, 5,
    -- layer=1 filter=37 channel=76
    11, 4, 0, -4, -14, -15, 27, 19, 19,
    -- layer=1 filter=37 channel=77
    -16, -19, -16, 20, 18, -2, 18, 19, 10,
    -- layer=1 filter=37 channel=78
    -1, -2, -19, 21, -21, -20, 6, 24, 10,
    -- layer=1 filter=37 channel=79
    14, -19, -48, 59, 67, 69, -53, -51, -9,
    -- layer=1 filter=37 channel=80
    -14, -7, 2, 3, 12, 7, -3, 10, -4,
    -- layer=1 filter=37 channel=81
    -8, -6, -30, 43, 40, 28, -18, 0, -2,
    -- layer=1 filter=37 channel=82
    -24, -10, -22, 20, 1, -2, 26, 30, 13,
    -- layer=1 filter=37 channel=83
    -28, -56, -61, 16, 65, 54, -12, 2, 28,
    -- layer=1 filter=37 channel=84
    -44, -28, -3, -42, -32, -41, 42, 23, -3,
    -- layer=1 filter=37 channel=85
    -2, 15, -9, 0, -23, 22, 22, -20, 41,
    -- layer=1 filter=37 channel=86
    -7, 5, 16, 11, 14, 25, -35, -11, -15,
    -- layer=1 filter=37 channel=87
    -24, 10, 0, 72, 67, 19, 55, 6, 6,
    -- layer=1 filter=37 channel=88
    14, 1, 23, -5, 0, 18, 53, 30, 34,
    -- layer=1 filter=37 channel=89
    -21, -25, -11, -9, -8, -22, 34, 36, 18,
    -- layer=1 filter=37 channel=90
    -23, -35, -61, -12, 21, 36, 3, 6, 31,
    -- layer=1 filter=37 channel=91
    -41, -40, -66, -15, -37, -51, 52, 38, 29,
    -- layer=1 filter=37 channel=92
    10, -46, -21, 6, 24, 39, 6, -30, -13,
    -- layer=1 filter=37 channel=93
    -16, -27, -18, 18, 2, -4, -2, -5, -6,
    -- layer=1 filter=37 channel=94
    -7, 0, -10, 7, -12, -16, 1, 5, 25,
    -- layer=1 filter=37 channel=95
    -45, -38, -24, -87, -73, -45, 37, 19, -8,
    -- layer=1 filter=37 channel=96
    -10, -16, -11, -5, -9, -8, 14, 1, -4,
    -- layer=1 filter=37 channel=97
    -21, -28, -23, 31, 11, 11, 7, 0, -3,
    -- layer=1 filter=37 channel=98
    -24, -60, -75, 80, 68, 57, -6, -7, 6,
    -- layer=1 filter=37 channel=99
    -14, -26, -47, -21, -37, -25, 26, 27, 9,
    -- layer=1 filter=37 channel=100
    15, 21, 24, -15, -10, 31, 25, 3, 6,
    -- layer=1 filter=37 channel=101
    -52, -38, -28, -12, -36, -40, 40, 28, 22,
    -- layer=1 filter=37 channel=102
    -11, -4, -16, -12, -36, -52, 48, 45, 30,
    -- layer=1 filter=37 channel=103
    -5, -7, -7, -37, -21, 8, 30, 35, 35,
    -- layer=1 filter=37 channel=104
    -23, 9, 13, -34, -29, 10, 15, -3, 29,
    -- layer=1 filter=37 channel=105
    -17, -18, -19, 4, -2, -26, 8, 14, 12,
    -- layer=1 filter=37 channel=106
    -49, -42, -19, -31, -42, -21, 67, 48, 37,
    -- layer=1 filter=37 channel=107
    12, -2, 0, 0, 8, 20, -6, -3, -8,
    -- layer=1 filter=37 channel=108
    -12, -54, -13, 3, 9, 43, -4, -26, 21,
    -- layer=1 filter=37 channel=109
    -11, 7, -2, 1, -4, 4, -8, 6, -7,
    -- layer=1 filter=37 channel=110
    -4, -22, -15, -11, -3, -12, 4, 20, 6,
    -- layer=1 filter=37 channel=111
    -1, -47, -21, -72, -42, -46, 26, 22, 16,
    -- layer=1 filter=37 channel=112
    -4, -2, 2, -22, 26, -4, 19, 2, 9,
    -- layer=1 filter=37 channel=113
    14, -34, -12, -11, -7, -10, 23, 43, 6,
    -- layer=1 filter=37 channel=114
    28, -3, -10, 60, 76, 78, -84, -108, -45,
    -- layer=1 filter=37 channel=115
    4, -23, -25, 9, -18, 1, -29, -8, -10,
    -- layer=1 filter=37 channel=116
    -7, -6, -1, -4, -6, -7, 11, 0, -6,
    -- layer=1 filter=37 channel=117
    -28, -1, -39, 20, 64, 22, 16, 27, 14,
    -- layer=1 filter=37 channel=118
    -14, -15, -14, -67, -47, -61, 60, 36, 6,
    -- layer=1 filter=37 channel=119
    -11, -40, -27, -19, -38, -16, 27, 1, 33,
    -- layer=1 filter=37 channel=120
    -21, -28, -33, 21, 8, -2, 20, 19, 7,
    -- layer=1 filter=37 channel=121
    -33, -26, -16, -32, 36, 66, -6, 27, 14,
    -- layer=1 filter=37 channel=122
    6, 5, -4, -5, -3, 3, -5, -1, -3,
    -- layer=1 filter=37 channel=123
    -17, -5, 17, -35, -3, 49, -28, 0, -14,
    -- layer=1 filter=37 channel=124
    -5, 11, 6, 20, 9, 2, -15, -4, 0,
    -- layer=1 filter=37 channel=125
    35, 17, 1, -65, -83, -8, 57, 59, 31,
    -- layer=1 filter=37 channel=126
    -75, -84, -70, 80, 78, 51, 18, 11, 26,
    -- layer=1 filter=37 channel=127
    -31, -35, -9, -100, -63, -60, 32, 24, 1,
    -- layer=1 filter=38 channel=0
    -1, -4, -11, 4, -7, -11, -10, 8, 1,
    -- layer=1 filter=38 channel=1
    0, -7, 5, -4, 2, -11, -1, 5, 8,
    -- layer=1 filter=38 channel=2
    1, -8, -5, 3, 0, -11, -4, -11, 4,
    -- layer=1 filter=38 channel=3
    -6, -9, 4, 7, 7, 4, -7, 0, 1,
    -- layer=1 filter=38 channel=4
    6, -3, -6, 7, 6, -4, 0, 0, 0,
    -- layer=1 filter=38 channel=5
    2, 6, -1, -6, 4, 0, 6, -10, 5,
    -- layer=1 filter=38 channel=6
    4, -6, 0, 6, -8, -3, 7, -2, -11,
    -- layer=1 filter=38 channel=7
    -15, -2, -12, 3, 8, 1, 4, -1, 5,
    -- layer=1 filter=38 channel=8
    0, -11, 8, -9, 6, -4, 3, -1, 4,
    -- layer=1 filter=38 channel=9
    -7, 0, 0, -5, 9, 4, 8, 9, -4,
    -- layer=1 filter=38 channel=10
    0, -9, 6, 4, 4, -3, 2, -7, 0,
    -- layer=1 filter=38 channel=11
    6, -3, -8, -5, -8, -7, 6, -4, -5,
    -- layer=1 filter=38 channel=12
    10, -4, 4, 0, 3, 8, 10, 7, 7,
    -- layer=1 filter=38 channel=13
    9, 9, -3, 1, 0, 8, -9, 0, -7,
    -- layer=1 filter=38 channel=14
    0, 6, -10, 4, 6, -4, -9, 0, -6,
    -- layer=1 filter=38 channel=15
    7, 0, -9, -5, -1, 7, 6, 2, 0,
    -- layer=1 filter=38 channel=16
    6, 1, -10, -5, 1, -6, 2, 4, 4,
    -- layer=1 filter=38 channel=17
    -11, 5, 2, 3, -12, -7, -7, 5, -5,
    -- layer=1 filter=38 channel=18
    3, -9, -11, 0, -12, -13, -5, 5, 4,
    -- layer=1 filter=38 channel=19
    -2, 1, -4, -3, -4, -9, -2, 7, -9,
    -- layer=1 filter=38 channel=20
    0, -6, 2, 7, 5, -2, -1, -11, 0,
    -- layer=1 filter=38 channel=21
    -5, -7, 0, 9, 0, 12, 10, -8, -3,
    -- layer=1 filter=38 channel=22
    -10, 7, -2, 3, -5, -10, -12, -12, -6,
    -- layer=1 filter=38 channel=23
    2, -8, -10, 2, 8, -3, -11, -4, -1,
    -- layer=1 filter=38 channel=24
    7, 7, 1, 2, -9, 5, -8, 4, -9,
    -- layer=1 filter=38 channel=25
    7, -13, -3, 5, -6, 4, 0, -11, -10,
    -- layer=1 filter=38 channel=26
    -8, -10, 2, 7, -2, 0, 5, -8, -9,
    -- layer=1 filter=38 channel=27
    3, -5, 4, 5, -8, -9, 4, 1, -5,
    -- layer=1 filter=38 channel=28
    9, 0, -7, 0, 0, 1, 0, -1, -6,
    -- layer=1 filter=38 channel=29
    -2, 1, -3, 7, -6, 8, 0, 6, 9,
    -- layer=1 filter=38 channel=30
    1, -7, -5, 4, -13, -1, -8, 7, -11,
    -- layer=1 filter=38 channel=31
    -13, -1, -13, -5, -8, 0, 2, 2, 0,
    -- layer=1 filter=38 channel=32
    -6, 2, 6, 6, 0, -1, 5, -4, -11,
    -- layer=1 filter=38 channel=33
    -10, -7, 0, 2, 0, 0, -8, -2, -6,
    -- layer=1 filter=38 channel=34
    5, 2, -4, 5, -4, -10, 8, -8, -7,
    -- layer=1 filter=38 channel=35
    -6, -11, -1, -10, 3, -11, 5, 0, -5,
    -- layer=1 filter=38 channel=36
    -10, -11, -13, 2, -5, -9, -7, -7, -4,
    -- layer=1 filter=38 channel=37
    -3, 0, -13, 8, 4, -12, -9, -7, 6,
    -- layer=1 filter=38 channel=38
    8, 4, 1, 3, 0, -2, -3, 8, -8,
    -- layer=1 filter=38 channel=39
    -2, 6, -2, -9, 4, -3, 3, -5, 4,
    -- layer=1 filter=38 channel=40
    3, 4, -9, 1, 0, -1, -13, -12, -5,
    -- layer=1 filter=38 channel=41
    -5, -4, 3, -3, -4, 9, -1, 1, -8,
    -- layer=1 filter=38 channel=42
    -3, -4, -10, -3, 8, -9, -10, -2, -4,
    -- layer=1 filter=38 channel=43
    6, -3, -1, -10, 8, 4, 4, 1, 4,
    -- layer=1 filter=38 channel=44
    6, -11, -4, 8, -5, -4, 7, -8, -7,
    -- layer=1 filter=38 channel=45
    7, 6, 1, 1, 8, -6, 0, -2, 0,
    -- layer=1 filter=38 channel=46
    -4, -12, -3, 4, 0, 2, 6, -6, 0,
    -- layer=1 filter=38 channel=47
    8, 5, -3, 7, -6, -11, -5, 7, 0,
    -- layer=1 filter=38 channel=48
    -2, 8, -8, -10, -4, -11, 4, 3, -9,
    -- layer=1 filter=38 channel=49
    -5, -10, -10, 5, -6, 10, 0, 0, 2,
    -- layer=1 filter=38 channel=50
    3, -3, -7, 5, -1, -2, -3, 4, -5,
    -- layer=1 filter=38 channel=51
    5, 2, -2, -6, 5, 2, 3, 4, -2,
    -- layer=1 filter=38 channel=52
    -5, 0, 0, 3, -4, 3, -6, -6, 0,
    -- layer=1 filter=38 channel=53
    -1, -5, 7, -10, -3, -7, 5, 0, 5,
    -- layer=1 filter=38 channel=54
    -9, -1, -7, -8, -1, 2, -7, -6, -5,
    -- layer=1 filter=38 channel=55
    -2, 4, 0, -11, 5, -11, 8, -6, -7,
    -- layer=1 filter=38 channel=56
    -2, 9, 0, 9, 8, 4, 8, -9, 0,
    -- layer=1 filter=38 channel=57
    -9, -4, 4, -4, 0, 1, -11, 4, 6,
    -- layer=1 filter=38 channel=58
    -6, 9, -8, 0, -11, -3, -4, 0, 6,
    -- layer=1 filter=38 channel=59
    2, 5, 4, -9, 0, 4, -11, 3, 3,
    -- layer=1 filter=38 channel=60
    -7, -8, 6, -5, -9, -5, 6, 7, 4,
    -- layer=1 filter=38 channel=61
    2, 7, 6, -8, 0, -6, 10, -11, -5,
    -- layer=1 filter=38 channel=62
    -2, 4, -2, -11, 2, -6, 5, 4, -9,
    -- layer=1 filter=38 channel=63
    -8, 2, -7, -4, -2, 1, 3, -4, -10,
    -- layer=1 filter=38 channel=64
    -9, -7, 5, -3, -6, -6, -3, 8, 0,
    -- layer=1 filter=38 channel=65
    -12, 0, -5, -4, 0, 8, -6, 7, 1,
    -- layer=1 filter=38 channel=66
    -11, -8, -12, 2, -4, -4, -10, -4, -8,
    -- layer=1 filter=38 channel=67
    -3, -1, -3, -7, -12, 0, 4, 7, 0,
    -- layer=1 filter=38 channel=68
    3, -6, 2, -3, -3, 1, 1, -4, 0,
    -- layer=1 filter=38 channel=69
    1, -5, 0, 0, -9, 5, 6, -2, -6,
    -- layer=1 filter=38 channel=70
    -4, 5, -11, 3, -13, -10, 6, 4, -11,
    -- layer=1 filter=38 channel=71
    -11, 1, 8, -8, 7, 4, -11, 6, -9,
    -- layer=1 filter=38 channel=72
    -8, 6, 5, 7, -9, 7, -5, -10, -4,
    -- layer=1 filter=38 channel=73
    -4, -7, -10, 1, -4, -3, -3, 0, -12,
    -- layer=1 filter=38 channel=74
    -6, 2, -2, 0, -7, 5, 6, 5, -11,
    -- layer=1 filter=38 channel=75
    1, -2, -7, -8, 0, 0, -2, 6, -6,
    -- layer=1 filter=38 channel=76
    -1, -7, 0, -1, 0, 7, 0, -8, -11,
    -- layer=1 filter=38 channel=77
    -3, 6, 0, -3, 2, -5, -7, -2, -3,
    -- layer=1 filter=38 channel=78
    -6, -7, 6, 5, 3, -3, 7, 0, -8,
    -- layer=1 filter=38 channel=79
    0, 2, -1, 0, 2, -11, -7, -8, 0,
    -- layer=1 filter=38 channel=80
    -8, 9, -7, -4, 5, 0, -11, 0, 4,
    -- layer=1 filter=38 channel=81
    9, -3, -3, 6, 1, -5, 2, 6, -11,
    -- layer=1 filter=38 channel=82
    -9, 2, 4, 2, 0, 7, 4, 0, 4,
    -- layer=1 filter=38 channel=83
    -3, -4, 7, -8, 3, 2, 4, 6, 6,
    -- layer=1 filter=38 channel=84
    -1, -3, -5, -8, -3, -2, -7, 7, -7,
    -- layer=1 filter=38 channel=85
    -10, 7, -8, -1, 6, 5, 2, -4, 7,
    -- layer=1 filter=38 channel=86
    2, -7, 0, 3, 0, 6, -2, -6, 2,
    -- layer=1 filter=38 channel=87
    7, 1, -11, -9, 0, -3, -5, 0, 9,
    -- layer=1 filter=38 channel=88
    4, -6, -5, -8, 0, -5, 4, -2, 7,
    -- layer=1 filter=38 channel=89
    -7, 0, -5, 8, 0, 4, -9, -4, 8,
    -- layer=1 filter=38 channel=90
    -6, -11, 8, -8, 7, -11, -4, -3, 6,
    -- layer=1 filter=38 channel=91
    6, 5, -3, -6, 0, -5, 4, -1, 8,
    -- layer=1 filter=38 channel=92
    -3, 0, 9, -7, -7, 3, -11, -1, -10,
    -- layer=1 filter=38 channel=93
    -9, -1, -6, 2, -7, 7, -1, -10, -6,
    -- layer=1 filter=38 channel=94
    5, 1, -10, -6, -3, 3, -8, -1, -3,
    -- layer=1 filter=38 channel=95
    -3, 2, -11, 0, 8, 4, -5, 0, -1,
    -- layer=1 filter=38 channel=96
    -5, -8, -10, 0, -6, 7, -9, 3, 7,
    -- layer=1 filter=38 channel=97
    -8, 7, -7, 2, 7, 0, 0, -4, 0,
    -- layer=1 filter=38 channel=98
    1, -1, 1, 0, -11, -9, -10, -7, 2,
    -- layer=1 filter=38 channel=99
    6, -5, 2, -1, -3, -3, -5, -10, -1,
    -- layer=1 filter=38 channel=100
    3, -11, -1, -6, -9, 6, 0, 2, 3,
    -- layer=1 filter=38 channel=101
    -5, -9, 1, 5, -3, 5, -3, -6, 0,
    -- layer=1 filter=38 channel=102
    -3, 0, 0, 7, -2, -2, 3, 2, -5,
    -- layer=1 filter=38 channel=103
    -8, -3, -11, -3, 4, -11, -3, -10, 0,
    -- layer=1 filter=38 channel=104
    5, 7, -9, 0, 5, 6, 0, 0, -5,
    -- layer=1 filter=38 channel=105
    4, 7, -10, -7, -8, 8, 8, 8, 8,
    -- layer=1 filter=38 channel=106
    3, -5, -6, -5, 5, -7, 5, -9, 1,
    -- layer=1 filter=38 channel=107
    4, -3, 0, -8, 0, -3, -1, 4, -2,
    -- layer=1 filter=38 channel=108
    -1, 6, -6, -6, -11, -3, 7, 3, -3,
    -- layer=1 filter=38 channel=109
    -4, 0, -1, 3, -9, -10, 8, -7, 7,
    -- layer=1 filter=38 channel=110
    -6, -3, 0, 8, -3, -3, 6, -8, -9,
    -- layer=1 filter=38 channel=111
    -8, -7, -4, -10, 7, -11, -5, -6, -7,
    -- layer=1 filter=38 channel=112
    6, 0, -11, 1, 8, -10, -2, 6, 6,
    -- layer=1 filter=38 channel=113
    4, -2, -1, 3, 7, -4, 1, 4, 0,
    -- layer=1 filter=38 channel=114
    -6, -6, 6, 5, 8, 8, -6, 7, 1,
    -- layer=1 filter=38 channel=115
    8, -3, 0, 3, 3, -10, -4, -11, -9,
    -- layer=1 filter=38 channel=116
    5, 10, 1, -7, 10, 4, 10, 0, 1,
    -- layer=1 filter=38 channel=117
    3, 6, -1, 0, 1, -10, 7, 5, -6,
    -- layer=1 filter=38 channel=118
    2, -4, 2, -4, 3, 2, 2, 9, 3,
    -- layer=1 filter=38 channel=119
    2, 2, -10, -4, -4, -7, -8, -4, -1,
    -- layer=1 filter=38 channel=120
    1, -3, -1, -4, -12, 1, -4, 7, 7,
    -- layer=1 filter=38 channel=121
    -9, -6, -9, 7, 8, 1, -1, -3, -6,
    -- layer=1 filter=38 channel=122
    8, 0, -10, 1, 4, -7, -4, 0, -4,
    -- layer=1 filter=38 channel=123
    -3, -5, -1, 0, -5, 0, -6, 5, 8,
    -- layer=1 filter=38 channel=124
    -12, 1, 4, 7, -2, 0, 6, -9, -6,
    -- layer=1 filter=38 channel=125
    -12, 3, -12, 2, -10, -4, -4, -1, -3,
    -- layer=1 filter=38 channel=126
    3, 4, 8, -6, -1, -6, 4, -5, -4,
    -- layer=1 filter=38 channel=127
    -13, -1, -8, -12, -15, -5, 0, 1, 5,
    -- layer=1 filter=39 channel=0
    -3, -12, -2, 12, 9, -8, -4, -2, 8,
    -- layer=1 filter=39 channel=1
    -6, -5, -2, 0, 0, 13, 38, 5, 2,
    -- layer=1 filter=39 channel=2
    -9, -22, -52, -7, -25, -21, -7, -16, -23,
    -- layer=1 filter=39 channel=3
    -2, 10, 0, 4, -3, -1, -16, 5, -7,
    -- layer=1 filter=39 channel=4
    -8, -6, 5, -2, 6, 0, 0, -7, 2,
    -- layer=1 filter=39 channel=5
    -2, -19, -22, -22, -35, -10, 23, -5, 13,
    -- layer=1 filter=39 channel=6
    0, -2, 1, -2, -26, -11, -26, -10, -9,
    -- layer=1 filter=39 channel=7
    6, 20, -27, 10, 0, 22, 0, 10, 7,
    -- layer=1 filter=39 channel=8
    -14, -14, -42, -16, -27, 4, 1, -23, 16,
    -- layer=1 filter=39 channel=9
    -21, -10, 9, -21, -36, -9, 2, -10, 2,
    -- layer=1 filter=39 channel=10
    -9, 13, -26, 2, -15, 22, -27, 0, -7,
    -- layer=1 filter=39 channel=11
    -6, -18, 2, -5, 5, 0, 0, -17, -19,
    -- layer=1 filter=39 channel=12
    -64, -35, -33, -19, -81, -12, -56, -48, 4,
    -- layer=1 filter=39 channel=13
    15, 12, 3, -3, -8, 10, 7, 4, -2,
    -- layer=1 filter=39 channel=14
    -29, 16, -39, -4, -51, -42, -33, -30, -11,
    -- layer=1 filter=39 channel=15
    -8, -44, -28, -19, -80, -31, 20, -33, -35,
    -- layer=1 filter=39 channel=16
    -5, -20, -52, -4, -18, -3, 10, -11, 12,
    -- layer=1 filter=39 channel=17
    7, 6, -4, 12, 11, 9, 7, -5, 1,
    -- layer=1 filter=39 channel=18
    -18, -26, -31, 16, 5, -18, -15, -3, 0,
    -- layer=1 filter=39 channel=19
    -18, -32, -12, -7, -23, 16, 36, 10, 51,
    -- layer=1 filter=39 channel=20
    16, 3, 6, 14, 12, 3, 23, 19, 2,
    -- layer=1 filter=39 channel=21
    -8, 2, -3, -20, 3, -9, 10, -10, 4,
    -- layer=1 filter=39 channel=22
    16, -3, 9, 3, -8, -4, 19, -13, 7,
    -- layer=1 filter=39 channel=23
    -36, -4, 8, -3, -7, 27, -4, -14, 20,
    -- layer=1 filter=39 channel=24
    -27, 1, 3, -15, -14, 0, -1, 8, -9,
    -- layer=1 filter=39 channel=25
    9, 18, -25, -8, 0, 11, 5, 11, 17,
    -- layer=1 filter=39 channel=26
    10, -2, 9, 5, 4, 16, 21, 13, -8,
    -- layer=1 filter=39 channel=27
    -31, -35, -39, -48, -35, -35, -57, -70, -66,
    -- layer=1 filter=39 channel=28
    -3, 21, -11, 3, 9, 6, -15, 9, 5,
    -- layer=1 filter=39 channel=29
    -12, -5, -9, -25, -16, -20, -22, -28, -31,
    -- layer=1 filter=39 channel=30
    -35, -43, -26, -8, -33, -3, 5, 17, -7,
    -- layer=1 filter=39 channel=31
    -5, -2, -23, -3, -29, -20, -16, -29, -8,
    -- layer=1 filter=39 channel=32
    -2, 9, 27, -2, 15, -4, 17, 7, -38,
    -- layer=1 filter=39 channel=33
    -1, -4, -4, -12, -4, -5, -13, 4, -4,
    -- layer=1 filter=39 channel=34
    -4, -21, -11, -28, -39, -10, -6, -19, -4,
    -- layer=1 filter=39 channel=35
    8, -6, 10, 2, -2, -4, 14, -4, -2,
    -- layer=1 filter=39 channel=36
    -10, -1, 8, 10, -5, -15, -14, -1, -13,
    -- layer=1 filter=39 channel=37
    2, -21, -35, -1, -20, 7, 28, -6, 14,
    -- layer=1 filter=39 channel=38
    16, 4, -7, -4, 8, -10, 11, 13, 0,
    -- layer=1 filter=39 channel=39
    9, 7, -9, 0, 1, 10, 3, -3, 5,
    -- layer=1 filter=39 channel=40
    2, 3, -5, 11, -12, 9, -7, 6, 15,
    -- layer=1 filter=39 channel=41
    -6, -1, 51, 7, -12, -11, 5, -13, -31,
    -- layer=1 filter=39 channel=42
    -10, -38, -34, 12, -22, -19, -11, -8, -26,
    -- layer=1 filter=39 channel=43
    -18, -9, -33, -8, -20, -5, 21, -20, 22,
    -- layer=1 filter=39 channel=44
    15, 15, 4, 0, 8, -3, 28, -5, -24,
    -- layer=1 filter=39 channel=45
    3, 7, -13, -12, -3, 4, 15, -10, -13,
    -- layer=1 filter=39 channel=46
    -18, -40, -26, -9, -52, -21, 48, 34, 51,
    -- layer=1 filter=39 channel=47
    -17, 0, 30, -20, -11, 15, -14, -11, -8,
    -- layer=1 filter=39 channel=48
    -8, 5, -1, -7, 0, 6, -2, 0, 0,
    -- layer=1 filter=39 channel=49
    5, -2, 17, 10, -3, 14, -7, -12, 6,
    -- layer=1 filter=39 channel=50
    10, 1, 6, 0, 1, 7, 0, 5, 0,
    -- layer=1 filter=39 channel=51
    -4, 11, -13, -9, 0, -15, -15, 8, -1,
    -- layer=1 filter=39 channel=52
    11, 4, 4, 11, 1, 0, 15, -4, 2,
    -- layer=1 filter=39 channel=53
    9, 9, 10, 4, 6, -1, 7, 21, 8,
    -- layer=1 filter=39 channel=54
    -12, 14, -31, 6, -17, 21, 7, -10, 11,
    -- layer=1 filter=39 channel=55
    0, -12, 6, -9, 0, 1, -29, -13, -16,
    -- layer=1 filter=39 channel=56
    -1, 5, -12, -5, -7, -8, -9, -1, -11,
    -- layer=1 filter=39 channel=57
    14, 17, -17, 9, -21, 0, -8, 15, -16,
    -- layer=1 filter=39 channel=58
    -35, 2, -18, -4, -28, 56, -9, 13, 1,
    -- layer=1 filter=39 channel=59
    0, -2, 2, 13, 0, -1, 11, 0, 12,
    -- layer=1 filter=39 channel=60
    -13, -3, -6, 2, -3, -19, 6, -3, -9,
    -- layer=1 filter=39 channel=61
    8, -9, 9, -1, -10, 2, -2, -12, -8,
    -- layer=1 filter=39 channel=62
    -3, -24, -51, 0, -13, 16, 23, 3, 21,
    -- layer=1 filter=39 channel=63
    -6, -10, 6, -4, 0, -7, -11, 2, 0,
    -- layer=1 filter=39 channel=64
    14, 10, 10, -11, 8, 5, 5, -5, 1,
    -- layer=1 filter=39 channel=65
    -12, -2, -10, 4, -1, 0, 1, 8, 9,
    -- layer=1 filter=39 channel=66
    4, -9, 10, 8, 1, 6, 7, 0, -5,
    -- layer=1 filter=39 channel=67
    24, 5, 17, 11, -4, 0, -22, -23, -19,
    -- layer=1 filter=39 channel=68
    24, 16, 14, 8, 24, -3, 33, 9, -20,
    -- layer=1 filter=39 channel=69
    -3, -11, -7, -23, -21, -7, 9, -24, 6,
    -- layer=1 filter=39 channel=70
    -18, -30, -5, -19, -33, -22, -67, -53, -50,
    -- layer=1 filter=39 channel=71
    -5, -10, -7, -17, -8, -6, 1, -7, 19,
    -- layer=1 filter=39 channel=72
    -33, -36, -21, -29, -31, -5, 32, 0, 25,
    -- layer=1 filter=39 channel=73
    -4, -1, -4, -6, 9, 6, -2, -11, -6,
    -- layer=1 filter=39 channel=74
    19, 5, 12, 4, 13, -11, 17, 11, -2,
    -- layer=1 filter=39 channel=75
    -45, -61, -71, -12, -66, -39, -18, 0, -4,
    -- layer=1 filter=39 channel=76
    7, -5, 8, 24, 19, -12, 13, 18, 6,
    -- layer=1 filter=39 channel=77
    -10, -9, 3, 2, -5, 5, -7, 0, 13,
    -- layer=1 filter=39 channel=78
    10, 1, -7, 5, 9, 9, 0, -4, -17,
    -- layer=1 filter=39 channel=79
    -7, -16, -30, -1, -27, 8, 24, -14, 19,
    -- layer=1 filter=39 channel=80
    -2, -7, -2, 4, 1, 7, -5, 0, 9,
    -- layer=1 filter=39 channel=81
    -8, -6, -5, -13, -7, 1, -4, -2, 2,
    -- layer=1 filter=39 channel=82
    7, -3, -11, -15, 2, 3, 8, -1, 8,
    -- layer=1 filter=39 channel=83
    12, -1, -5, -2, -33, -9, 19, -21, -5,
    -- layer=1 filter=39 channel=84
    0, -15, 1, 8, 17, -8, 12, 5, 8,
    -- layer=1 filter=39 channel=85
    -26, 4, -4, -11, -17, 33, 1, -14, 5,
    -- layer=1 filter=39 channel=86
    13, 0, 17, 2, 12, -1, 14, -2, 9,
    -- layer=1 filter=39 channel=87
    -31, -39, 1, -32, -17, -5, 22, -28, 15,
    -- layer=1 filter=39 channel=88
    0, -9, -2, 0, 7, 12, 12, 16, 18,
    -- layer=1 filter=39 channel=89
    0, -18, -2, 0, 3, 0, 5, 5, 6,
    -- layer=1 filter=39 channel=90
    16, 5, 9, 9, -9, 10, 28, -5, -23,
    -- layer=1 filter=39 channel=91
    6, 19, 13, 16, 1, 0, -5, 11, 12,
    -- layer=1 filter=39 channel=92
    -13, -46, 3, -35, -71, -80, -37, -26, -109,
    -- layer=1 filter=39 channel=93
    -1, 9, 8, 5, -2, 8, 0, 6, 14,
    -- layer=1 filter=39 channel=94
    -3, 3, -10, 16, -1, 8, -1, 6, 16,
    -- layer=1 filter=39 channel=95
    -16, -38, -20, 0, -9, -24, 19, 6, 1,
    -- layer=1 filter=39 channel=96
    -5, 1, 5, -3, 2, -5, 0, 6, -6,
    -- layer=1 filter=39 channel=97
    -6, -1, -5, 4, 11, 3, 7, 9, -3,
    -- layer=1 filter=39 channel=98
    7, -8, -28, 8, -6, 10, 4, -12, 2,
    -- layer=1 filter=39 channel=99
    -4, -7, -18, 9, 10, -17, -29, 11, -10,
    -- layer=1 filter=39 channel=100
    -4, -2, 7, -14, 8, -26, 14, -2, -9,
    -- layer=1 filter=39 channel=101
    9, 14, 9, 8, -4, 5, 8, 3, 1,
    -- layer=1 filter=39 channel=102
    3, 0, -13, 11, 6, 1, 4, 8, 6,
    -- layer=1 filter=39 channel=103
    0, 2, -11, -8, -17, -6, -14, -17, 0,
    -- layer=1 filter=39 channel=104
    -32, -10, -5, 2, -19, 28, 6, -4, -6,
    -- layer=1 filter=39 channel=105
    1, 9, -9, 12, -5, -1, 9, 1, 6,
    -- layer=1 filter=39 channel=106
    5, 4, 24, 0, -1, -7, 18, 0, -13,
    -- layer=1 filter=39 channel=107
    6, 0, -4, -21, -15, -9, -6, -18, -13,
    -- layer=1 filter=39 channel=108
    -5, -4, 37, 8, 2, 0, 5, 2, -38,
    -- layer=1 filter=39 channel=109
    -7, -5, -5, -1, -8, 6, 1, -10, 6,
    -- layer=1 filter=39 channel=110
    6, 7, -10, 7, 2, 3, -9, 0, 7,
    -- layer=1 filter=39 channel=111
    -8, -21, -32, 20, 11, 10, -11, 21, 15,
    -- layer=1 filter=39 channel=112
    -11, -12, -35, 33, 22, -9, -25, -5, 10,
    -- layer=1 filter=39 channel=113
    -7, -31, -28, -14, -32, -36, -21, -15, -17,
    -- layer=1 filter=39 channel=114
    -49, -68, -65, -70, -80, -61, -39, -87, -31,
    -- layer=1 filter=39 channel=115
    1, 4, -3, 9, 1, -1, -1, -1, 5,
    -- layer=1 filter=39 channel=116
    -2, 1, -10, 5, -11, 7, 4, -5, -7,
    -- layer=1 filter=39 channel=117
    -32, -44, -61, 21, -18, 18, -55, -7, -9,
    -- layer=1 filter=39 channel=118
    -3, -12, -16, 5, 7, 5, 9, 20, 3,
    -- layer=1 filter=39 channel=119
    -7, 7, 9, -2, 4, 14, 16, -5, -31,
    -- layer=1 filter=39 channel=120
    2, 9, 4, -7, -9, 10, 4, 13, 12,
    -- layer=1 filter=39 channel=121
    -49, -56, -35, -26, -82, -40, -6, 8, -17,
    -- layer=1 filter=39 channel=122
    2, -3, -8, -3, 7, 5, -5, 3, 2,
    -- layer=1 filter=39 channel=123
    -40, -46, -20, -33, -37, -19, -1, -10, -14,
    -- layer=1 filter=39 channel=124
    1, -11, -1, -7, -6, 1, 0, -3, -7,
    -- layer=1 filter=39 channel=125
    10, 4, 1, -7, -23, -19, -25, -36, -34,
    -- layer=1 filter=39 channel=126
    -17, -10, -15, -13, -32, -12, 16, -37, 9,
    -- layer=1 filter=39 channel=127
    -8, -35, -31, 22, 3, -12, 14, 13, 12,
    -- layer=1 filter=40 channel=0
    11, 21, 21, 11, 15, 14, 6, 5, 15,
    -- layer=1 filter=40 channel=1
    1, -19, -13, -4, 16, -1, -16, 11, 13,
    -- layer=1 filter=40 channel=2
    -6, 22, 15, 1, 27, 23, -36, -24, 11,
    -- layer=1 filter=40 channel=3
    -3, 0, -3, 9, -7, -4, 11, -9, 0,
    -- layer=1 filter=40 channel=4
    -1, -8, -4, -2, -2, -12, 6, -5, 6,
    -- layer=1 filter=40 channel=5
    -46, -53, -25, -17, -8, 18, 4, 22, 17,
    -- layer=1 filter=40 channel=6
    -17, -32, -17, -84, -67, -86, -13, -21, -35,
    -- layer=1 filter=40 channel=7
    -47, -79, -21, -29, -48, 11, -8, -5, 24,
    -- layer=1 filter=40 channel=8
    -49, -72, -28, 12, 8, 37, 13, 39, 31,
    -- layer=1 filter=40 channel=9
    -13, 14, -25, -3, -5, -21, 15, 18, -4,
    -- layer=1 filter=40 channel=10
    -44, -70, -12, -21, -36, 24, 26, -27, 28,
    -- layer=1 filter=40 channel=11
    -4, 1, -3, 7, 17, -7, 2, -14, -2,
    -- layer=1 filter=40 channel=12
    11, 9, 31, -38, 7, -12, -10, 26, 13,
    -- layer=1 filter=40 channel=13
    -22, -32, -39, -29, -32, -39, -13, -29, -51,
    -- layer=1 filter=40 channel=14
    -63, -49, -10, 25, 30, 5, 5, 7, 3,
    -- layer=1 filter=40 channel=15
    -43, -25, -34, -17, -11, -21, 7, 0, 7,
    -- layer=1 filter=40 channel=16
    -37, -70, -46, 25, 12, 43, 36, 33, 22,
    -- layer=1 filter=40 channel=17
    14, 10, 9, 8, -2, 0, -8, -17, -2,
    -- layer=1 filter=40 channel=18
    11, -6, 11, 34, 37, 29, 8, 6, 4,
    -- layer=1 filter=40 channel=19
    -17, -9, -45, 22, -13, -32, 9, 8, -11,
    -- layer=1 filter=40 channel=20
    -7, 3, -3, -29, -24, -34, -31, -19, -30,
    -- layer=1 filter=40 channel=21
    -51, -44, -22, -37, -41, -41, -6, -23, -12,
    -- layer=1 filter=40 channel=22
    -37, -38, -33, -20, -36, -47, 6, -22, -16,
    -- layer=1 filter=40 channel=23
    -12, -35, -41, -36, -12, -36, -15, -7, -13,
    -- layer=1 filter=40 channel=24
    -27, -31, -49, -28, -17, -10, 22, 20, 7,
    -- layer=1 filter=40 channel=25
    -67, -92, -45, -40, -67, 15, -1, -5, -2,
    -- layer=1 filter=40 channel=26
    0, -29, -52, -2, -11, -36, 21, 6, -10,
    -- layer=1 filter=40 channel=27
    -9, -2, -7, 0, 16, -2, -22, -2, -1,
    -- layer=1 filter=40 channel=28
    -39, -64, -7, -24, -60, 0, 11, -21, 34,
    -- layer=1 filter=40 channel=29
    -5, 6, -3, -26, -10, -15, -23, -17, -28,
    -- layer=1 filter=40 channel=30
    34, -10, 12, 32, 47, 17, 34, 12, 10,
    -- layer=1 filter=40 channel=31
    -16, -30, -8, -6, -3, -28, -23, -7, -27,
    -- layer=1 filter=40 channel=32
    27, -38, -26, -3, -1, -7, 23, -5, -16,
    -- layer=1 filter=40 channel=33
    -5, 0, 8, 4, 5, 6, 5, 14, -4,
    -- layer=1 filter=40 channel=34
    -3, -6, 8, -3, -8, -9, -17, -2, -13,
    -- layer=1 filter=40 channel=35
    -5, -6, -5, -9, -14, 0, -14, -8, -9,
    -- layer=1 filter=40 channel=36
    17, 19, 15, 22, 13, 11, 3, -1, 8,
    -- layer=1 filter=40 channel=37
    -29, -48, -35, 5, 8, 24, 14, 21, 13,
    -- layer=1 filter=40 channel=38
    -12, -3, -11, -28, -30, -40, -20, -39, -35,
    -- layer=1 filter=40 channel=39
    8, -5, 2, -3, 0, 0, 8, 8, 2,
    -- layer=1 filter=40 channel=40
    -40, -47, -47, -16, -16, -26, -7, -1, -18,
    -- layer=1 filter=40 channel=41
    65, -4, -38, 2, 14, 2, 48, 8, 12,
    -- layer=1 filter=40 channel=42
    8, 1, 41, -34, 22, 17, -51, -55, -26,
    -- layer=1 filter=40 channel=43
    -53, -95, -45, -15, -14, 19, 21, 14, 20,
    -- layer=1 filter=40 channel=44
    -16, -45, -43, 14, -13, -20, 43, -10, 0,
    -- layer=1 filter=40 channel=45
    -26, -20, -17, -19, 0, -13, 0, 13, -5,
    -- layer=1 filter=40 channel=46
    -31, -2, -18, 20, -7, -35, -26, 14, -20,
    -- layer=1 filter=40 channel=47
    -18, -39, -54, -21, -30, -44, -25, 4, -22,
    -- layer=1 filter=40 channel=48
    -19, -21, -17, -26, -6, -14, 0, -15, -6,
    -- layer=1 filter=40 channel=49
    -24, -17, -1, -26, -19, -13, -25, -26, -29,
    -- layer=1 filter=40 channel=50
    0, 0, -6, 3, -15, -11, -16, -14, -9,
    -- layer=1 filter=40 channel=51
    -22, -31, -27, -11, -42, -20, 2, -28, 16,
    -- layer=1 filter=40 channel=52
    10, 0, -14, 9, 2, 12, 16, 0, 20,
    -- layer=1 filter=40 channel=53
    3, 6, 11, -4, -16, 3, 0, 1, -18,
    -- layer=1 filter=40 channel=54
    -87, -60, -23, -26, -46, 14, 12, 3, 2,
    -- layer=1 filter=40 channel=55
    -20, -8, -26, -5, -8, -10, -12, -8, -16,
    -- layer=1 filter=40 channel=56
    0, -10, -2, -5, 4, 9, 0, 2, -1,
    -- layer=1 filter=40 channel=57
    -57, -107, -40, -31, -61, 0, 21, -31, 22,
    -- layer=1 filter=40 channel=58
    -72, -68, -65, -63, -49, -31, 5, -9, -27,
    -- layer=1 filter=40 channel=59
    -9, -1, -3, 0, -7, 3, 5, 2, -9,
    -- layer=1 filter=40 channel=60
    -7, -17, -17, -20, 1, -22, -13, -6, -7,
    -- layer=1 filter=40 channel=61
    -1, -3, -9, -5, 11, -2, 4, -6, -1,
    -- layer=1 filter=40 channel=62
    -59, -75, -32, 18, -7, 27, 23, 25, 16,
    -- layer=1 filter=40 channel=63
    11, -3, -1, 28, 21, 22, 0, 0, 8,
    -- layer=1 filter=40 channel=64
    0, 12, -4, 6, 4, 2, 0, 12, 3,
    -- layer=1 filter=40 channel=65
    -16, -10, 0, -6, -6, -24, -2, -25, -7,
    -- layer=1 filter=40 channel=66
    20, 9, 7, 9, 13, 9, -1, -7, 7,
    -- layer=1 filter=40 channel=67
    -6, -18, -27, -44, -36, -38, 19, -5, -11,
    -- layer=1 filter=40 channel=68
    1, -40, -57, -6, -15, -15, 49, -14, 3,
    -- layer=1 filter=40 channel=69
    -44, -59, -58, 4, 9, 11, 17, 37, 20,
    -- layer=1 filter=40 channel=70
    -30, -23, -23, -15, -44, -10, -17, 16, -41,
    -- layer=1 filter=40 channel=71
    -12, -14, -3, -13, -5, -3, 9, 25, 8,
    -- layer=1 filter=40 channel=72
    15, -15, -23, 24, 10, -30, 23, 10, 10,
    -- layer=1 filter=40 channel=73
    -12, -9, 6, -5, -8, -12, -3, -6, 4,
    -- layer=1 filter=40 channel=74
    0, -13, -21, -6, -5, 1, 33, -14, 3,
    -- layer=1 filter=40 channel=75
    0, -9, 13, 8, 27, -2, 6, 46, 36,
    -- layer=1 filter=40 channel=76
    33, 0, -3, 11, 25, 6, 23, -16, -13,
    -- layer=1 filter=40 channel=77
    -11, -10, 1, -7, -22, -18, -2, -9, -14,
    -- layer=1 filter=40 channel=78
    4, 2, 15, 2, 5, 18, 0, -9, 12,
    -- layer=1 filter=40 channel=79
    -55, -74, -29, 25, 1, 28, 10, 28, 18,
    -- layer=1 filter=40 channel=80
    3, 7, 6, -6, -2, -9, 2, -10, -8,
    -- layer=1 filter=40 channel=81
    -36, -36, -29, -10, -2, 4, 12, 15, 12,
    -- layer=1 filter=40 channel=82
    -43, -23, -12, -40, -25, -21, -9, -38, -26,
    -- layer=1 filter=40 channel=83
    -30, -27, -37, 0, -2, -15, 6, 2, -12,
    -- layer=1 filter=40 channel=84
    17, -11, -5, 12, 30, 23, 38, 0, -2,
    -- layer=1 filter=40 channel=85
    -41, -39, -59, -54, -52, -38, -8, -16, -39,
    -- layer=1 filter=40 channel=86
    17, 11, 10, 0, -10, -6, -6, -13, 2,
    -- layer=1 filter=40 channel=87
    13, 4, -38, 12, -7, -43, 1, 15, -42,
    -- layer=1 filter=40 channel=88
    -22, -3, 4, -36, -21, -13, -9, -19, -9,
    -- layer=1 filter=40 channel=89
    -33, -21, -31, -18, -11, -30, 0, -15, -22,
    -- layer=1 filter=40 channel=90
    -32, -52, -97, -8, -36, -38, 34, 1, -7,
    -- layer=1 filter=40 channel=91
    -1, -2, 5, -15, -13, -13, 0, -11, -11,
    -- layer=1 filter=40 channel=92
    1, -18, -85, -20, -7, -18, 49, -17, 13,
    -- layer=1 filter=40 channel=93
    -2, -7, -4, -11, -16, 8, -6, 10, -1,
    -- layer=1 filter=40 channel=94
    24, 24, 17, 22, 10, 28, -6, 8, 4,
    -- layer=1 filter=40 channel=95
    26, 2, 13, 41, 37, 28, 7, 3, 11,
    -- layer=1 filter=40 channel=96
    11, 4, 0, -8, 14, 12, 5, -2, 14,
    -- layer=1 filter=40 channel=97
    4, 6, 3, 13, -2, 6, 8, 0, 0,
    -- layer=1 filter=40 channel=98
    -44, -58, -17, 4, -5, 9, 12, 7, 13,
    -- layer=1 filter=40 channel=99
    -46, -74, -27, -19, -48, 9, 52, -48, 39,
    -- layer=1 filter=40 channel=100
    4, -3, 4, 11, 10, -2, -7, -28, -19,
    -- layer=1 filter=40 channel=101
    -9, -1, 12, -25, -26, -24, -15, -30, -24,
    -- layer=1 filter=40 channel=102
    34, 30, 40, 9, 19, 26, 10, 1, 0,
    -- layer=1 filter=40 channel=103
    5, 15, -2, 7, 21, -5, -19, -23, -14,
    -- layer=1 filter=40 channel=104
    -22, -10, -22, -8, 5, -20, -12, -11, -34,
    -- layer=1 filter=40 channel=105
    19, 5, 19, 9, 8, 19, -2, 5, 13,
    -- layer=1 filter=40 channel=106
    -28, -27, -13, -38, -20, -22, -18, -21, -29,
    -- layer=1 filter=40 channel=107
    -6, 1, 13, 0, -2, -2, 5, -5, 4,
    -- layer=1 filter=40 channel=108
    -13, -86, -76, -2, -32, -25, 7, -5, -14,
    -- layer=1 filter=40 channel=109
    -7, 0, 0, 3, 5, -4, -7, 6, -9,
    -- layer=1 filter=40 channel=110
    5, -4, 8, -6, -1, 12, -3, 1, -5,
    -- layer=1 filter=40 channel=111
    37, -7, 29, 24, 55, 56, 35, 4, 23,
    -- layer=1 filter=40 channel=112
    3, -9, 6, 33, 40, 40, 13, 13, 7,
    -- layer=1 filter=40 channel=113
    -48, -32, -23, -47, -47, -34, -42, -74, -51,
    -- layer=1 filter=40 channel=114
    -32, -48, -34, -11, 7, 13, 14, 27, 14,
    -- layer=1 filter=40 channel=115
    9, 11, 19, -9, -1, 20, -9, -14, 19,
    -- layer=1 filter=40 channel=116
    8, 6, -6, -10, -6, -11, 4, 8, 2,
    -- layer=1 filter=40 channel=117
    0, -23, 33, 4, 34, 29, 45, 11, 19,
    -- layer=1 filter=40 channel=118
    29, -2, 4, 29, 25, 33, 21, -10, 16,
    -- layer=1 filter=40 channel=119
    14, -42, -62, -3, -5, -23, 16, -9, -18,
    -- layer=1 filter=40 channel=120
    -27, -48, -24, -44, -51, -27, -23, -30, -16,
    -- layer=1 filter=40 channel=121
    -7, 0, -10, 25, 15, -10, -15, -6, -21,
    -- layer=1 filter=40 channel=122
    8, -9, -3, 2, -1, -5, 7, -5, -4,
    -- layer=1 filter=40 channel=123
    -3, 0, -7, 14, 19, 4, 0, -1, -6,
    -- layer=1 filter=40 channel=124
    -1, -4, -7, -13, -2, -17, -6, -3, 2,
    -- layer=1 filter=40 channel=125
    -37, -50, -24, -20, -8, -37, -26, -66, -40,
    -- layer=1 filter=40 channel=126
    -39, -48, -20, -25, -26, -9, 24, 12, 17,
    -- layer=1 filter=40 channel=127
    31, 1, 18, 30, 53, 24, 28, 12, 21,
    -- layer=1 filter=41 channel=0
    0, 6, -10, 0, -5, 1, -10, 0, 4,
    -- layer=1 filter=41 channel=1
    -10, 2, -7, -12, 8, 0, -6, -7, -7,
    -- layer=1 filter=41 channel=2
    0, 3, -10, 1, -3, -8, 4, 10, -7,
    -- layer=1 filter=41 channel=3
    0, 8, 0, 2, 9, 9, -9, 4, 3,
    -- layer=1 filter=41 channel=4
    2, 1, -1, 2, -6, -10, 4, 1, -12,
    -- layer=1 filter=41 channel=5
    -9, -3, -3, 3, -13, -12, -10, 2, -8,
    -- layer=1 filter=41 channel=6
    -2, -12, 2, -6, -11, -12, -8, 0, -9,
    -- layer=1 filter=41 channel=7
    -11, -6, -5, -5, -7, -11, -5, -7, -6,
    -- layer=1 filter=41 channel=8
    -1, -4, -1, -3, 5, -10, -9, -4, 8,
    -- layer=1 filter=41 channel=9
    -2, 1, -7, -2, 4, -9, 0, -10, 6,
    -- layer=1 filter=41 channel=10
    -4, -11, 2, -5, -15, -9, 3, -1, 0,
    -- layer=1 filter=41 channel=11
    -10, 5, -6, 4, -5, -3, 5, 1, -5,
    -- layer=1 filter=41 channel=12
    6, -3, -1, 7, -7, -6, -1, -3, 0,
    -- layer=1 filter=41 channel=13
    2, -14, 2, -8, -4, 0, -4, -5, 0,
    -- layer=1 filter=41 channel=14
    -4, 6, -2, -6, -3, 7, -9, 0, -10,
    -- layer=1 filter=41 channel=15
    4, -6, -2, -14, -8, 2, 8, 5, -2,
    -- layer=1 filter=41 channel=16
    3, 1, 10, -2, 0, -8, -2, 3, -10,
    -- layer=1 filter=41 channel=17
    3, -7, -1, -9, -10, -2, -5, -9, 4,
    -- layer=1 filter=41 channel=18
    -6, 6, -12, -3, -12, -2, 7, 1, 7,
    -- layer=1 filter=41 channel=19
    -2, -1, -2, -7, -2, -2, 0, -1, -2,
    -- layer=1 filter=41 channel=20
    1, 1, -2, 0, -4, -4, 3, -9, -8,
    -- layer=1 filter=41 channel=21
    6, -3, 2, -11, 4, 0, -4, -7, -9,
    -- layer=1 filter=41 channel=22
    1, -2, -5, -1, 3, 1, 8, -2, -1,
    -- layer=1 filter=41 channel=23
    9, -11, -3, 2, 8, -1, -11, 0, 8,
    -- layer=1 filter=41 channel=24
    4, -1, -11, -11, -7, -6, 0, -5, 0,
    -- layer=1 filter=41 channel=25
    2, -2, -6, 1, 0, -5, -12, -5, 2,
    -- layer=1 filter=41 channel=26
    -2, -7, -5, -9, 3, -15, 4, -3, -9,
    -- layer=1 filter=41 channel=27
    -6, -3, 1, 3, 0, 4, -6, 7, 11,
    -- layer=1 filter=41 channel=28
    5, -10, 12, -11, -7, -3, 4, 7, 6,
    -- layer=1 filter=41 channel=29
    2, 4, 9, 6, 4, 7, 4, 1, -2,
    -- layer=1 filter=41 channel=30
    1, 1, -2, 2, -13, 1, 1, 0, -2,
    -- layer=1 filter=41 channel=31
    -4, -4, -13, -2, 0, -12, 2, -12, -14,
    -- layer=1 filter=41 channel=32
    4, -2, -10, 3, -3, -3, -3, 5, -4,
    -- layer=1 filter=41 channel=33
    -8, -7, 2, 8, -3, 6, 0, 9, -4,
    -- layer=1 filter=41 channel=34
    -1, -10, -12, -4, -6, 0, -11, -4, 0,
    -- layer=1 filter=41 channel=35
    2, -5, 2, 7, 7, -1, 0, -7, 6,
    -- layer=1 filter=41 channel=36
    -9, 7, -11, 0, 0, -11, 4, -4, 0,
    -- layer=1 filter=41 channel=37
    -10, 7, 10, 2, -3, -7, 4, 7, 6,
    -- layer=1 filter=41 channel=38
    -2, -1, 1, -10, -1, -8, -8, -3, -8,
    -- layer=1 filter=41 channel=39
    2, -9, -10, 0, 5, -9, 6, 2, -10,
    -- layer=1 filter=41 channel=40
    -11, -4, 1, -13, -17, -10, 6, -20, -4,
    -- layer=1 filter=41 channel=41
    10, 1, 0, 1, -11, -2, -3, 3, 1,
    -- layer=1 filter=41 channel=42
    -9, 6, -4, -5, 6, -2, -3, 1, 1,
    -- layer=1 filter=41 channel=43
    -5, -2, 0, 0, -12, 1, 7, 0, -7,
    -- layer=1 filter=41 channel=44
    6, 7, -6, 6, 0, -2, -4, -9, -6,
    -- layer=1 filter=41 channel=45
    -1, -1, -7, -8, 0, -8, -7, 7, 1,
    -- layer=1 filter=41 channel=46
    -3, -9, 2, -9, 10, 6, 2, 4, -6,
    -- layer=1 filter=41 channel=47
    -10, -8, -2, 3, 0, 7, 11, -2, 3,
    -- layer=1 filter=41 channel=48
    -4, 1, -9, 2, 4, 2, 6, 2, 5,
    -- layer=1 filter=41 channel=49
    5, -9, 4, 2, -8, -3, 6, 2, -6,
    -- layer=1 filter=41 channel=50
    -3, -5, -4, 3, 7, -7, -11, 6, 5,
    -- layer=1 filter=41 channel=51
    -3, 7, -10, -11, -8, -11, 3, -1, 5,
    -- layer=1 filter=41 channel=52
    -4, 0, -6, 0, 5, 6, 1, -4, -1,
    -- layer=1 filter=41 channel=53
    -5, 0, 2, -4, 0, -8, -5, 8, 5,
    -- layer=1 filter=41 channel=54
    1, 7, 8, -6, -10, -8, -11, -10, 3,
    -- layer=1 filter=41 channel=55
    -5, 2, 0, -16, 5, -6, -7, 10, -5,
    -- layer=1 filter=41 channel=56
    7, 0, -8, 8, 1, -9, 0, 8, 5,
    -- layer=1 filter=41 channel=57
    -1, 4, -11, 4, -6, -8, 1, -6, -8,
    -- layer=1 filter=41 channel=58
    5, -2, 7, -12, -4, 5, 5, -3, -8,
    -- layer=1 filter=41 channel=59
    8, -6, 0, 7, 3, 7, -4, -11, -11,
    -- layer=1 filter=41 channel=60
    -5, 7, -7, 5, -9, -7, -10, 7, -2,
    -- layer=1 filter=41 channel=61
    2, -7, 0, 9, -3, -5, 1, -7, 7,
    -- layer=1 filter=41 channel=62
    -3, 6, -10, 6, -8, 0, 0, -3, -2,
    -- layer=1 filter=41 channel=63
    -2, -12, 7, 3, 1, 4, 5, -9, -5,
    -- layer=1 filter=41 channel=64
    2, 2, 0, 0, 6, -10, -2, -9, -3,
    -- layer=1 filter=41 channel=65
    7, -9, -2, -1, -2, 3, 6, 5, -4,
    -- layer=1 filter=41 channel=66
    -7, 0, 6, 6, 0, 8, -13, -11, -7,
    -- layer=1 filter=41 channel=67
    -1, 0, 7, -1, -3, -2, -5, -1, -1,
    -- layer=1 filter=41 channel=68
    -3, 5, -4, 5, 3, -8, -9, 9, -13,
    -- layer=1 filter=41 channel=69
    9, -4, -7, 3, -11, -14, -4, 6, -13,
    -- layer=1 filter=41 channel=70
    -7, 0, 4, -8, -10, -4, 5, 6, -10,
    -- layer=1 filter=41 channel=71
    -9, -3, 10, -4, -5, -2, -10, -2, 2,
    -- layer=1 filter=41 channel=72
    4, 5, 9, -11, 4, 1, -8, 2, -1,
    -- layer=1 filter=41 channel=73
    10, -8, -5, -10, -5, 3, 0, 2, 7,
    -- layer=1 filter=41 channel=74
    0, 7, -8, 4, 5, 4, -8, 7, -4,
    -- layer=1 filter=41 channel=75
    -7, 3, 2, 3, 1, 0, -10, -12, 0,
    -- layer=1 filter=41 channel=76
    9, -2, 1, -1, -4, -5, -11, -9, -4,
    -- layer=1 filter=41 channel=77
    -4, -9, 3, -2, -2, -7, -7, -3, 0,
    -- layer=1 filter=41 channel=78
    -6, -10, 3, -1, -8, 1, 2, 3, 0,
    -- layer=1 filter=41 channel=79
    -9, -10, -11, -5, -5, 0, 0, -13, -15,
    -- layer=1 filter=41 channel=80
    2, -9, 3, 0, -6, -6, -6, -5, -7,
    -- layer=1 filter=41 channel=81
    0, 6, 1, -14, -6, 2, -6, 2, 0,
    -- layer=1 filter=41 channel=82
    5, -6, -6, 4, -1, -9, 12, -10, 0,
    -- layer=1 filter=41 channel=83
    -11, -5, 0, 8, 4, -13, -4, -2, 4,
    -- layer=1 filter=41 channel=84
    8, 3, -7, -10, 0, 1, 9, -6, 4,
    -- layer=1 filter=41 channel=85
    8, -4, 0, 0, -11, 0, 4, -5, 5,
    -- layer=1 filter=41 channel=86
    -9, 0, -7, -4, -9, -4, -12, -2, -7,
    -- layer=1 filter=41 channel=87
    0, -6, -8, -10, 7, -9, 5, 3, -1,
    -- layer=1 filter=41 channel=88
    6, 2, 9, 0, -4, 1, 0, -1, -10,
    -- layer=1 filter=41 channel=89
    4, -8, -10, -2, -11, 1, -11, -3, -1,
    -- layer=1 filter=41 channel=90
    4, -2, 1, 0, -2, -11, 0, 2, 1,
    -- layer=1 filter=41 channel=91
    5, -3, -1, -13, -15, 2, -3, -7, -12,
    -- layer=1 filter=41 channel=92
    -3, 8, 3, -9, 0, 2, -9, -3, -7,
    -- layer=1 filter=41 channel=93
    -14, 6, -12, -7, -11, -3, -8, 8, -8,
    -- layer=1 filter=41 channel=94
    -1, 8, -3, 0, 7, 4, -4, 7, -1,
    -- layer=1 filter=41 channel=95
    -7, 2, -3, -5, 3, 7, 0, 6, -9,
    -- layer=1 filter=41 channel=96
    -8, -7, -8, 4, 1, 1, -1, -12, -2,
    -- layer=1 filter=41 channel=97
    4, -5, 8, -7, -10, -7, -4, 0, -4,
    -- layer=1 filter=41 channel=98
    -5, -3, 3, -4, -7, -4, -10, -6, -11,
    -- layer=1 filter=41 channel=99
    -6, -8, -3, -13, 5, -6, -9, -4, -6,
    -- layer=1 filter=41 channel=100
    -3, -6, -3, -4, -10, -5, 0, -2, 6,
    -- layer=1 filter=41 channel=101
    -3, 7, -7, 2, -7, 5, 0, -4, 0,
    -- layer=1 filter=41 channel=102
    3, -1, -4, -1, -11, -1, 1, 4, -10,
    -- layer=1 filter=41 channel=103
    -9, 8, -2, -7, 2, 7, -7, -1, -7,
    -- layer=1 filter=41 channel=104
    -8, 0, 6, 2, -2, -5, -7, 7, -6,
    -- layer=1 filter=41 channel=105
    7, 0, 6, -11, 7, 2, -10, -10, -3,
    -- layer=1 filter=41 channel=106
    0, -5, 0, -10, -10, 1, 1, -4, 1,
    -- layer=1 filter=41 channel=107
    8, 4, -10, -1, 7, -2, 8, 8, -7,
    -- layer=1 filter=41 channel=108
    -10, -11, 1, -3, -11, -5, 0, -7, 1,
    -- layer=1 filter=41 channel=109
    0, 6, -10, -11, 10, 2, -5, 3, -9,
    -- layer=1 filter=41 channel=110
    -7, -6, 0, 1, 0, -9, 1, -5, -6,
    -- layer=1 filter=41 channel=111
    -10, 5, -2, 5, 5, 3, -7, 2, 5,
    -- layer=1 filter=41 channel=112
    -7, -9, 2, -4, 3, 0, -1, 3, -6,
    -- layer=1 filter=41 channel=113
    7, -15, 6, -2, -6, -8, -6, -8, -10,
    -- layer=1 filter=41 channel=114
    -1, -9, -8, 0, -8, 8, -1, 7, 2,
    -- layer=1 filter=41 channel=115
    -11, -2, -5, 6, -9, -2, -2, -9, 3,
    -- layer=1 filter=41 channel=116
    -8, -5, -7, 4, 5, -3, -10, -3, -9,
    -- layer=1 filter=41 channel=117
    1, 3, -6, -2, -2, 0, 1, 7, -6,
    -- layer=1 filter=41 channel=118
    -7, 4, 1, -2, -4, -4, -10, 1, 2,
    -- layer=1 filter=41 channel=119
    -3, 2, -11, 9, -3, 3, 0, -10, -5,
    -- layer=1 filter=41 channel=120
    -3, 8, 2, -13, -8, -11, -3, 4, 0,
    -- layer=1 filter=41 channel=121
    -4, 9, 4, -3, 2, 4, 2, 1, -4,
    -- layer=1 filter=41 channel=122
    10, -10, 5, -4, -10, -5, 7, -4, 9,
    -- layer=1 filter=41 channel=123
    1, 8, -5, -8, -6, 3, -11, -3, -11,
    -- layer=1 filter=41 channel=124
    -9, 0, 1, -5, -6, -10, 0, 5, -10,
    -- layer=1 filter=41 channel=125
    -12, -11, -2, -6, -7, -11, -8, -11, 1,
    -- layer=1 filter=41 channel=126
    -4, 0, -11, -7, -8, -4, -7, 6, 5,
    -- layer=1 filter=41 channel=127
    -7, -14, -2, 4, 5, -6, -3, -4, 9,
    -- layer=1 filter=42 channel=0
    7, -7, 4, 12, 3, 6, 16, 7, -3,
    -- layer=1 filter=42 channel=1
    2, -5, -5, 9, 4, 1, 16, -13, 12,
    -- layer=1 filter=42 channel=2
    6, 3, 6, 9, 4, 20, -9, -23, 0,
    -- layer=1 filter=42 channel=3
    -8, 0, -6, -10, 1, 4, -14, 4, -15,
    -- layer=1 filter=42 channel=4
    4, 5, 4, -4, 1, -10, 1, 7, -1,
    -- layer=1 filter=42 channel=5
    -8, -5, 4, 18, -17, -12, 11, -19, 13,
    -- layer=1 filter=42 channel=6
    -5, -12, -3, -15, -4, -6, -9, -3, -3,
    -- layer=1 filter=42 channel=7
    -14, -23, 14, -16, 14, 21, -3, 0, 0,
    -- layer=1 filter=42 channel=8
    -5, -8, -12, 20, 9, -7, 17, -2, 18,
    -- layer=1 filter=42 channel=9
    8, 8, 4, 3, 19, -21, 8, -9, 16,
    -- layer=1 filter=42 channel=10
    -17, -7, 5, -15, 9, 7, -8, -1, -9,
    -- layer=1 filter=42 channel=11
    -21, -31, -33, -15, -31, -24, 3, -25, -29,
    -- layer=1 filter=42 channel=12
    29, -15, -14, -15, -53, -52, 21, -3, 12,
    -- layer=1 filter=42 channel=13
    -10, -4, -15, 9, 0, 2, 3, 8, -4,
    -- layer=1 filter=42 channel=14
    -15, 10, -8, -11, -19, -1, 5, -16, -21,
    -- layer=1 filter=42 channel=15
    -2, -10, -5, 29, -10, 4, 16, -22, -17,
    -- layer=1 filter=42 channel=16
    4, -3, 1, 2, -8, -10, -10, -8, 5,
    -- layer=1 filter=42 channel=17
    8, -7, -15, 10, -10, -4, 0, 1, -1,
    -- layer=1 filter=42 channel=18
    -31, -30, -44, -4, -14, -12, -16, -20, -9,
    -- layer=1 filter=42 channel=19
    -9, -24, 14, 21, -2, -8, -6, 37, 23,
    -- layer=1 filter=42 channel=20
    -3, -4, 8, 10, 14, -2, 9, 0, 2,
    -- layer=1 filter=42 channel=21
    4, -2, -10, 0, 9, -4, -2, -8, 3,
    -- layer=1 filter=42 channel=22
    0, -17, -11, 3, -13, 3, 5, -1, 10,
    -- layer=1 filter=42 channel=23
    16, -19, 11, 6, -5, -7, 0, 22, -29,
    -- layer=1 filter=42 channel=24
    -3, 14, 0, 4, -1, 1, -8, 1, 10,
    -- layer=1 filter=42 channel=25
    -20, -29, -1, 0, 5, 0, -21, 9, 9,
    -- layer=1 filter=42 channel=26
    -6, -6, -8, 4, -11, 5, 2, 0, -10,
    -- layer=1 filter=42 channel=27
    26, 24, 28, 8, 3, 22, -2, -14, -8,
    -- layer=1 filter=42 channel=28
    -20, -19, 7, -16, 8, 15, -3, 11, 16,
    -- layer=1 filter=42 channel=29
    9, 5, 7, 9, 12, 10, -15, 5, 0,
    -- layer=1 filter=42 channel=30
    -16, -23, -28, 17, 3, -16, 17, -1, 11,
    -- layer=1 filter=42 channel=31
    -27, -10, -22, -15, -26, -37, -21, -10, -6,
    -- layer=1 filter=42 channel=32
    -7, -7, 1, 7, 7, 6, 7, 17, 7,
    -- layer=1 filter=42 channel=33
    -9, 4, -14, -5, 9, -10, 6, -2, -8,
    -- layer=1 filter=42 channel=34
    -6, 2, 17, -6, 2, 15, -4, 1, 0,
    -- layer=1 filter=42 channel=35
    3, 6, 0, 7, 19, 3, 6, 3, 15,
    -- layer=1 filter=42 channel=36
    -41, -38, -41, -31, -30, -25, -30, -33, -30,
    -- layer=1 filter=42 channel=37
    -15, -14, -6, -4, -15, -19, 2, -3, -2,
    -- layer=1 filter=42 channel=38
    -1, -2, -14, 14, 0, 0, 3, 1, 10,
    -- layer=1 filter=42 channel=39
    -5, -5, -8, 9, -19, -10, 0, 9, -9,
    -- layer=1 filter=42 channel=40
    -15, -12, -12, -4, -6, -20, -7, -11, -6,
    -- layer=1 filter=42 channel=41
    14, 10, 31, 0, 17, -25, -7, -15, 24,
    -- layer=1 filter=42 channel=42
    -2, 0, -4, -5, -14, -5, -6, -13, -27,
    -- layer=1 filter=42 channel=43
    -3, -12, 3, 18, 7, 20, 12, -12, 10,
    -- layer=1 filter=42 channel=44
    -6, -2, 4, 10, 4, 4, 27, 16, 1,
    -- layer=1 filter=42 channel=45
    -8, 1, -10, 3, 8, -4, 20, -2, 2,
    -- layer=1 filter=42 channel=46
    -25, -28, 15, 0, -25, -32, -15, 13, 18,
    -- layer=1 filter=42 channel=47
    7, -9, 25, 2, 15, 0, -22, 18, -5,
    -- layer=1 filter=42 channel=48
    -9, 0, -3, 1, 1, -3, 0, 2, 10,
    -- layer=1 filter=42 channel=49
    -3, -2, -1, 4, 3, 1, -3, 1, -9,
    -- layer=1 filter=42 channel=50
    -11, 14, -6, -2, -8, 4, -3, 3, 5,
    -- layer=1 filter=42 channel=51
    -6, -11, 6, -1, -2, 2, 7, 8, -10,
    -- layer=1 filter=42 channel=52
    5, 12, 9, -3, -2, 4, -6, 4, 8,
    -- layer=1 filter=42 channel=53
    -3, 5, -1, 5, 1, -2, 0, -4, -10,
    -- layer=1 filter=42 channel=54
    0, -16, 16, 1, -2, 1, -23, 12, 0,
    -- layer=1 filter=42 channel=55
    -5, -7, -4, -24, -35, -15, -26, -17, -28,
    -- layer=1 filter=42 channel=56
    8, 1, -6, 1, 1, -3, 2, -4, 0,
    -- layer=1 filter=42 channel=57
    -23, -23, 1, -26, 1, 0, -11, -2, -13,
    -- layer=1 filter=42 channel=58
    -6, 5, 13, 8, 22, 3, -26, 46, -20,
    -- layer=1 filter=42 channel=59
    -2, -2, 17, 1, 1, 14, 9, 1, 14,
    -- layer=1 filter=42 channel=60
    5, 8, 0, -13, 5, 6, 13, 1, -5,
    -- layer=1 filter=42 channel=61
    6, -17, -6, -17, 0, 0, -12, 2, -2,
    -- layer=1 filter=42 channel=62
    -3, -5, -14, 24, -14, -11, 6, -4, 7,
    -- layer=1 filter=42 channel=63
    -10, -22, -2, -8, -4, -5, 10, -15, 2,
    -- layer=1 filter=42 channel=64
    0, -6, 5, -7, -4, 0, -4, 13, 16,
    -- layer=1 filter=42 channel=65
    14, -1, 4, 5, -3, 4, 14, -5, 2,
    -- layer=1 filter=42 channel=66
    -4, 6, 5, 6, 2, 2, -4, 1, -9,
    -- layer=1 filter=42 channel=67
    -27, -27, -20, -23, -32, -24, -61, -60, -43,
    -- layer=1 filter=42 channel=68
    -9, 1, -13, -8, 16, 8, 31, 4, 14,
    -- layer=1 filter=42 channel=69
    -9, 12, 0, 15, -18, -2, 1, -14, 1,
    -- layer=1 filter=42 channel=70
    -19, -33, -3, -29, -35, -26, -39, -30, -22,
    -- layer=1 filter=42 channel=71
    0, -6, 7, 7, -11, 8, -11, -13, 0,
    -- layer=1 filter=42 channel=72
    -6, -13, -22, 11, -12, -16, -3, -7, 11,
    -- layer=1 filter=42 channel=73
    5, 1, 3, -9, 6, 4, -3, 3, -5,
    -- layer=1 filter=42 channel=74
    -8, 3, -1, 2, 8, -4, 22, -9, 0,
    -- layer=1 filter=42 channel=75
    -15, -29, -10, 2, -12, -16, 0, 6, -34,
    -- layer=1 filter=42 channel=76
    -7, -8, -12, 16, 24, -11, 16, 6, 9,
    -- layer=1 filter=42 channel=77
    3, 5, 0, 3, 9, 5, 8, -9, -4,
    -- layer=1 filter=42 channel=78
    -8, 3, 5, -1, 11, 0, 6, 4, 12,
    -- layer=1 filter=42 channel=79
    2, 5, -8, 9, 6, 5, 7, -3, 11,
    -- layer=1 filter=42 channel=80
    -4, -5, -3, 5, -4, -8, -2, 5, 5,
    -- layer=1 filter=42 channel=81
    5, 17, 16, 2, 2, 6, -10, -6, 7,
    -- layer=1 filter=42 channel=82
    12, 5, -4, -1, 7, 11, 3, -1, 15,
    -- layer=1 filter=42 channel=83
    1, -4, -14, 22, 0, 12, 14, 10, 0,
    -- layer=1 filter=42 channel=84
    -18, 0, -20, 8, 16, -8, 16, -12, 5,
    -- layer=1 filter=42 channel=85
    -4, 0, 27, 3, 5, 0, -17, 17, -6,
    -- layer=1 filter=42 channel=86
    -20, -23, -6, -9, -19, -23, -20, -21, -2,
    -- layer=1 filter=42 channel=87
    -3, -13, 10, -4, -2, -26, -9, -3, -4,
    -- layer=1 filter=42 channel=88
    2, 5, -6, -12, -4, -11, 0, -10, -5,
    -- layer=1 filter=42 channel=89
    3, 12, 11, 7, 2, -7, 6, 0, 12,
    -- layer=1 filter=42 channel=90
    -8, 0, -21, 2, 9, 3, 10, 14, -8,
    -- layer=1 filter=42 channel=91
    8, -5, 11, 3, 6, 6, 3, 4, 7,
    -- layer=1 filter=42 channel=92
    -2, -8, 0, -13, 10, -7, -4, -9, 4,
    -- layer=1 filter=42 channel=93
    14, 18, 9, -1, -1, 13, 7, 15, 4,
    -- layer=1 filter=42 channel=94
    -6, -8, -11, 0, 5, -7, 1, -3, 6,
    -- layer=1 filter=42 channel=95
    -4, -21, -10, 8, 14, -15, 14, 9, 8,
    -- layer=1 filter=42 channel=96
    -13, 6, -1, 4, -1, -4, -12, -5, 0,
    -- layer=1 filter=42 channel=97
    7, -2, -9, 13, -7, 0, 13, 7, 0,
    -- layer=1 filter=42 channel=98
    4, -2, -24, 12, -6, -3, 15, 3, 7,
    -- layer=1 filter=42 channel=99
    -7, 6, -20, 2, 13, 12, 30, 3, 22,
    -- layer=1 filter=42 channel=100
    -19, -29, -26, -15, 0, -33, 9, -17, -1,
    -- layer=1 filter=42 channel=101
    -4, 0, 10, 15, 13, 9, 18, 1, 9,
    -- layer=1 filter=42 channel=102
    16, 9, -7, 22, 3, 1, 21, 17, 4,
    -- layer=1 filter=42 channel=103
    -14, -12, -19, -5, -11, -21, -12, -7, -18,
    -- layer=1 filter=42 channel=104
    17, -27, 10, 7, -17, -13, 9, 2, -13,
    -- layer=1 filter=42 channel=105
    8, 6, -4, 6, 11, 4, 0, -2, -2,
    -- layer=1 filter=42 channel=106
    4, 11, -13, -1, 1, 3, 4, 17, 9,
    -- layer=1 filter=42 channel=107
    -7, 0, -4, -8, -1, 4, 2, -9, 0,
    -- layer=1 filter=42 channel=108
    8, 3, 0, -3, 6, 15, -1, 6, 3,
    -- layer=1 filter=42 channel=109
    7, -7, -4, -8, -13, -9, 1, 5, 3,
    -- layer=1 filter=42 channel=110
    -6, 0, 2, -7, 2, -7, 0, -6, 10,
    -- layer=1 filter=42 channel=111
    -17, -4, -22, 16, -2, -6, 17, 13, 14,
    -- layer=1 filter=42 channel=112
    -3, -8, -24, 9, 1, 5, 26, 0, -10,
    -- layer=1 filter=42 channel=113
    -19, -6, 1, -3, 13, 6, -11, -2, -4,
    -- layer=1 filter=42 channel=114
    -26, -18, -19, -12, -31, -52, -39, -46, -14,
    -- layer=1 filter=42 channel=115
    -15, -29, -2, -9, -18, -10, -18, -16, -5,
    -- layer=1 filter=42 channel=116
    -10, -5, 0, -6, 3, -7, 8, 6, -6,
    -- layer=1 filter=42 channel=117
    -2, -10, -33, -13, -11, -4, 28, 6, -14,
    -- layer=1 filter=42 channel=118
    -15, -3, -26, 8, 13, -9, 19, -5, 12,
    -- layer=1 filter=42 channel=119
    8, 16, 13, 6, 6, 15, 6, 24, 0,
    -- layer=1 filter=42 channel=120
    -4, 5, -1, 0, -5, -1, -4, 0, 7,
    -- layer=1 filter=42 channel=121
    -17, -24, -15, 2, -21, -9, 4, 1, -9,
    -- layer=1 filter=42 channel=122
    9, -10, -4, 2, -1, -2, -1, 3, -3,
    -- layer=1 filter=42 channel=123
    -20, -18, -3, -9, -23, -26, -4, 0, -11,
    -- layer=1 filter=42 channel=124
    5, 1, -1, 2, -10, 1, -4, 0, -11,
    -- layer=1 filter=42 channel=125
    -11, -25, -2, -16, -20, -18, -23, -6, -22,
    -- layer=1 filter=42 channel=126
    17, 4, -3, 5, -17, 24, 30, 16, 1,
    -- layer=1 filter=42 channel=127
    -17, -21, -27, 9, -1, -7, 19, -12, 15,
    -- layer=1 filter=43 channel=0
    6, 1, -1, 8, -9, -12, 22, 20, 5,
    -- layer=1 filter=43 channel=1
    -11, 41, 38, 26, 0, 32, 6, -2, 22,
    -- layer=1 filter=43 channel=2
    33, 30, 45, 22, 27, 11, 17, 26, 24,
    -- layer=1 filter=43 channel=3
    -5, -3, 9, 7, 4, 4, -1, 6, -1,
    -- layer=1 filter=43 channel=4
    -10, -1, 10, -2, -9, -4, -1, -5, 0,
    -- layer=1 filter=43 channel=5
    -19, 42, 47, 20, 0, 50, 31, 10, 17,
    -- layer=1 filter=43 channel=6
    -11, -4, 0, 4, 2, 31, -3, -41, -46,
    -- layer=1 filter=43 channel=7
    -35, -74, -13, -42, -175, -57, -45, -115, -51,
    -- layer=1 filter=43 channel=8
    8, 65, 41, 42, 17, 26, 17, 2, 25,
    -- layer=1 filter=43 channel=9
    -3, -7, 24, 1, 1, 23, 19, -7, -2,
    -- layer=1 filter=43 channel=10
    -17, -63, -20, -47, -154, -28, -34, -96, -38,
    -- layer=1 filter=43 channel=11
    -2, -9, -20, -9, -3, -2, 18, 7, -7,
    -- layer=1 filter=43 channel=12
    1, 31, 22, 21, 43, 12, 2, -9, 9,
    -- layer=1 filter=43 channel=13
    -4, 43, 5, -25, 14, -10, -7, -25, -9,
    -- layer=1 filter=43 channel=14
    -13, 0, -3, -44, -61, -63, -41, -39, -34,
    -- layer=1 filter=43 channel=15
    -19, 60, 79, 0, -1, 52, 38, -36, -16,
    -- layer=1 filter=43 channel=16
    -4, 42, 43, 26, 12, 36, 15, 13, 22,
    -- layer=1 filter=43 channel=17
    25, 8, 0, 11, 12, 5, 31, 27, 20,
    -- layer=1 filter=43 channel=18
    -44, -46, -27, -62, -48, -55, -31, -51, -34,
    -- layer=1 filter=43 channel=19
    -36, -32, -14, -37, -10, -2, -5, -39, -46,
    -- layer=1 filter=43 channel=20
    11, 22, 7, 5, 8, 11, 17, 0, 9,
    -- layer=1 filter=43 channel=21
    -25, -18, -19, -6, -31, -28, -14, -20, -6,
    -- layer=1 filter=43 channel=22
    -2, 45, 21, 17, -23, -9, 7, -8, 7,
    -- layer=1 filter=43 channel=23
    -10, -12, 8, 20, -15, 12, -5, -3, 6,
    -- layer=1 filter=43 channel=24
    0, 31, 14, -12, 14, 14, 10, -17, 21,
    -- layer=1 filter=43 channel=25
    -10, -31, -5, -1, -70, 14, -17, -18, -3,
    -- layer=1 filter=43 channel=26
    5, 64, 3, -7, 14, 6, 8, -7, 4,
    -- layer=1 filter=43 channel=27
    -9, -28, -42, -31, -34, -32, -16, -29, -35,
    -- layer=1 filter=43 channel=28
    -4, -44, -17, -27, -109, -69, -25, -72, -27,
    -- layer=1 filter=43 channel=29
    -12, -16, -41, -31, -24, -27, -22, -25, -26,
    -- layer=1 filter=43 channel=30
    -82, -59, -37, -78, -73, -80, -26, -75, -72,
    -- layer=1 filter=43 channel=31
    -18, -21, -17, -40, -43, -65, -72, -49, -64,
    -- layer=1 filter=43 channel=32
    -31, 30, -19, -44, -46, -12, 20, -87, -27,
    -- layer=1 filter=43 channel=33
    -9, 2, 10, -6, -9, 1, 1, -5, -5,
    -- layer=1 filter=43 channel=34
    15, 25, 30, 19, 0, 34, 0, -10, -8,
    -- layer=1 filter=43 channel=35
    -12, -8, -2, -5, -11, -11, 0, 2, 2,
    -- layer=1 filter=43 channel=36
    18, -1, -4, 17, 19, 1, 25, 28, 10,
    -- layer=1 filter=43 channel=37
    -12, 48, 35, 11, 18, 40, 15, 4, 17,
    -- layer=1 filter=43 channel=38
    -1, 2, -10, 0, 0, 0, -7, -14, -19,
    -- layer=1 filter=43 channel=39
    -3, -4, -16, 11, 15, 2, 15, 16, 12,
    -- layer=1 filter=43 channel=40
    -67, -53, -21, -58, -76, -97, -38, -95, -82,
    -- layer=1 filter=43 channel=41
    -16, 29, 3, 3, -43, -49, 27, -7, 7,
    -- layer=1 filter=43 channel=42
    54, 52, 32, 1, 38, 29, 6, 29, 24,
    -- layer=1 filter=43 channel=43
    -12, 28, 25, 24, -30, 12, -7, -5, 32,
    -- layer=1 filter=43 channel=44
    -11, 58, -20, -28, -12, -2, 23, -85, -20,
    -- layer=1 filter=43 channel=45
    -32, 41, 4, -30, 20, 9, -9, -36, -25,
    -- layer=1 filter=43 channel=46
    1, 20, 59, -14, 1, 43, 0, -1, -20,
    -- layer=1 filter=43 channel=47
    -36, -20, -3, 17, -52, -1, -16, -35, -5,
    -- layer=1 filter=43 channel=48
    -24, -34, -35, -13, -22, -14, -19, -19, -26,
    -- layer=1 filter=43 channel=49
    26, 7, 11, 19, 17, 6, -9, 6, -5,
    -- layer=1 filter=43 channel=50
    13, 7, 25, 3, -4, 0, 15, 13, -3,
    -- layer=1 filter=43 channel=51
    4, -37, -13, -22, -48, -33, -2, -48, -20,
    -- layer=1 filter=43 channel=52
    5, 10, 9, 17, 5, 11, 9, -4, 1,
    -- layer=1 filter=43 channel=53
    5, -1, 9, 9, 7, 0, 3, 4, -2,
    -- layer=1 filter=43 channel=54
    -9, -21, -12, -20, -38, 42, -12, -7, -11,
    -- layer=1 filter=43 channel=55
    9, 6, 16, 20, 13, 21, 9, 22, 12,
    -- layer=1 filter=43 channel=56
    -8, 9, -8, 2, 0, 0, 5, -3, 0,
    -- layer=1 filter=43 channel=57
    4, -44, -13, -38, -103, -35, -28, -91, -54,
    -- layer=1 filter=43 channel=58
    -44, -78, 0, -43, -92, 16, -73, -32, -48,
    -- layer=1 filter=43 channel=59
    -4, 2, -5, -5, -4, 0, 5, -9, -2,
    -- layer=1 filter=43 channel=60
    -4, -10, -16, 0, -8, -7, 0, -19, -5,
    -- layer=1 filter=43 channel=61
    -1, 1, 4, 7, -3, 0, -8, 0, -1,
    -- layer=1 filter=43 channel=62
    -18, 49, 27, 9, 6, 40, -5, 1, 39,
    -- layer=1 filter=43 channel=63
    6, -4, -10, -5, 0, -16, 19, 7, 7,
    -- layer=1 filter=43 channel=64
    -13, 1, 0, 0, -7, -9, -7, -7, 2,
    -- layer=1 filter=43 channel=65
    -14, -38, -40, -14, -23, -26, -29, -13, -26,
    -- layer=1 filter=43 channel=66
    8, -8, -15, 12, 0, -3, 24, 7, 10,
    -- layer=1 filter=43 channel=67
    -30, -31, -43, -55, -13, 0, -25, -29, -15,
    -- layer=1 filter=43 channel=68
    -19, 32, -51, -66, -31, -31, -2, -94, -17,
    -- layer=1 filter=43 channel=69
    -19, 64, 52, 23, 29, 44, 43, -16, -2,
    -- layer=1 filter=43 channel=70
    26, 47, 3, -37, -10, 11, -32, -26, -6,
    -- layer=1 filter=43 channel=71
    -13, -2, -3, -13, -23, 0, -7, 4, -14,
    -- layer=1 filter=43 channel=72
    -35, -24, -5, -21, -44, -22, -9, -11, -8,
    -- layer=1 filter=43 channel=73
    0, -7, 1, -7, 9, -10, 6, 10, -5,
    -- layer=1 filter=43 channel=74
    -40, 38, 0, -36, -11, -47, -20, -40, -34,
    -- layer=1 filter=43 channel=75
    -45, 3, -7, 7, -21, -72, -47, -34, 2,
    -- layer=1 filter=43 channel=76
    8, 8, -20, 6, -7, -7, 17, 1, -4,
    -- layer=1 filter=43 channel=77
    -28, -26, -37, -36, -22, -25, -16, -17, -10,
    -- layer=1 filter=43 channel=78
    11, 6, 0, 9, -14, 2, 6, 2, -7,
    -- layer=1 filter=43 channel=79
    0, 32, 50, 27, 16, 33, 22, 4, 31,
    -- layer=1 filter=43 channel=80
    9, -6, 0, -8, 8, 8, 7, 0, 3,
    -- layer=1 filter=43 channel=81
    -3, -16, -14, -16, -2, -8, -3, -5, 6,
    -- layer=1 filter=43 channel=82
    -31, -9, -11, -17, -14, -10, -27, -25, -19,
    -- layer=1 filter=43 channel=83
    -20, 44, 33, -13, 8, 1, 3, -19, 18,
    -- layer=1 filter=43 channel=84
    -78, -35, -25, -70, -109, -95, -76, -115, -44,
    -- layer=1 filter=43 channel=85
    -34, -19, -1, -19, -69, -15, -24, -46, 14,
    -- layer=1 filter=43 channel=86
    12, -1, 10, 14, 10, 7, 20, 14, 25,
    -- layer=1 filter=43 channel=87
    -13, -32, 47, 10, 0, 31, 8, 6, -14,
    -- layer=1 filter=43 channel=88
    4, 13, -9, 0, 9, 0, 2, -10, 5,
    -- layer=1 filter=43 channel=89
    -55, -28, -37, -17, -22, -38, -19, -25, -32,
    -- layer=1 filter=43 channel=90
    -6, 79, -2, -26, 12, 11, 9, -56, -7,
    -- layer=1 filter=43 channel=91
    1, -9, -1, 4, -13, -7, -3, -10, -18,
    -- layer=1 filter=43 channel=92
    -15, 27, -60, 1, 7, -7, 41, -16, -1,
    -- layer=1 filter=43 channel=93
    -6, 6, -6, 0, 2, 8, 4, 5, 17,
    -- layer=1 filter=43 channel=94
    -3, -23, -13, -7, -3, -17, 24, 10, 15,
    -- layer=1 filter=43 channel=95
    -70, -67, -37, -75, -101, -86, -97, -111, -49,
    -- layer=1 filter=43 channel=96
    10, 10, 13, 5, 12, 6, 10, 8, 4,
    -- layer=1 filter=43 channel=97
    3, 7, -3, 8, 12, 5, 22, 25, 23,
    -- layer=1 filter=43 channel=98
    11, 48, 32, 30, 1, 1, -11, -9, 23,
    -- layer=1 filter=43 channel=99
    -58, -59, -66, -107, -83, -136, -28, -98, -89,
    -- layer=1 filter=43 channel=100
    -16, -17, -12, -9, -22, -23, 16, -4, -5,
    -- layer=1 filter=43 channel=101
    -9, 1, -1, -11, -16, -23, -12, -15, -20,
    -- layer=1 filter=43 channel=102
    3, -16, -22, -4, 0, -20, 17, 8, -9,
    -- layer=1 filter=43 channel=103
    -11, -32, -26, -29, -36, -28, -17, -24, -26,
    -- layer=1 filter=43 channel=104
    -20, 0, -16, 27, -11, -5, 7, -9, 16,
    -- layer=1 filter=43 channel=105
    -1, 0, -20, 3, 13, 1, 10, 12, 10,
    -- layer=1 filter=43 channel=106
    2, 28, -6, -29, -14, -18, -17, -24, -20,
    -- layer=1 filter=43 channel=107
    3, -3, 5, 0, -3, -5, 9, 4, -2,
    -- layer=1 filter=43 channel=108
    -6, 68, -11, -34, -2, 8, 7, -81, -12,
    -- layer=1 filter=43 channel=109
    -8, 5, 6, 1, 1, -9, -7, 4, -3,
    -- layer=1 filter=43 channel=110
    1, -2, -1, 7, 5, 2, 7, -4, -1,
    -- layer=1 filter=43 channel=111
    -37, -42, 0, -63, -61, -76, -44, -93, -55,
    -- layer=1 filter=43 channel=112
    -10, -10, 22, -58, -49, -39, -40, -66, -25,
    -- layer=1 filter=43 channel=113
    60, 43, 16, 23, 18, 16, 13, 4, -8,
    -- layer=1 filter=43 channel=114
    -24, 28, 48, 37, 20, 32, 46, 4, -7,
    -- layer=1 filter=43 channel=115
    0, -15, -13, 15, 4, -8, 24, 23, 25,
    -- layer=1 filter=43 channel=116
    -8, 0, -1, 1, 10, -1, 8, 6, -3,
    -- layer=1 filter=43 channel=117
    -18, -28, 27, -73, -57, -57, -60, -94, -58,
    -- layer=1 filter=43 channel=118
    -67, -21, -12, -67, -75, -79, -30, -86, -54,
    -- layer=1 filter=43 channel=119
    1, 39, -32, -43, -25, -34, -1, -90, 2,
    -- layer=1 filter=43 channel=120
    -16, -25, -8, -3, -36, -8, 0, -3, -8,
    -- layer=1 filter=43 channel=121
    -9, -31, -15, -20, -8, -18, -22, -13, -22,
    -- layer=1 filter=43 channel=122
    5, -4, 3, -9, -6, -6, -9, 2, 3,
    -- layer=1 filter=43 channel=123
    9, -15, -26, -20, -13, -33, -3, -1, -24,
    -- layer=1 filter=43 channel=124
    4, -9, 0, 3, -7, -6, -15, -13, -14,
    -- layer=1 filter=43 channel=125
    27, 35, 7, -3, -14, 35, -5, 19, 1,
    -- layer=1 filter=43 channel=126
    18, 63, 33, 28, -5, -17, -6, -12, 41,
    -- layer=1 filter=43 channel=127
    -77, -40, -33, -80, -70, -85, -63, -100, -53,
    -- layer=1 filter=44 channel=0
    5, -8, 0, -7, -7, 3, 15, 11, -2,
    -- layer=1 filter=44 channel=1
    -3, -19, -20, -13, 1, 33, 11, 26, 9,
    -- layer=1 filter=44 channel=2
    12, 13, -1, 25, 0, 30, -5, -24, -12,
    -- layer=1 filter=44 channel=3
    3, 6, 4, -1, 3, -1, 1, 0, 10,
    -- layer=1 filter=44 channel=4
    -14, 3, 1, 3, -2, 12, 1, 1, -3,
    -- layer=1 filter=44 channel=5
    -2, -16, -20, 7, 8, 30, 30, 37, 40,
    -- layer=1 filter=44 channel=6
    -7, 19, 21, 15, 52, 39, -3, 24, 36,
    -- layer=1 filter=44 channel=7
    -32, -61, -31, -27, -44, -32, 8, -17, -37,
    -- layer=1 filter=44 channel=8
    21, 25, -6, 5, 33, 45, 20, 13, -18,
    -- layer=1 filter=44 channel=9
    13, 29, 17, 56, 53, 39, 14, -4, -6,
    -- layer=1 filter=44 channel=10
    -24, -80, -45, -30, -16, -27, 32, 34, -4,
    -- layer=1 filter=44 channel=11
    5, 21, 26, -36, -64, -53, 1, -22, 13,
    -- layer=1 filter=44 channel=12
    -2, 16, 38, 97, 85, 78, -17, -27, -29,
    -- layer=1 filter=44 channel=13
    -18, 11, -4, -1, 23, 21, -27, -2, -7,
    -- layer=1 filter=44 channel=14
    1, -61, -18, -12, 2, -4, 17, -15, -63,
    -- layer=1 filter=44 channel=15
    -30, -26, 13, -27, -12, 6, -33, 6, 19,
    -- layer=1 filter=44 channel=16
    13, 33, 8, 6, 30, 33, -12, -19, -11,
    -- layer=1 filter=44 channel=17
    -17, -26, -29, -20, -25, -19, 2, -22, -41,
    -- layer=1 filter=44 channel=18
    16, 23, 30, -5, 6, 9, -44, -54, -39,
    -- layer=1 filter=44 channel=19
    -21, 1, 4, 40, 28, -17, -18, -33, -5,
    -- layer=1 filter=44 channel=20
    -4, 1, 14, 19, 29, 18, -17, -7, 3,
    -- layer=1 filter=44 channel=21
    1, 4, 3, 6, 36, 29, 7, 25, 9,
    -- layer=1 filter=44 channel=22
    0, 18, 13, 7, 24, 17, -25, -20, -34,
    -- layer=1 filter=44 channel=23
    26, -39, -37, 52, -73, -16, 1, -84, 0,
    -- layer=1 filter=44 channel=24
    -13, 17, -6, 16, 17, 14, 7, 10, 6,
    -- layer=1 filter=44 channel=25
    -12, -41, -12, -6, 0, 11, 16, 11, -8,
    -- layer=1 filter=44 channel=26
    9, 30, 1, -3, -5, -22, -36, -41, -38,
    -- layer=1 filter=44 channel=27
    68, 41, 41, 34, 10, 23, 66, 31, 45,
    -- layer=1 filter=44 channel=28
    -28, -30, 5, -32, 0, 19, -2, 3, -38,
    -- layer=1 filter=44 channel=29
    7, 8, -11, 5, 9, 6, 7, 8, 7,
    -- layer=1 filter=44 channel=30
    2, -3, 21, 16, 27, -4, 2, -8, -23,
    -- layer=1 filter=44 channel=31
    23, 12, 20, 33, 29, 44, 29, -3, 28,
    -- layer=1 filter=44 channel=32
    -25, -36, -42, 0, -51, -18, -19, -30, -22,
    -- layer=1 filter=44 channel=33
    6, 5, 2, -10, 1, 3, -9, 1, -4,
    -- layer=1 filter=44 channel=34
    -48, -39, -6, -30, -29, -1, -21, -30, -11,
    -- layer=1 filter=44 channel=35
    0, 0, 9, -2, -5, 8, 1, -7, 7,
    -- layer=1 filter=44 channel=36
    21, -11, 13, -34, -78, -41, 17, -10, 20,
    -- layer=1 filter=44 channel=37
    -30, -4, 0, -20, 11, 17, 16, 35, 40,
    -- layer=1 filter=44 channel=38
    1, 0, 4, 12, 34, 33, 2, 11, 11,
    -- layer=1 filter=44 channel=39
    11, 16, 6, -41, -24, -3, 17, 5, 19,
    -- layer=1 filter=44 channel=40
    23, 10, 15, 11, 35, 30, -1, 10, 19,
    -- layer=1 filter=44 channel=41
    -7, 11, -31, 42, -19, -29, -12, -15, -8,
    -- layer=1 filter=44 channel=42
    18, -1, 8, 30, 10, 31, 4, -11, 12,
    -- layer=1 filter=44 channel=43
    8, 31, -1, 12, 18, 35, 5, 3, -30,
    -- layer=1 filter=44 channel=44
    -33, -8, -22, -24, -42, -29, -20, -17, -15,
    -- layer=1 filter=44 channel=45
    -23, 23, -14, 3, 14, 26, 5, 17, 1,
    -- layer=1 filter=44 channel=46
    -13, -10, 13, 65, 49, 6, 15, 13, 40,
    -- layer=1 filter=44 channel=47
    25, -45, 33, 26, -1, 49, 13, 8, 40,
    -- layer=1 filter=44 channel=48
    -9, 1, 0, 6, 38, 17, 8, 27, 13,
    -- layer=1 filter=44 channel=49
    0, -10, 13, 11, 28, 36, 4, 8, 25,
    -- layer=1 filter=44 channel=50
    -14, -14, -9, -10, 3, -2, -12, -22, -11,
    -- layer=1 filter=44 channel=51
    -1, 5, -17, 18, 42, 18, 10, 24, 7,
    -- layer=1 filter=44 channel=52
    -14, 0, -16, 9, -23, 0, -11, -2, -22,
    -- layer=1 filter=44 channel=53
    -1, 3, 4, -7, -11, -4, -6, -13, -7,
    -- layer=1 filter=44 channel=54
    -25, -46, -38, -3, -22, -9, 11, 9, -14,
    -- layer=1 filter=44 channel=55
    -13, -59, -13, -82, -93, -68, 8, -7, 23,
    -- layer=1 filter=44 channel=56
    -2, 2, -6, 7, 0, 4, -7, -5, 1,
    -- layer=1 filter=44 channel=57
    0, -49, -8, 0, 4, -5, 23, 15, -15,
    -- layer=1 filter=44 channel=58
    20, -60, -31, 26, -34, -39, 52, 0, 2,
    -- layer=1 filter=44 channel=59
    -16, -3, 1, -4, 1, -5, -2, 4, -16,
    -- layer=1 filter=44 channel=60
    -11, -35, -18, 2, -4, 0, -4, 8, -7,
    -- layer=1 filter=44 channel=61
    2, 10, 14, 0, -5, -2, 14, 1, -9,
    -- layer=1 filter=44 channel=62
    -11, 3, -22, -15, 14, 19, -8, -3, -23,
    -- layer=1 filter=44 channel=63
    -12, -8, -20, -55, -74, -52, -10, -44, -2,
    -- layer=1 filter=44 channel=64
    -23, -25, -5, -4, 19, 8, -4, 17, 12,
    -- layer=1 filter=44 channel=65
    -10, 16, 11, 14, 30, 24, -8, 7, -2,
    -- layer=1 filter=44 channel=66
    -3, -21, -5, -27, -39, -15, 14, 1, 23,
    -- layer=1 filter=44 channel=67
    -11, 19, 6, 35, 78, 59, 32, 61, 60,
    -- layer=1 filter=44 channel=68
    -55, 6, -27, -46, -52, -26, -25, -15, 6,
    -- layer=1 filter=44 channel=69
    -10, 7, 17, -28, -9, 25, -6, -24, 4,
    -- layer=1 filter=44 channel=70
    19, -2, 7, 17, 52, 19, 35, 66, 80,
    -- layer=1 filter=44 channel=71
    -6, 9, -33, 6, 14, 4, 2, 13, -2,
    -- layer=1 filter=44 channel=72
    -9, 10, 15, 57, 49, 17, 0, -36, -26,
    -- layer=1 filter=44 channel=73
    3, -5, -6, -9, 3, -12, -7, -2, 0,
    -- layer=1 filter=44 channel=74
    -7, 35, 12, -6, 37, 19, 0, 1, 26,
    -- layer=1 filter=44 channel=75
    3, 4, 4, 26, 11, 24, -36, -45, -40,
    -- layer=1 filter=44 channel=76
    11, 8, 11, 10, -11, -10, -3, -18, -11,
    -- layer=1 filter=44 channel=77
    -23, 13, -10, -15, 27, 35, 3, 16, 19,
    -- layer=1 filter=44 channel=78
    19, -5, 7, -6, 9, -15, 19, 29, -16,
    -- layer=1 filter=44 channel=79
    12, 14, 8, 11, 13, 24, -4, -17, -16,
    -- layer=1 filter=44 channel=80
    18, -10, -10, -10, 25, 4, 0, -34, -19,
    -- layer=1 filter=44 channel=81
    5, 20, -4, -1, 12, 26, -3, 2, 6,
    -- layer=1 filter=44 channel=82
    -4, 17, -20, 16, 45, 32, 5, 30, 12,
    -- layer=1 filter=44 channel=83
    -23, -10, -4, -18, -8, 37, 17, 19, 7,
    -- layer=1 filter=44 channel=84
    23, 33, 15, -12, -10, -27, -58, -40, -34,
    -- layer=1 filter=44 channel=85
    0, -17, -30, 50, 17, 15, 46, 2, 15,
    -- layer=1 filter=44 channel=86
    -11, -30, -11, -68, -84, -51, -11, -11, 13,
    -- layer=1 filter=44 channel=87
    -8, 28, 47, 53, 90, 25, 57, 34, 49,
    -- layer=1 filter=44 channel=88
    -15, 4, -20, 12, 37, 15, 11, 15, 5,
    -- layer=1 filter=44 channel=89
    5, 27, 1, 21, 31, 23, 7, 22, 28,
    -- layer=1 filter=44 channel=90
    -54, -21, -35, -39, -57, -22, -19, -25, 2,
    -- layer=1 filter=44 channel=91
    -14, -1, 1, 0, 31, 27, -7, 13, 23,
    -- layer=1 filter=44 channel=92
    3, -26, 45, -50, -18, 26, -45, -38, 2,
    -- layer=1 filter=44 channel=93
    -14, -3, -9, -5, 20, 0, -6, 12, -1,
    -- layer=1 filter=44 channel=94
    -6, -18, -8, -18, -21, -23, -5, -40, -11,
    -- layer=1 filter=44 channel=95
    -9, 2, -4, -37, -6, -23, -39, -25, -34,
    -- layer=1 filter=44 channel=96
    -30, -17, -13, -13, -7, -22, -7, -2, 1,
    -- layer=1 filter=44 channel=97
    4, -13, -7, -10, -11, -1, -4, -8, -18,
    -- layer=1 filter=44 channel=98
    13, 28, -4, 8, 24, 22, 17, 0, -15,
    -- layer=1 filter=44 channel=99
    -26, -19, -19, -28, 3, 13, 10, 19, -20,
    -- layer=1 filter=44 channel=100
    -16, 14, 15, 7, -45, -26, 35, -22, 33,
    -- layer=1 filter=44 channel=101
    -10, 5, 10, 15, 20, 20, 4, 19, 4,
    -- layer=1 filter=44 channel=102
    -19, -17, -20, -12, -5, -8, -6, -3, 9,
    -- layer=1 filter=44 channel=103
    6, -8, 0, -19, -15, -8, 2, -6, -36,
    -- layer=1 filter=44 channel=104
    24, -9, -19, 23, -11, -7, 10, -25, -3,
    -- layer=1 filter=44 channel=105
    -11, -25, -21, -31, -28, -15, 0, -4, -17,
    -- layer=1 filter=44 channel=106
    3, 10, 12, 14, 13, 25, -4, 7, 21,
    -- layer=1 filter=44 channel=107
    11, -4, -10, 12, -4, 7, -1, 11, -9,
    -- layer=1 filter=44 channel=108
    -4, -17, -33, 3, -30, -22, -6, 0, -10,
    -- layer=1 filter=44 channel=109
    -5, -8, 1, 7, 2, -8, 0, -2, -10,
    -- layer=1 filter=44 channel=110
    13, -9, -5, 3, -8, -6, 3, 9, 4,
    -- layer=1 filter=44 channel=111
    13, 5, 2, -38, 8, -21, -18, -17, -25,
    -- layer=1 filter=44 channel=112
    28, 22, 3, -20, -12, -3, -20, 6, -1,
    -- layer=1 filter=44 channel=113
    -4, -9, 5, 38, 18, 12, 8, 10, -12,
    -- layer=1 filter=44 channel=114
    21, 21, 34, -15, -8, 8, 8, 25, 14,
    -- layer=1 filter=44 channel=115
    -2, -38, -15, -28, -66, -51, -8, -38, -34,
    -- layer=1 filter=44 channel=116
    -8, -5, 7, 7, 4, -5, -3, -6, 0,
    -- layer=1 filter=44 channel=117
    51, 0, -9, -15, 0, 2, -18, -9, -56,
    -- layer=1 filter=44 channel=118
    -5, 14, 7, -11, 13, 7, -11, -16, 11,
    -- layer=1 filter=44 channel=119
    -38, -44, -51, -21, -36, -29, -21, -26, -23,
    -- layer=1 filter=44 channel=120
    -19, -14, -7, -1, 41, 38, 9, 12, 13,
    -- layer=1 filter=44 channel=121
    -29, -52, -22, -7, 1, -34, 9, -21, -23,
    -- layer=1 filter=44 channel=122
    5, -8, 7, 0, 9, -8, -10, 4, 3,
    -- layer=1 filter=44 channel=123
    -14, -48, -18, -26, -31, -33, -21, -37, -19,
    -- layer=1 filter=44 channel=124
    3, 10, 12, 5, -10, 0, 0, 0, -5,
    -- layer=1 filter=44 channel=125
    12, -14, 0, -8, 60, 9, 49, 60, 74,
    -- layer=1 filter=44 channel=126
    -20, 8, -13, 20, 37, 58, 61, 64, 21,
    -- layer=1 filter=44 channel=127
    9, 39, 7, -12, -2, -2, -31, -13, -10,
    -- layer=1 filter=45 channel=0
    -3, -6, -4, 1, -1, -2, 1, -2, -10,
    -- layer=1 filter=45 channel=1
    -3, -3, 4, 6, 2, -1, 7, 5, -3,
    -- layer=1 filter=45 channel=2
    11, 11, 11, 5, 8, 5, -2, 0, -5,
    -- layer=1 filter=45 channel=3
    -1, -3, 4, -10, 0, 2, 0, -1, -2,
    -- layer=1 filter=45 channel=4
    5, 9, -5, 6, -5, 7, -1, -4, -1,
    -- layer=1 filter=45 channel=5
    6, 3, -2, -8, 0, 0, -6, 4, -5,
    -- layer=1 filter=45 channel=6
    -9, -12, 1, 5, 8, -10, 1, -3, -9,
    -- layer=1 filter=45 channel=7
    -5, 1, -11, -8, -12, -5, -12, -10, 3,
    -- layer=1 filter=45 channel=8
    7, -7, 6, -5, 7, 3, 5, -8, 0,
    -- layer=1 filter=45 channel=9
    6, 2, -2, 3, -11, -13, 0, 3, 5,
    -- layer=1 filter=45 channel=10
    0, -1, -7, -6, -5, -7, 0, -3, -12,
    -- layer=1 filter=45 channel=11
    -14, 7, -10, -10, 0, -8, -1, -8, -11,
    -- layer=1 filter=45 channel=12
    6, 7, -9, -5, -5, -8, 6, -2, 6,
    -- layer=1 filter=45 channel=13
    -7, 6, 0, -10, 0, -7, -1, 6, -10,
    -- layer=1 filter=45 channel=14
    5, 0, -3, -4, 0, 5, 3, 1, -6,
    -- layer=1 filter=45 channel=15
    5, -1, 3, -1, -4, 0, -10, 2, -2,
    -- layer=1 filter=45 channel=16
    -3, -3, 9, -3, -10, 5, -13, -9, -3,
    -- layer=1 filter=45 channel=17
    -6, -11, 6, -8, 7, 5, 9, -4, 0,
    -- layer=1 filter=45 channel=18
    -9, -2, -10, -4, 0, -10, -1, -12, 4,
    -- layer=1 filter=45 channel=19
    2, 9, 5, -4, 6, -3, 5, -6, -8,
    -- layer=1 filter=45 channel=20
    3, -9, 1, 8, -1, -9, 4, -1, 5,
    -- layer=1 filter=45 channel=21
    -9, -1, -7, -3, 5, -9, -3, -8, 6,
    -- layer=1 filter=45 channel=22
    -7, -8, -4, -13, -4, -11, 1, -6, -11,
    -- layer=1 filter=45 channel=23
    -9, -7, -2, -6, -8, -9, -10, -11, 1,
    -- layer=1 filter=45 channel=24
    -5, -6, -1, -4, -5, 5, 4, 7, 4,
    -- layer=1 filter=45 channel=25
    -12, -11, 4, 0, 4, -10, -13, -9, -7,
    -- layer=1 filter=45 channel=26
    7, 9, 6, 0, -11, -10, -2, -2, 8,
    -- layer=1 filter=45 channel=27
    9, -4, -3, -7, 6, -3, -6, -1, -1,
    -- layer=1 filter=45 channel=28
    4, 0, 0, -3, 1, 0, 8, 3, 8,
    -- layer=1 filter=45 channel=29
    -3, 5, 2, -9, 7, 3, -9, -1, -1,
    -- layer=1 filter=45 channel=30
    -10, -1, 2, -2, 8, -6, -9, -4, 3,
    -- layer=1 filter=45 channel=31
    1, 0, 4, 0, 0, -1, -2, -1, -12,
    -- layer=1 filter=45 channel=32
    -9, 0, 5, -9, 8, 6, 6, 5, 6,
    -- layer=1 filter=45 channel=33
    -7, -4, 6, 11, 0, 9, -1, 1, 4,
    -- layer=1 filter=45 channel=34
    -11, 4, 6, -7, -6, 5, 8, 8, -5,
    -- layer=1 filter=45 channel=35
    1, -2, -11, -1, -8, -6, -8, 9, 8,
    -- layer=1 filter=45 channel=36
    -10, -1, 7, 1, -10, 7, 0, -11, 7,
    -- layer=1 filter=45 channel=37
    6, -9, 6, 4, -12, -4, 1, -6, -10,
    -- layer=1 filter=45 channel=38
    4, 3, -6, 2, 1, -2, -4, 5, -3,
    -- layer=1 filter=45 channel=39
    -4, -5, -11, 1, 2, -11, -7, -5, -2,
    -- layer=1 filter=45 channel=40
    8, -4, -4, -11, 8, 0, 4, -5, 0,
    -- layer=1 filter=45 channel=41
    -10, -3, 0, -8, -9, -4, -1, -8, -4,
    -- layer=1 filter=45 channel=42
    -3, 1, 2, -1, 10, 0, -5, 8, -5,
    -- layer=1 filter=45 channel=43
    -2, 9, 0, -4, 2, 3, -9, -6, 4,
    -- layer=1 filter=45 channel=44
    6, -5, -9, 0, -9, 8, 1, -9, -9,
    -- layer=1 filter=45 channel=45
    5, 8, 0, 0, -4, 0, -2, 8, 3,
    -- layer=1 filter=45 channel=46
    -1, 0, -9, -9, -7, -1, 0, -10, -12,
    -- layer=1 filter=45 channel=47
    0, -4, -7, 9, -15, -8, -4, -11, -4,
    -- layer=1 filter=45 channel=48
    -6, -3, 1, -3, 6, 0, -10, -11, 1,
    -- layer=1 filter=45 channel=49
    -9, 1, -8, 0, -11, -6, -5, -4, 0,
    -- layer=1 filter=45 channel=50
    -4, 6, -3, 2, -8, 2, -11, -6, -7,
    -- layer=1 filter=45 channel=51
    0, 9, 1, -1, -2, -9, 5, 0, -4,
    -- layer=1 filter=45 channel=52
    3, -7, 2, -2, -1, -4, -9, -8, 6,
    -- layer=1 filter=45 channel=53
    -9, -8, -1, 4, 4, -10, -6, 0, -5,
    -- layer=1 filter=45 channel=54
    1, -7, 0, 0, -7, -4, 3, 7, 4,
    -- layer=1 filter=45 channel=55
    -9, 2, -3, 0, -7, -9, 7, -5, -1,
    -- layer=1 filter=45 channel=56
    -4, 2, -3, -3, 4, -1, 8, 0, 8,
    -- layer=1 filter=45 channel=57
    -8, 2, -9, -12, 1, 1, -6, 3, 3,
    -- layer=1 filter=45 channel=58
    -4, -5, 4, -6, -9, 0, 0, -4, -9,
    -- layer=1 filter=45 channel=59
    7, 6, -4, -8, -2, -7, 5, 8, -6,
    -- layer=1 filter=45 channel=60
    0, -4, 1, -8, 12, 8, 1, 1, 0,
    -- layer=1 filter=45 channel=61
    -1, -5, -11, -2, 1, 2, -8, 9, 3,
    -- layer=1 filter=45 channel=62
    -6, -9, 0, -3, -13, -1, 6, 0, -7,
    -- layer=1 filter=45 channel=63
    5, -2, 0, -1, -5, 7, 6, -5, 6,
    -- layer=1 filter=45 channel=64
    0, -6, 5, -6, -2, 0, 0, -6, -8,
    -- layer=1 filter=45 channel=65
    -2, 1, -7, 8, 9, 2, 3, -11, 0,
    -- layer=1 filter=45 channel=66
    0, 0, 7, 0, 1, 2, 0, 5, -9,
    -- layer=1 filter=45 channel=67
    7, -8, -3, 6, -1, -5, 7, -10, -2,
    -- layer=1 filter=45 channel=68
    -3, 9, 8, 3, -12, -4, 1, 1, 0,
    -- layer=1 filter=45 channel=69
    0, -3, -3, -2, -10, 1, -9, -9, -5,
    -- layer=1 filter=45 channel=70
    -6, -7, -8, 6, 6, 7, 4, -4, 3,
    -- layer=1 filter=45 channel=71
    3, -3, -3, 2, 7, 8, 3, -2, -5,
    -- layer=1 filter=45 channel=72
    -1, -3, 0, -5, -11, 8, 2, -3, -2,
    -- layer=1 filter=45 channel=73
    -2, -10, -2, -10, -5, -5, 2, -5, -7,
    -- layer=1 filter=45 channel=74
    5, 6, 4, 0, 8, -11, -10, -4, 1,
    -- layer=1 filter=45 channel=75
    5, 2, -6, -6, -8, 3, 5, 0, 4,
    -- layer=1 filter=45 channel=76
    -3, -10, 2, 7, 7, -9, -7, -11, 5,
    -- layer=1 filter=45 channel=77
    2, 8, -11, -1, 0, 2, 8, -7, -9,
    -- layer=1 filter=45 channel=78
    0, 7, -7, 6, -7, -7, 0, 4, 8,
    -- layer=1 filter=45 channel=79
    4, 2, -1, 4, -10, -12, 2, -10, 3,
    -- layer=1 filter=45 channel=80
    2, -12, -8, -10, 6, -7, 7, -9, -1,
    -- layer=1 filter=45 channel=81
    -12, -7, -9, -11, -3, -11, -4, 0, 9,
    -- layer=1 filter=45 channel=82
    0, -7, 7, 3, 8, 8, -5, 9, -9,
    -- layer=1 filter=45 channel=83
    -6, -1, -1, 7, 4, 7, -2, -7, 1,
    -- layer=1 filter=45 channel=84
    -2, -6, -7, 0, -2, 3, -5, 5, 1,
    -- layer=1 filter=45 channel=85
    4, -5, -8, 0, -11, 0, 3, -8, -8,
    -- layer=1 filter=45 channel=86
    0, -7, 6, 0, -1, -8, 6, 2, -6,
    -- layer=1 filter=45 channel=87
    7, 3, 1, 1, 7, -2, 0, 7, -3,
    -- layer=1 filter=45 channel=88
    -5, -4, 0, 4, -9, -2, -9, -9, -5,
    -- layer=1 filter=45 channel=89
    -7, 1, -6, 7, -1, 4, -10, -3, -3,
    -- layer=1 filter=45 channel=90
    5, -1, 3, -5, -2, -2, 7, 4, -3,
    -- layer=1 filter=45 channel=91
    1, 2, -7, -9, -9, 2, 0, -7, -1,
    -- layer=1 filter=45 channel=92
    7, -2, 2, 7, -8, 5, 6, -8, -2,
    -- layer=1 filter=45 channel=93
    -5, 5, 8, -4, -10, -5, 7, 2, -9,
    -- layer=1 filter=45 channel=94
    2, 8, -6, 1, -8, 5, -10, -4, 4,
    -- layer=1 filter=45 channel=95
    0, 0, 7, 0, -4, 3, -12, 5, 0,
    -- layer=1 filter=45 channel=96
    -8, -7, 3, 0, 0, 0, 5, 8, -8,
    -- layer=1 filter=45 channel=97
    7, 8, -9, 7, -11, -10, 1, 8, 5,
    -- layer=1 filter=45 channel=98
    -13, -10, -6, -13, -16, 5, -6, -1, -4,
    -- layer=1 filter=45 channel=99
    3, 0, 0, -2, -9, -7, -10, -3, 8,
    -- layer=1 filter=45 channel=100
    1, -11, -5, -10, -1, -12, -3, -4, -7,
    -- layer=1 filter=45 channel=101
    -5, 5, -2, 7, 2, -8, 3, 3, -4,
    -- layer=1 filter=45 channel=102
    -8, -10, -7, -5, 8, 6, -11, 8, 1,
    -- layer=1 filter=45 channel=103
    -5, -4, 4, 3, -6, 2, -8, -11, 5,
    -- layer=1 filter=45 channel=104
    7, 2, 1, -5, 7, 3, 0, 8, -2,
    -- layer=1 filter=45 channel=105
    7, -6, -8, -1, -2, -8, 6, -4, -7,
    -- layer=1 filter=45 channel=106
    8, -3, 0, -1, -11, -6, 3, -7, -14,
    -- layer=1 filter=45 channel=107
    -7, 2, 0, 4, -8, 0, -2, 2, -8,
    -- layer=1 filter=45 channel=108
    1, 0, -5, -8, -1, -2, -11, -15, -8,
    -- layer=1 filter=45 channel=109
    8, -1, -4, 1, -2, -9, 3, -6, -6,
    -- layer=1 filter=45 channel=110
    0, 8, 6, -3, -7, 5, -3, -8, -6,
    -- layer=1 filter=45 channel=111
    2, 3, -1, -6, -1, -8, 0, 1, -11,
    -- layer=1 filter=45 channel=112
    -7, -9, 0, 3, 1, -3, -3, -3, -3,
    -- layer=1 filter=45 channel=113
    -1, 2, -7, -1, 0, -6, 9, -4, 11,
    -- layer=1 filter=45 channel=114
    -3, -4, -3, -5, 0, -3, 9, -5, -4,
    -- layer=1 filter=45 channel=115
    -8, -1, -9, 5, 8, 9, -6, 8, 8,
    -- layer=1 filter=45 channel=116
    -7, 3, 0, -6, -1, -6, -10, -4, -2,
    -- layer=1 filter=45 channel=117
    4, -10, 2, -8, 4, 0, 10, -3, -3,
    -- layer=1 filter=45 channel=118
    -6, -5, -8, 6, -9, 4, -8, 5, -13,
    -- layer=1 filter=45 channel=119
    -9, -9, -7, -10, -11, -4, 7, -1, -10,
    -- layer=1 filter=45 channel=120
    -7, -1, -9, -8, -1, -1, -12, -4, 6,
    -- layer=1 filter=45 channel=121
    -4, -13, 0, -10, 6, 5, -13, -14, -7,
    -- layer=1 filter=45 channel=122
    6, 6, -4, -1, 3, -3, -3, -9, 1,
    -- layer=1 filter=45 channel=123
    -9, -10, 1, 1, -4, -4, 8, -9, -9,
    -- layer=1 filter=45 channel=124
    4, -2, 3, -10, -1, -9, 0, 2, -8,
    -- layer=1 filter=45 channel=125
    8, -5, -12, 2, 2, 1, -8, -3, 0,
    -- layer=1 filter=45 channel=126
    -5, 8, 0, 0, -7, 1, -4, 0, 2,
    -- layer=1 filter=45 channel=127
    -11, -6, -11, -9, -5, 3, -5, -4, -1,
    -- layer=1 filter=46 channel=0
    -18, -16, 0, 6, 14, 5, -18, -5, 10,
    -- layer=1 filter=46 channel=1
    28, 31, 5, 18, 4, -8, -37, -7, -13,
    -- layer=1 filter=46 channel=2
    45, 44, 46, 42, 31, 21, 15, 11, -25,
    -- layer=1 filter=46 channel=3
    11, 13, 7, 10, -1, 5, 11, -1, 19,
    -- layer=1 filter=46 channel=4
    10, 2, 5, -2, -2, -15, 14, 13, 0,
    -- layer=1 filter=46 channel=5
    18, 39, 2, 24, 3, -9, 2, 17, -2,
    -- layer=1 filter=46 channel=6
    -14, -22, -22, 0, -3, 15, 28, 26, 15,
    -- layer=1 filter=46 channel=7
    -27, -15, -7, -41, -38, -21, -20, -30, 0,
    -- layer=1 filter=46 channel=8
    35, 32, 3, 47, 9, -1, 4, 18, 10,
    -- layer=1 filter=46 channel=9
    -7, -13, -5, -57, -42, -19, -1, -16, -50,
    -- layer=1 filter=46 channel=10
    -3, -29, 11, -14, -35, -14, 8, -4, 8,
    -- layer=1 filter=46 channel=11
    -17, -30, -21, 8, 3, -4, 3, -3, 2,
    -- layer=1 filter=46 channel=12
    21, 37, 26, -32, -5, -49, -7, -30, -50,
    -- layer=1 filter=46 channel=13
    4, -4, 15, -14, -1, 10, -17, -2, 1,
    -- layer=1 filter=46 channel=14
    -7, 0, 0, -26, -38, -17, -5, -53, -5,
    -- layer=1 filter=46 channel=15
    22, -2, -26, 46, -14, -11, -17, 2, -22,
    -- layer=1 filter=46 channel=16
    49, 40, 22, 26, 19, 6, 20, 11, 1,
    -- layer=1 filter=46 channel=17
    -1, 2, 6, 4, 17, 23, -19, -10, -9,
    -- layer=1 filter=46 channel=18
    6, 15, 23, 13, 41, 5, 29, 11, 14,
    -- layer=1 filter=46 channel=19
    39, 43, 38, 61, 46, 32, 36, 60, 26,
    -- layer=1 filter=46 channel=20
    12, 8, 18, 11, 20, 30, -4, 5, 9,
    -- layer=1 filter=46 channel=21
    -8, 5, -3, 12, -1, 1, -17, -20, -11,
    -- layer=1 filter=46 channel=22
    19, 22, 2, 43, 27, 49, -12, 4, 0,
    -- layer=1 filter=46 channel=23
    -33, -27, -17, -88, -72, -31, -73, -57, -71,
    -- layer=1 filter=46 channel=24
    12, -3, -1, -1, -1, 3, 1, -25, -8,
    -- layer=1 filter=46 channel=25
    6, 36, 33, -13, 0, 13, 11, 0, 13,
    -- layer=1 filter=46 channel=26
    12, 0, -8, -16, -31, -20, -4, -53, -15,
    -- layer=1 filter=46 channel=27
    26, 21, 6, 47, 38, 30, 69, 56, 36,
    -- layer=1 filter=46 channel=28
    0, -6, 8, -19, -35, -6, -17, -25, 7,
    -- layer=1 filter=46 channel=29
    -11, -8, -15, 2, 9, -1, 13, 2, 13,
    -- layer=1 filter=46 channel=30
    11, 7, 10, 20, 35, -11, 49, 54, -2,
    -- layer=1 filter=46 channel=31
    31, 33, 30, 18, 32, 28, 7, 9, 8,
    -- layer=1 filter=46 channel=32
    -33, -68, -48, -75, -104, -56, -8, -108, -44,
    -- layer=1 filter=46 channel=33
    11, 13, -12, 2, 19, 5, -1, 0, 4,
    -- layer=1 filter=46 channel=34
    16, 12, -23, 14, -13, -10, 4, -3, -8,
    -- layer=1 filter=46 channel=35
    7, 4, -18, -15, -12, -25, -16, -13, -22,
    -- layer=1 filter=46 channel=36
    -18, -18, -26, -2, -7, 3, -1, 3, 7,
    -- layer=1 filter=46 channel=37
    42, 43, 19, 22, 21, 10, 29, 21, 38,
    -- layer=1 filter=46 channel=38
    -10, -4, -11, -7, 7, 15, 7, 15, 9,
    -- layer=1 filter=46 channel=39
    -16, -2, -5, 3, -1, -5, -12, -19, -1,
    -- layer=1 filter=46 channel=40
    17, -3, 9, 20, 16, 22, 33, 30, 17,
    -- layer=1 filter=46 channel=41
    -6, -42, -6, -70, -77, -76, -10, -40, -92,
    -- layer=1 filter=46 channel=42
    33, 53, 39, 44, 49, 24, 21, 5, -6,
    -- layer=1 filter=46 channel=43
    35, 48, 20, 15, 12, 11, 0, 17, 0,
    -- layer=1 filter=46 channel=44
    -52, -73, -52, -63, -89, -52, -17, -89, -39,
    -- layer=1 filter=46 channel=45
    -10, 3, -22, -3, -6, -1, -18, -17, -6,
    -- layer=1 filter=46 channel=46
    84, 84, 45, 91, 62, 28, 73, 46, 8,
    -- layer=1 filter=46 channel=47
    -38, -76, -27, -77, -77, -42, -70, -60, -32,
    -- layer=1 filter=46 channel=48
    -9, -16, -5, 1, 4, 4, 2, 7, 6,
    -- layer=1 filter=46 channel=49
    2, 3, 2, -4, 21, 11, 8, -5, -6,
    -- layer=1 filter=46 channel=50
    14, 6, 9, 7, 9, 8, 9, -2, 18,
    -- layer=1 filter=46 channel=51
    -24, -23, -2, -16, -9, -9, -4, -1, 5,
    -- layer=1 filter=46 channel=52
    9, 13, 5, 28, 18, 12, 7, 8, -6,
    -- layer=1 filter=46 channel=53
    22, 23, 28, 15, 23, 20, 19, 30, 33,
    -- layer=1 filter=46 channel=54
    35, 35, 27, -1, -2, -1, 24, 13, 12,
    -- layer=1 filter=46 channel=55
    -15, -18, -22, 21, 2, -11, 8, 16, 8,
    -- layer=1 filter=46 channel=56
    -2, 4, 0, 4, -9, -6, -14, 4, -1,
    -- layer=1 filter=46 channel=57
    7, -10, 24, 7, 3, 16, 19, 7, 44,
    -- layer=1 filter=46 channel=58
    -61, -76, 7, -124, -100, -73, -59, -64, -81,
    -- layer=1 filter=46 channel=59
    25, 12, 5, 34, 3, 7, -9, -9, -34,
    -- layer=1 filter=46 channel=60
    6, 2, 8, 4, 19, 23, 4, 9, 4,
    -- layer=1 filter=46 channel=61
    -5, 9, 8, 13, 0, 6, 6, 7, -5,
    -- layer=1 filter=46 channel=62
    40, 56, 31, 33, 23, 10, 18, 14, 7,
    -- layer=1 filter=46 channel=63
    -27, -20, -15, -5, 1, -12, 23, 11, 11,
    -- layer=1 filter=46 channel=64
    0, 17, 9, 7, 12, 21, -7, -1, 4,
    -- layer=1 filter=46 channel=65
    -13, -8, 10, 2, -6, 10, -10, -4, 3,
    -- layer=1 filter=46 channel=66
    0, -6, -10, -4, 10, 6, -6, 0, 7,
    -- layer=1 filter=46 channel=67
    -12, -14, -23, 31, 38, 29, 28, 44, 26,
    -- layer=1 filter=46 channel=68
    -60, -97, -56, -97, -92, -74, -24, -118, -71,
    -- layer=1 filter=46 channel=69
    18, 20, -10, 4, -11, -8, 11, 9, 0,
    -- layer=1 filter=46 channel=70
    15, -2, -9, 23, 27, 8, 33, 13, 20,
    -- layer=1 filter=46 channel=71
    0, 19, -6, 19, -6, 6, 28, 27, 0,
    -- layer=1 filter=46 channel=72
    27, 17, 23, 37, 29, 5, 62, 54, 21,
    -- layer=1 filter=46 channel=73
    -3, 5, 10, 3, -6, 12, -4, 8, 1,
    -- layer=1 filter=46 channel=74
    -16, -18, -5, -19, 0, -8, 6, -19, 3,
    -- layer=1 filter=46 channel=75
    0, -4, 0, -12, 3, -18, 25, 0, -11,
    -- layer=1 filter=46 channel=76
    -44, -37, -15, -18, 4, -11, 13, -1, -1,
    -- layer=1 filter=46 channel=77
    -11, -12, -4, -1, 7, 6, -14, -9, 9,
    -- layer=1 filter=46 channel=78
    -15, -13, -13, -17, -15, -11, -4, -1, 0,
    -- layer=1 filter=46 channel=79
    39, 36, 29, 29, 20, 4, -9, 6, 9,
    -- layer=1 filter=46 channel=80
    5, -6, 3, 25, 9, -2, -2, -7, -9,
    -- layer=1 filter=46 channel=81
    17, -2, -15, 23, 18, 5, 11, 1, 1,
    -- layer=1 filter=46 channel=82
    -17, -4, -9, -2, 11, 10, -19, -17, -14,
    -- layer=1 filter=46 channel=83
    -24, -3, -3, -3, -6, -25, -38, -13, -8,
    -- layer=1 filter=46 channel=84
    34, 28, 37, 19, 40, 0, 36, 18, -2,
    -- layer=1 filter=46 channel=85
    -36, -26, -3, -96, -99, -57, -84, -48, -59,
    -- layer=1 filter=46 channel=86
    -8, 11, 6, 12, 15, 6, 9, 9, 2,
    -- layer=1 filter=46 channel=87
    55, 59, 34, 21, 26, -14, 44, 47, 10,
    -- layer=1 filter=46 channel=88
    23, 7, -3, 19, 19, 30, 15, 24, 28,
    -- layer=1 filter=46 channel=89
    -9, -20, -22, -13, -4, -7, -4, 0, -20,
    -- layer=1 filter=46 channel=90
    -45, -76, -66, -76, -96, -67, -46, -120, -74,
    -- layer=1 filter=46 channel=91
    -13, 5, -5, -6, 24, 8, -1, 23, 27,
    -- layer=1 filter=46 channel=92
    11, -71, -11, -37, -7, -39, -42, -59, -47,
    -- layer=1 filter=46 channel=93
    -10, -2, 6, 3, 1, 1, -7, -8, -5,
    -- layer=1 filter=46 channel=94
    -15, -18, -1, -1, 13, 8, -7, -4, 7,
    -- layer=1 filter=46 channel=95
    24, 22, 21, 5, 27, -5, 48, 8, 15,
    -- layer=1 filter=46 channel=96
    -2, -5, 2, 13, 18, 11, -9, 11, -11,
    -- layer=1 filter=46 channel=97
    4, -3, -5, 6, 1, 17, -21, -10, 6,
    -- layer=1 filter=46 channel=98
    39, 37, 21, 30, 29, 12, 6, 9, -4,
    -- layer=1 filter=46 channel=99
    -46, -102, -57, -53, -85, -54, -48, -76, -15,
    -- layer=1 filter=46 channel=100
    -27, -19, -16, 3, -3, -1, 11, -1, 11,
    -- layer=1 filter=46 channel=101
    -17, -8, -10, -6, 18, 23, 3, 13, 0,
    -- layer=1 filter=46 channel=102
    -29, -25, -8, 8, 3, 21, -10, 1, 8,
    -- layer=1 filter=46 channel=103
    -9, -4, -10, 10, 15, 6, -2, 17, 3,
    -- layer=1 filter=46 channel=104
    -30, 3, 17, -61, -50, -21, -51, -1, -45,
    -- layer=1 filter=46 channel=105
    -11, 1, 1, 8, 8, 12, -6, -7, 7,
    -- layer=1 filter=46 channel=106
    -8, -18, -8, -3, 8, 0, 15, -1, -2,
    -- layer=1 filter=46 channel=107
    -9, 4, -26, 2, 3, 8, 10, 5, 9,
    -- layer=1 filter=46 channel=108
    -20, -77, -66, -57, -95, -75, -29, -116, -69,
    -- layer=1 filter=46 channel=109
    -6, -6, 1, 4, 7, 0, -3, 1, 7,
    -- layer=1 filter=46 channel=110
    -10, 0, -1, -2, 1, -5, -16, 4, -3,
    -- layer=1 filter=46 channel=111
    22, 5, 18, 23, 23, -7, 31, 12, 3,
    -- layer=1 filter=46 channel=112
    24, 38, 20, 27, 43, 14, 21, -21, -9,
    -- layer=1 filter=46 channel=113
    19, 45, 41, 27, 22, 36, 7, 18, 6,
    -- layer=1 filter=46 channel=114
    44, 24, 7, 26, -4, -9, 12, 24, 0,
    -- layer=1 filter=46 channel=115
    -13, 5, 12, 7, 19, 30, -9, 14, 25,
    -- layer=1 filter=46 channel=116
    -7, -4, 0, 4, 3, 5, -9, -1, -8,
    -- layer=1 filter=46 channel=117
    78, 53, 59, 65, 56, 21, 23, -13, 1,
    -- layer=1 filter=46 channel=118
    17, 1, -1, -10, 2, 0, 32, 3, -10,
    -- layer=1 filter=46 channel=119
    -38, -86, -65, -93, -97, -93, -16, -130, -70,
    -- layer=1 filter=46 channel=120
    0, 1, -7, -13, 2, -2, -8, -21, 11,
    -- layer=1 filter=46 channel=121
    30, 27, 8, 55, 40, 14, 77, 46, 34,
    -- layer=1 filter=46 channel=122
    5, 0, 2, -6, -4, 0, 3, -2, 4,
    -- layer=1 filter=46 channel=123
    0, 6, -6, 39, 25, 8, 50, 47, 19,
    -- layer=1 filter=46 channel=124
    -12, -5, -3, -4, 4, 8, -1, 0, 0,
    -- layer=1 filter=46 channel=125
    0, 0, -9, 9, 28, 0, 37, 19, 22,
    -- layer=1 filter=46 channel=126
    17, 38, 7, 65, 37, 17, -16, -12, -10,
    -- layer=1 filter=46 channel=127
    9, 18, 15, 17, 30, 10, 48, 23, 11,
    -- layer=1 filter=47 channel=0
    -3, -12, 6, 7, 0, 1, 6, 1, -1,
    -- layer=1 filter=47 channel=1
    8, 7, -1, 2, 8, -8, 9, -4, -8,
    -- layer=1 filter=47 channel=2
    -2, 8, 6, -7, -5, -1, 1, 3, -2,
    -- layer=1 filter=47 channel=3
    6, -10, -1, -7, -2, 3, -2, -7, 5,
    -- layer=1 filter=47 channel=4
    -9, -4, 6, -6, 1, 7, 9, -9, -8,
    -- layer=1 filter=47 channel=5
    -9, 6, -5, -7, 7, 0, -6, -9, 1,
    -- layer=1 filter=47 channel=6
    6, -9, 3, 5, 0, 0, -9, 0, 0,
    -- layer=1 filter=47 channel=7
    -7, -12, -8, -5, 0, -9, -4, 5, -11,
    -- layer=1 filter=47 channel=8
    6, 0, 7, 0, 0, -5, 4, 3, 6,
    -- layer=1 filter=47 channel=9
    7, -11, 7, -13, 0, -10, -5, -4, 3,
    -- layer=1 filter=47 channel=10
    -11, 4, -6, -6, 6, -10, -6, 4, -9,
    -- layer=1 filter=47 channel=11
    0, -1, 6, -4, 6, 5, 4, -5, 6,
    -- layer=1 filter=47 channel=12
    5, 1, 4, -6, 1, -2, -5, -11, -5,
    -- layer=1 filter=47 channel=13
    -8, -5, 7, -8, -1, -3, -4, -8, 0,
    -- layer=1 filter=47 channel=14
    4, 7, -10, -4, -1, -3, -5, 2, -1,
    -- layer=1 filter=47 channel=15
    -2, -7, -5, -3, 1, -6, -10, 7, -9,
    -- layer=1 filter=47 channel=16
    4, 4, 2, -11, -11, -10, -8, 6, 1,
    -- layer=1 filter=47 channel=17
    5, 3, 1, 2, -4, 7, 2, -8, 7,
    -- layer=1 filter=47 channel=18
    2, 0, -2, 0, -11, 10, 0, -7, 7,
    -- layer=1 filter=47 channel=19
    8, -8, 0, 6, -2, -10, -1, -4, 6,
    -- layer=1 filter=47 channel=20
    -6, -2, -7, -11, -9, 3, 7, -11, 2,
    -- layer=1 filter=47 channel=21
    -7, 7, 4, 3, 7, 7, -3, 5, 1,
    -- layer=1 filter=47 channel=22
    -4, 1, -2, -5, 9, -8, -2, 4, -9,
    -- layer=1 filter=47 channel=23
    -2, -8, 7, -6, 9, -4, 8, 2, 2,
    -- layer=1 filter=47 channel=24
    5, 4, -2, -6, 7, 4, 3, -11, -13,
    -- layer=1 filter=47 channel=25
    -2, -6, 0, 5, 3, -7, 3, 6, -6,
    -- layer=1 filter=47 channel=26
    -6, -8, -11, -5, 4, 0, 3, -2, -5,
    -- layer=1 filter=47 channel=27
    -4, 3, 1, 9, -6, -10, -8, 3, -11,
    -- layer=1 filter=47 channel=28
    -10, -4, -7, 1, -10, -7, -8, -10, 8,
    -- layer=1 filter=47 channel=29
    4, -1, 0, -7, -1, -8, 2, -9, 6,
    -- layer=1 filter=47 channel=30
    6, 0, 2, 0, 6, -1, -7, -12, -9,
    -- layer=1 filter=47 channel=31
    1, -10, -13, -7, 0, -12, 5, 3, 0,
    -- layer=1 filter=47 channel=32
    5, -12, 2, 0, -3, 8, 5, -6, 7,
    -- layer=1 filter=47 channel=33
    2, -8, 5, 0, -8, -3, 7, -2, -4,
    -- layer=1 filter=47 channel=34
    4, 0, -6, 7, -5, -3, 0, 1, -5,
    -- layer=1 filter=47 channel=35
    -1, -5, -10, 7, -9, 0, -6, 3, -1,
    -- layer=1 filter=47 channel=36
    -1, -8, 4, -3, 9, -5, -3, 7, 8,
    -- layer=1 filter=47 channel=37
    -8, -10, -16, -2, -9, 8, 9, -10, -4,
    -- layer=1 filter=47 channel=38
    7, -2, -11, -5, 6, -11, -9, -8, 0,
    -- layer=1 filter=47 channel=39
    -11, 9, -5, -5, -10, -4, -3, -3, -1,
    -- layer=1 filter=47 channel=40
    5, -3, -8, 0, 0, 4, 8, -7, -2,
    -- layer=1 filter=47 channel=41
    5, 1, 6, 8, -3, 2, 0, 1, 3,
    -- layer=1 filter=47 channel=42
    -10, 9, 9, -6, 2, -8, 7, 0, -4,
    -- layer=1 filter=47 channel=43
    6, -7, 5, 0, 7, -9, 1, -8, 4,
    -- layer=1 filter=47 channel=44
    -9, 6, -10, 8, 4, -1, -4, -3, -6,
    -- layer=1 filter=47 channel=45
    -2, 2, 7, 7, 7, -8, -4, -10, 5,
    -- layer=1 filter=47 channel=46
    3, 6, -5, 6, 8, 0, 7, -5, 5,
    -- layer=1 filter=47 channel=47
    2, -4, -7, -13, -13, -8, -6, -8, -12,
    -- layer=1 filter=47 channel=48
    3, -3, 8, 5, -9, 7, 3, -2, -5,
    -- layer=1 filter=47 channel=49
    -9, -12, 0, 7, -9, -11, 1, 4, -5,
    -- layer=1 filter=47 channel=50
    0, 0, 1, -7, 8, -1, 5, -1, 0,
    -- layer=1 filter=47 channel=51
    -7, 5, 4, 7, 6, 6, 6, 2, 3,
    -- layer=1 filter=47 channel=52
    -2, 0, -5, -7, 6, -4, 1, -10, 9,
    -- layer=1 filter=47 channel=53
    7, 0, -3, 1, 3, 4, 8, -5, -4,
    -- layer=1 filter=47 channel=54
    4, -1, 0, 8, 0, -11, 8, -8, -2,
    -- layer=1 filter=47 channel=55
    -4, 5, 7, -8, -7, -4, -9, 8, -6,
    -- layer=1 filter=47 channel=56
    -5, -4, 7, 0, -1, 4, -9, -5, 2,
    -- layer=1 filter=47 channel=57
    9, 7, 4, -7, 4, -2, -3, -5, 0,
    -- layer=1 filter=47 channel=58
    -12, 1, -5, -4, -2, 8, 0, -4, 4,
    -- layer=1 filter=47 channel=59
    8, 0, -7, -3, -1, 4, 9, 6, 5,
    -- layer=1 filter=47 channel=60
    -1, 6, -7, -7, -3, -1, -10, 0, 1,
    -- layer=1 filter=47 channel=61
    -1, 7, 5, 0, 0, 8, 1, -1, -2,
    -- layer=1 filter=47 channel=62
    0, -9, -3, 1, -8, 9, 4, -4, -13,
    -- layer=1 filter=47 channel=63
    -5, -1, 1, -1, 6, -7, 5, -9, 3,
    -- layer=1 filter=47 channel=64
    -11, -9, -6, 9, 8, 0, -6, -6, -9,
    -- layer=1 filter=47 channel=65
    2, -2, -5, -3, -2, -7, -1, -7, 2,
    -- layer=1 filter=47 channel=66
    -2, 2, -3, -9, 7, -8, 8, -3, -9,
    -- layer=1 filter=47 channel=67
    0, 1, 4, 7, 5, -5, 3, 10, 4,
    -- layer=1 filter=47 channel=68
    -7, 2, -8, 2, -3, -1, -6, 1, -1,
    -- layer=1 filter=47 channel=69
    -6, 4, -10, 7, -1, 2, 0, -9, -6,
    -- layer=1 filter=47 channel=70
    4, -8, -9, -5, -1, -10, -4, 1, 8,
    -- layer=1 filter=47 channel=71
    -5, 3, -9, 6, 0, 1, -2, 5, 3,
    -- layer=1 filter=47 channel=72
    5, -10, 1, 2, -6, -8, -9, -9, -11,
    -- layer=1 filter=47 channel=73
    -4, 7, -1, -7, -2, -9, 9, -11, 7,
    -- layer=1 filter=47 channel=74
    1, 7, 5, 0, -5, -8, -1, -2, -8,
    -- layer=1 filter=47 channel=75
    5, -4, 0, -4, -7, 0, 0, -7, 3,
    -- layer=1 filter=47 channel=76
    7, -11, 8, 4, 9, 3, 4, 1, 3,
    -- layer=1 filter=47 channel=77
    -1, -9, 8, -6, 4, 5, -7, -11, -1,
    -- layer=1 filter=47 channel=78
    7, 2, -10, -1, -7, -4, -4, -5, -4,
    -- layer=1 filter=47 channel=79
    -9, 0, -6, -7, 4, 7, -12, 8, 7,
    -- layer=1 filter=47 channel=80
    4, -3, 4, 8, 9, 1, -3, -10, -7,
    -- layer=1 filter=47 channel=81
    1, -3, 1, -9, -5, 6, 3, 1, -2,
    -- layer=1 filter=47 channel=82
    1, 0, -9, -9, -7, 1, 0, 3, -6,
    -- layer=1 filter=47 channel=83
    -3, 1, 8, 8, -3, 2, -1, -1, -2,
    -- layer=1 filter=47 channel=84
    -11, 1, -4, 3, 4, -3, 0, 6, -6,
    -- layer=1 filter=47 channel=85
    7, -8, -1, 4, 4, -8, -2, -9, 8,
    -- layer=1 filter=47 channel=86
    1, -7, 9, -11, 0, -7, -5, 2, -11,
    -- layer=1 filter=47 channel=87
    3, 4, -2, 0, 7, 3, 7, 4, 2,
    -- layer=1 filter=47 channel=88
    -6, 6, -4, 0, 0, -5, -4, -5, 4,
    -- layer=1 filter=47 channel=89
    -2, -9, -9, -11, 5, 0, 2, 1, -2,
    -- layer=1 filter=47 channel=90
    -5, -1, 4, -9, 9, -10, 1, -4, 9,
    -- layer=1 filter=47 channel=91
    -6, -7, 6, 0, -9, 8, -4, -8, 7,
    -- layer=1 filter=47 channel=92
    0, 3, 7, -5, 3, 7, 9, -5, 4,
    -- layer=1 filter=47 channel=93
    -6, -8, 7, 0, 6, 5, -2, 1, -8,
    -- layer=1 filter=47 channel=94
    -5, 1, -11, 5, 0, 1, 4, 6, -3,
    -- layer=1 filter=47 channel=95
    -6, 5, 3, -2, -10, 4, 0, -1, 0,
    -- layer=1 filter=47 channel=96
    -6, -4, 2, 7, 2, -6, 0, 5, 3,
    -- layer=1 filter=47 channel=97
    1, 2, 6, -8, 6, -2, -10, 6, 2,
    -- layer=1 filter=47 channel=98
    -10, -6, 3, 5, 3, -13, -13, 1, -6,
    -- layer=1 filter=47 channel=99
    -9, 8, 0, 1, 2, 6, 8, -11, -9,
    -- layer=1 filter=47 channel=100
    4, 3, 3, -6, 7, -7, 2, 5, 9,
    -- layer=1 filter=47 channel=101
    0, -6, 3, 0, -11, -6, -7, 8, -3,
    -- layer=1 filter=47 channel=102
    -6, -6, -7, -3, -9, 0, -4, -9, -7,
    -- layer=1 filter=47 channel=103
    2, 0, 5, 5, 3, 0, 5, -6, -7,
    -- layer=1 filter=47 channel=104
    -7, -1, 0, 9, 8, -5, -9, 5, -9,
    -- layer=1 filter=47 channel=105
    6, 4, -6, 1, 0, 6, -7, -6, -4,
    -- layer=1 filter=47 channel=106
    -6, -13, 5, -12, -8, 7, -6, 0, -3,
    -- layer=1 filter=47 channel=107
    -2, 0, 1, -10, 4, 5, -4, -7, -2,
    -- layer=1 filter=47 channel=108
    -6, 5, -9, -11, 4, -4, 10, -8, 1,
    -- layer=1 filter=47 channel=109
    4, 6, -3, -10, -2, 7, 0, -9, -2,
    -- layer=1 filter=47 channel=110
    -10, -10, -7, -10, -2, -4, 7, 0, -8,
    -- layer=1 filter=47 channel=111
    0, 4, 8, -3, -4, -13, -6, -9, -10,
    -- layer=1 filter=47 channel=112
    1, 6, 8, -1, -1, -1, -8, -6, -9,
    -- layer=1 filter=47 channel=113
    -4, -5, -2, -7, -4, 0, 1, -4, -8,
    -- layer=1 filter=47 channel=114
    2, -2, -2, -6, -1, 8, -1, -3, -10,
    -- layer=1 filter=47 channel=115
    8, 2, 6, -10, -1, -9, 0, 0, 0,
    -- layer=1 filter=47 channel=116
    6, -8, -3, 8, -9, -10, 0, 8, -5,
    -- layer=1 filter=47 channel=117
    9, -9, -7, -9, -1, -2, 0, -2, -2,
    -- layer=1 filter=47 channel=118
    -3, -6, 2, -6, 5, -4, 5, 0, -6,
    -- layer=1 filter=47 channel=119
    -8, 2, 3, 7, 7, -6, -6, 7, 2,
    -- layer=1 filter=47 channel=120
    -11, 6, -6, -9, -7, -2, 5, -7, -2,
    -- layer=1 filter=47 channel=121
    -3, -10, 0, 5, -11, 0, 0, -2, 3,
    -- layer=1 filter=47 channel=122
    -1, 5, 10, -3, -1, -3, -6, -1, 2,
    -- layer=1 filter=47 channel=123
    -3, -6, -7, -6, -1, 0, 0, -1, -10,
    -- layer=1 filter=47 channel=124
    5, -9, -3, -5, 8, 8, -4, 8, 7,
    -- layer=1 filter=47 channel=125
    5, 3, -3, -4, -10, -4, 5, -8, -3,
    -- layer=1 filter=47 channel=126
    -5, 0, 7, 9, -9, -10, -7, 10, 8,
    -- layer=1 filter=47 channel=127
    5, 1, -10, 8, 4, 1, 3, 5, -8,
    -- layer=1 filter=48 channel=0
    -8, -2, 2, -1, 2, -6, -4, 0, 5,
    -- layer=1 filter=48 channel=1
    -3, 3, 0, -7, 1, -3, 0, -7, 3,
    -- layer=1 filter=48 channel=2
    4, 7, -8, -3, -8, 3, -8, 0, 1,
    -- layer=1 filter=48 channel=3
    10, -8, 4, -7, -7, -7, -2, 6, 1,
    -- layer=1 filter=48 channel=4
    8, -3, -8, -6, -4, -2, 2, 4, 5,
    -- layer=1 filter=48 channel=5
    7, 0, 6, 4, 5, -3, 6, -6, 3,
    -- layer=1 filter=48 channel=6
    2, 4, -3, -9, -11, 0, -1, -3, -9,
    -- layer=1 filter=48 channel=7
    -10, -8, 0, -7, 1, -10, -10, 0, 3,
    -- layer=1 filter=48 channel=8
    -2, -4, -5, 4, -2, 3, -1, -2, -1,
    -- layer=1 filter=48 channel=9
    -10, -11, -6, 6, -3, -4, 4, 6, -5,
    -- layer=1 filter=48 channel=10
    0, 6, -11, -5, 1, 4, 6, 5, 1,
    -- layer=1 filter=48 channel=11
    2, -3, -6, 5, 6, -2, 7, 0, -10,
    -- layer=1 filter=48 channel=12
    -6, 4, -10, 7, -8, -5, 2, 6, 9,
    -- layer=1 filter=48 channel=13
    2, -2, -9, 8, -9, -10, 1, -11, -8,
    -- layer=1 filter=48 channel=14
    5, 4, 2, -11, 6, 4, 3, 7, -4,
    -- layer=1 filter=48 channel=15
    2, -11, 0, -1, -3, -5, -12, -8, -2,
    -- layer=1 filter=48 channel=16
    8, 8, 8, 8, -9, 0, -12, -11, 1,
    -- layer=1 filter=48 channel=17
    7, 0, -5, -3, 3, -10, 0, 4, 0,
    -- layer=1 filter=48 channel=18
    9, -4, 5, -12, 4, -1, -3, 0, 1,
    -- layer=1 filter=48 channel=19
    -2, -8, 0, 0, 0, 2, 0, -6, 7,
    -- layer=1 filter=48 channel=20
    -12, -3, 2, 3, -7, -10, 5, 8, 5,
    -- layer=1 filter=48 channel=21
    -5, 7, -11, 4, 1, 7, 6, -3, 5,
    -- layer=1 filter=48 channel=22
    -1, 5, 5, 6, -1, -5, 0, 8, 3,
    -- layer=1 filter=48 channel=23
    -7, 0, -6, 2, 0, 0, -1, 8, 7,
    -- layer=1 filter=48 channel=24
    -11, -1, -8, 1, 6, 1, 0, 4, -1,
    -- layer=1 filter=48 channel=25
    3, 8, -6, -10, -12, -6, 4, -10, -10,
    -- layer=1 filter=48 channel=26
    4, 0, -11, -9, 5, -1, -9, 0, -7,
    -- layer=1 filter=48 channel=27
    5, 9, -7, -6, -8, -10, -2, 0, -1,
    -- layer=1 filter=48 channel=28
    1, 0, 7, 7, 1, -1, -9, 8, -2,
    -- layer=1 filter=48 channel=29
    1, 0, -10, -7, -5, -11, 9, -3, -6,
    -- layer=1 filter=48 channel=30
    3, 0, -7, 0, 7, 8, 0, 0, 3,
    -- layer=1 filter=48 channel=31
    0, 0, -1, 0, -11, 5, -1, 4, 9,
    -- layer=1 filter=48 channel=32
    3, 3, -3, -5, 2, -3, -4, 2, -11,
    -- layer=1 filter=48 channel=33
    5, -11, 9, 5, 8, 2, 7, -10, 7,
    -- layer=1 filter=48 channel=34
    2, -3, -6, -2, 1, -11, 4, -5, 7,
    -- layer=1 filter=48 channel=35
    -7, -5, 0, -4, -10, -10, 7, 6, 9,
    -- layer=1 filter=48 channel=36
    -7, 0, -3, -9, 0, 4, -2, 6, -5,
    -- layer=1 filter=48 channel=37
    0, -5, -6, 3, 3, -6, 3, -5, -12,
    -- layer=1 filter=48 channel=38
    0, -13, -8, 2, -11, -6, 0, -5, 0,
    -- layer=1 filter=48 channel=39
    6, -11, -5, 3, -2, -4, 2, 1, 3,
    -- layer=1 filter=48 channel=40
    -16, 1, -3, -3, -8, -8, 0, 4, -3,
    -- layer=1 filter=48 channel=41
    0, 0, -3, 0, -4, -11, -2, -9, 8,
    -- layer=1 filter=48 channel=42
    7, -2, 2, -2, -10, -8, 7, -2, 7,
    -- layer=1 filter=48 channel=43
    -11, 0, -9, -6, -1, -6, -6, -7, 5,
    -- layer=1 filter=48 channel=44
    -10, 6, -4, 0, -9, -8, 2, 7, -8,
    -- layer=1 filter=48 channel=45
    -9, 4, -9, -10, -9, -3, 8, 1, -9,
    -- layer=1 filter=48 channel=46
    5, -6, 0, 5, 4, -9, 1, -9, 0,
    -- layer=1 filter=48 channel=47
    7, -11, -4, 3, -6, -1, -10, 6, -4,
    -- layer=1 filter=48 channel=48
    8, -11, -3, -8, -8, 6, 1, 2, -1,
    -- layer=1 filter=48 channel=49
    -8, -6, -4, 6, -10, -1, 0, -4, -5,
    -- layer=1 filter=48 channel=50
    -3, 7, -5, 6, -2, 4, -10, 2, 1,
    -- layer=1 filter=48 channel=51
    -3, 3, 2, -3, 1, -4, 8, -3, 5,
    -- layer=1 filter=48 channel=52
    -2, 9, 0, 0, 0, -10, 0, -6, 5,
    -- layer=1 filter=48 channel=53
    0, 6, -5, -2, -7, -12, 5, 5, -6,
    -- layer=1 filter=48 channel=54
    8, 3, 0, 3, 0, 7, 0, 0, -6,
    -- layer=1 filter=48 channel=55
    6, -7, -5, 9, 4, -6, -5, -12, 2,
    -- layer=1 filter=48 channel=56
    0, 1, -6, -7, -9, 1, 4, -6, -2,
    -- layer=1 filter=48 channel=57
    -1, -4, 0, 2, -6, -11, 5, 3, -1,
    -- layer=1 filter=48 channel=58
    7, -8, -10, -3, -7, 2, -2, -9, -1,
    -- layer=1 filter=48 channel=59
    -10, -10, -1, -10, 5, -8, 5, 7, -2,
    -- layer=1 filter=48 channel=60
    0, 9, 9, 5, 9, 6, -4, 4, 0,
    -- layer=1 filter=48 channel=61
    3, -10, 3, 7, 6, -3, 3, -8, -3,
    -- layer=1 filter=48 channel=62
    7, 5, -2, 7, -7, 3, 0, -8, -5,
    -- layer=1 filter=48 channel=63
    -4, 3, 6, -11, -4, 5, 3, 5, -8,
    -- layer=1 filter=48 channel=64
    0, -10, -7, -7, -10, 7, -4, -11, -1,
    -- layer=1 filter=48 channel=65
    7, -7, -11, 2, 5, 4, 4, 3, 0,
    -- layer=1 filter=48 channel=66
    -11, 3, -10, -5, 0, -5, -7, 9, -11,
    -- layer=1 filter=48 channel=67
    -5, 7, 8, -5, -2, 0, 2, 4, 8,
    -- layer=1 filter=48 channel=68
    7, -10, 4, 6, -1, -7, -5, 4, -8,
    -- layer=1 filter=48 channel=69
    -6, 1, 0, -6, 0, 9, 3, -10, -7,
    -- layer=1 filter=48 channel=70
    -11, 1, -9, 1, 1, 6, -4, 0, 2,
    -- layer=1 filter=48 channel=71
    3, -7, 7, 8, -11, 8, -9, 8, 1,
    -- layer=1 filter=48 channel=72
    -2, 1, -4, 5, -1, -7, 1, -5, -5,
    -- layer=1 filter=48 channel=73
    -4, 1, -1, 1, 0, -6, -5, 7, -10,
    -- layer=1 filter=48 channel=74
    0, 2, -8, 8, 5, -2, -9, 4, 0,
    -- layer=1 filter=48 channel=75
    6, 8, -4, -5, 4, 8, 3, 3, -10,
    -- layer=1 filter=48 channel=76
    8, -11, -9, -11, 0, -3, 1, 8, -6,
    -- layer=1 filter=48 channel=77
    -5, 0, 1, -11, -5, 7, 0, -11, -10,
    -- layer=1 filter=48 channel=78
    -5, -5, -9, 0, -7, -1, -7, 0, -8,
    -- layer=1 filter=48 channel=79
    -6, -5, -1, 2, -8, -9, -5, 5, 5,
    -- layer=1 filter=48 channel=80
    9, 0, 9, 7, -6, -6, 4, 9, 2,
    -- layer=1 filter=48 channel=81
    8, -10, -6, -9, 8, 0, 9, 1, -11,
    -- layer=1 filter=48 channel=82
    -9, 0, 1, 1, -4, -1, -5, 3, -4,
    -- layer=1 filter=48 channel=83
    -10, 8, -10, 0, -11, 4, 7, -3, -1,
    -- layer=1 filter=48 channel=84
    -1, -8, 8, -8, -4, -5, -8, 6, 7,
    -- layer=1 filter=48 channel=85
    -9, -9, -7, -10, -9, -9, 1, 7, 5,
    -- layer=1 filter=48 channel=86
    -12, 9, 7, -1, -4, 1, 7, 4, -8,
    -- layer=1 filter=48 channel=87
    -3, -4, 0, -2, -11, -4, 4, -6, 6,
    -- layer=1 filter=48 channel=88
    8, 8, -5, 10, -2, 0, 0, 11, 1,
    -- layer=1 filter=48 channel=89
    -3, -7, 5, -5, -5, -3, -8, 8, -9,
    -- layer=1 filter=48 channel=90
    -1, 3, 4, 2, 0, -7, -3, -7, -9,
    -- layer=1 filter=48 channel=91
    6, 8, 5, 4, -6, 0, 7, 1, 8,
    -- layer=1 filter=48 channel=92
    2, -4, 8, 1, 0, 3, -5, 3, -5,
    -- layer=1 filter=48 channel=93
    -6, -10, -6, -2, 7, 3, 2, -2, 4,
    -- layer=1 filter=48 channel=94
    -5, 7, -4, 7, -8, 5, 8, 3, -5,
    -- layer=1 filter=48 channel=95
    -9, -2, -3, -7, 5, -9, -5, -7, -1,
    -- layer=1 filter=48 channel=96
    -1, 6, -11, -8, 2, -10, -4, 0, -10,
    -- layer=1 filter=48 channel=97
    1, 6, -10, -1, 2, -11, -9, 1, 3,
    -- layer=1 filter=48 channel=98
    0, 4, -6, -6, 5, 6, 8, 2, 0,
    -- layer=1 filter=48 channel=99
    -11, -6, 8, 2, -10, 3, 1, 6, -6,
    -- layer=1 filter=48 channel=100
    -1, 3, 3, 8, 3, 6, 5, 2, 8,
    -- layer=1 filter=48 channel=101
    0, 5, -3, 0, -6, -3, 8, -4, -1,
    -- layer=1 filter=48 channel=102
    5, -11, 3, 3, -4, -8, -9, -8, 2,
    -- layer=1 filter=48 channel=103
    8, -9, -1, 1, 4, 7, -10, -8, -1,
    -- layer=1 filter=48 channel=104
    6, -9, -8, 1, 5, 0, 6, -3, 4,
    -- layer=1 filter=48 channel=105
    1, 3, -6, -10, -2, -11, 7, -6, -4,
    -- layer=1 filter=48 channel=106
    5, -11, 0, 0, 8, -5, -1, -11, -5,
    -- layer=1 filter=48 channel=107
    7, 0, -8, 5, 1, -9, 3, -10, -8,
    -- layer=1 filter=48 channel=108
    -9, -7, 8, 4, -3, 3, 5, -6, 2,
    -- layer=1 filter=48 channel=109
    3, -9, 1, -2, 8, 1, -9, -3, 6,
    -- layer=1 filter=48 channel=110
    3, -11, -9, 3, -6, 3, 0, -7, 2,
    -- layer=1 filter=48 channel=111
    3, -5, 0, -5, 8, 3, 10, 3, 5,
    -- layer=1 filter=48 channel=112
    3, -7, 7, 7, -1, -3, 1, -4, 0,
    -- layer=1 filter=48 channel=113
    -12, -1, -1, 0, -8, -7, 2, -8, 4,
    -- layer=1 filter=48 channel=114
    -6, 0, -11, 1, -9, 7, -4, 0, 0,
    -- layer=1 filter=48 channel=115
    -9, 3, 0, -2, -1, 0, 4, 0, -10,
    -- layer=1 filter=48 channel=116
    -2, -6, -1, -2, 0, 5, -10, -8, -2,
    -- layer=1 filter=48 channel=117
    6, 2, 7, 0, 1, -4, 0, -7, -6,
    -- layer=1 filter=48 channel=118
    0, -8, -10, 0, -10, 5, 1, -6, -3,
    -- layer=1 filter=48 channel=119
    -8, 8, 0, -7, -11, -7, -3, -3, -6,
    -- layer=1 filter=48 channel=120
    -11, 6, -6, -1, 4, 0, -1, -3, -4,
    -- layer=1 filter=48 channel=121
    7, -13, 0, -9, 6, -2, 0, -8, -10,
    -- layer=1 filter=48 channel=122
    -3, 8, 8, -2, -7, 1, 0, 6, -9,
    -- layer=1 filter=48 channel=123
    -1, -9, -4, -5, 8, 0, 1, -9, -3,
    -- layer=1 filter=48 channel=124
    5, -4, -7, 0, -6, -10, 1, -8, 5,
    -- layer=1 filter=48 channel=125
    2, 2, -3, -14, 7, 1, 1, 8, -9,
    -- layer=1 filter=48 channel=126
    0, 3, 3, -8, -3, -5, 5, 5, 2,
    -- layer=1 filter=48 channel=127
    8, -6, 0, -3, -8, -8, -3, 7, -2,
    -- layer=1 filter=49 channel=0
    -8, -21, -20, -9, -9, 4, -31, 0, -1,
    -- layer=1 filter=49 channel=1
    24, 33, -14, 13, -6, 11, 0, -23, -24,
    -- layer=1 filter=49 channel=2
    -3, 40, 20, 17, 23, 12, 21, 24, 7,
    -- layer=1 filter=49 channel=3
    -1, 10, 6, -7, -1, 0, 9, 0, 6,
    -- layer=1 filter=49 channel=4
    0, -10, -22, 10, 0, -9, 0, 1, 2,
    -- layer=1 filter=49 channel=5
    35, 42, 22, -4, 21, 45, 16, -7, 9,
    -- layer=1 filter=49 channel=6
    33, 51, 22, 8, -8, -8, 19, -60, -4,
    -- layer=1 filter=49 channel=7
    76, 24, 21, 39, -34, 7, -12, -1, 25,
    -- layer=1 filter=49 channel=8
    7, 16, -33, -31, 10, 22, -10, -13, 0,
    -- layer=1 filter=49 channel=9
    5, 11, -45, -7, 6, -15, 17, 8, -15,
    -- layer=1 filter=49 channel=10
    79, 19, 35, 38, -24, 13, -14, -11, 12,
    -- layer=1 filter=49 channel=11
    5, 13, -7, 31, 36, 30, 4, 33, 44,
    -- layer=1 filter=49 channel=12
    -11, 41, 30, -32, 23, 12, 28, 17, -56,
    -- layer=1 filter=49 channel=13
    -22, -14, -43, -48, -53, -54, -12, -53, -48,
    -- layer=1 filter=49 channel=14
    18, 16, 34, 24, -15, 13, -10, -5, 15,
    -- layer=1 filter=49 channel=15
    25, 3, 48, -16, 1, 46, -19, -43, -40,
    -- layer=1 filter=49 channel=16
    -11, -10, -42, -16, -7, 3, 7, 0, 13,
    -- layer=1 filter=49 channel=17
    -21, -21, -24, -18, 14, -8, -12, -17, -5,
    -- layer=1 filter=49 channel=18
    16, 18, 12, 32, 36, 3, 9, 18, 40,
    -- layer=1 filter=49 channel=19
    -11, 4, 11, -34, -24, -25, 8, 24, -6,
    -- layer=1 filter=49 channel=20
    -41, -47, -28, -77, -87, -63, -19, -56, -50,
    -- layer=1 filter=49 channel=21
    7, 29, 15, 5, -15, 0, 1, -13, -22,
    -- layer=1 filter=49 channel=22
    -32, -52, -43, 6, -7, -11, 5, -29, -21,
    -- layer=1 filter=49 channel=23
    6, -9, 22, -17, -11, 10, 30, -7, 32,
    -- layer=1 filter=49 channel=24
    2, 30, -17, -22, 13, 6, -8, -14, 3,
    -- layer=1 filter=49 channel=25
    68, 6, 2, 16, -34, -5, -20, 14, 38,
    -- layer=1 filter=49 channel=26
    19, 17, -23, -1, 23, 12, 24, -4, 17,
    -- layer=1 filter=49 channel=27
    19, 38, 13, 51, 73, 62, 36, 50, 39,
    -- layer=1 filter=49 channel=28
    47, -6, 10, 50, -16, 11, -3, -1, 8,
    -- layer=1 filter=49 channel=29
    -6, 12, -3, 7, 14, 9, -1, 18, 14,
    -- layer=1 filter=49 channel=30
    8, 5, 2, -31, -3, -54, -21, -20, -9,
    -- layer=1 filter=49 channel=31
    16, 45, 36, -18, 10, -6, 5, -16, 14,
    -- layer=1 filter=49 channel=32
    36, 12, 16, 14, -5, 10, 29, -19, -27,
    -- layer=1 filter=49 channel=33
    9, -10, 5, 8, 14, 10, 19, 20, 9,
    -- layer=1 filter=49 channel=34
    -3, 4, -22, 3, -17, -13, 1, -2, -10,
    -- layer=1 filter=49 channel=35
    14, 17, 8, 9, 5, 6, 16, 6, 10,
    -- layer=1 filter=49 channel=36
    2, -5, -2, 22, 40, 43, 4, 26, 39,
    -- layer=1 filter=49 channel=37
    47, 37, 13, -4, 17, 29, 3, 0, 16,
    -- layer=1 filter=49 channel=38
    -21, 3, -5, -56, -95, -71, -27, -56, -29,
    -- layer=1 filter=49 channel=39
    -21, -24, -22, -5, 6, 13, -1, 16, 20,
    -- layer=1 filter=49 channel=40
    -23, 7, -1, -11, -26, -31, 6, -23, 7,
    -- layer=1 filter=49 channel=41
    50, 18, 2, 30, 27, 1, 24, -4, -11,
    -- layer=1 filter=49 channel=42
    -21, 0, 9, -9, 3, 3, 5, 7, -7,
    -- layer=1 filter=49 channel=43
    34, 2, -34, -16, -21, 21, -6, -18, 3,
    -- layer=1 filter=49 channel=44
    25, 35, 4, 2, 20, 21, 23, -6, -19,
    -- layer=1 filter=49 channel=45
    -14, -1, -4, -38, -4, 14, -4, -38, -33,
    -- layer=1 filter=49 channel=46
    -19, 4, 29, -10, -42, 10, 19, 53, -25,
    -- layer=1 filter=49 channel=47
    18, 7, 50, 17, 13, -24, 45, -31, -7,
    -- layer=1 filter=49 channel=48
    26, 7, 24, -31, -14, -27, -21, -27, 4,
    -- layer=1 filter=49 channel=49
    -4, -14, -6, -17, -15, -27, -12, -9, 3,
    -- layer=1 filter=49 channel=50
    25, -9, 11, 5, 2, 6, 35, 9, 2,
    -- layer=1 filter=49 channel=51
    39, -6, 3, -18, -98, -23, -45, -66, -6,
    -- layer=1 filter=49 channel=52
    14, -11, -17, 15, -14, -31, -5, -22, -9,
    -- layer=1 filter=49 channel=53
    7, -12, 19, 1, 10, 13, 6, 0, 14,
    -- layer=1 filter=49 channel=54
    81, 10, 19, -3, -12, 11, 1, 26, 46,
    -- layer=1 filter=49 channel=55
    12, 18, 4, 44, 68, 48, 32, 43, 28,
    -- layer=1 filter=49 channel=56
    -8, -3, 6, -8, 7, 2, 2, -9, 1,
    -- layer=1 filter=49 channel=57
    37, -24, 13, 16, -36, -15, -28, -39, 10,
    -- layer=1 filter=49 channel=58
    43, -4, 8, -3, 12, -2, 24, -11, 37,
    -- layer=1 filter=49 channel=59
    -4, 8, 2, -1, -1, 9, -8, -1, 11,
    -- layer=1 filter=49 channel=60
    -25, -2, -17, 2, -14, 2, -29, -29, -11,
    -- layer=1 filter=49 channel=61
    -11, -2, 7, 1, -6, -9, 2, 8, 4,
    -- layer=1 filter=49 channel=62
    18, 12, -26, -35, -4, 21, -11, -23, 15,
    -- layer=1 filter=49 channel=63
    6, -1, -4, 36, 19, 10, 3, 18, 15,
    -- layer=1 filter=49 channel=64
    -11, 6, -15, 5, -10, 12, -1, -10, -21,
    -- layer=1 filter=49 channel=65
    4, 27, 6, -18, -12, 0, 12, -7, 19,
    -- layer=1 filter=49 channel=66
    -3, 1, -14, 4, 11, 16, -3, -3, -4,
    -- layer=1 filter=49 channel=67
    74, 70, 64, 16, -25, 27, 7, -15, 25,
    -- layer=1 filter=49 channel=68
    51, 38, 0, 19, 14, 30, 11, 16, -7,
    -- layer=1 filter=49 channel=69
    -2, 0, -30, -26, 8, 26, 12, 3, -3,
    -- layer=1 filter=49 channel=70
    50, 103, 75, -23, 26, 30, 27, -20, 8,
    -- layer=1 filter=49 channel=71
    11, 2, 3, -23, -21, 8, 5, 10, -4,
    -- layer=1 filter=49 channel=72
    13, 6, 16, 17, 24, 8, 45, 13, 0,
    -- layer=1 filter=49 channel=73
    -2, 4, 9, 7, -1, 0, 0, 7, 11,
    -- layer=1 filter=49 channel=74
    11, 38, -27, -13, -34, 12, -41, -15, -11,
    -- layer=1 filter=49 channel=75
    -2, 20, 19, -9, -34, -30, 1, 7, -29,
    -- layer=1 filter=49 channel=76
    24, -8, -20, -3, -1, -37, -20, -9, -23,
    -- layer=1 filter=49 channel=77
    35, 45, 11, 15, -15, -2, -8, -12, -11,
    -- layer=1 filter=49 channel=78
    16, 6, 6, 25, 0, -7, -3, 7, 11,
    -- layer=1 filter=49 channel=79
    -7, -15, -34, -41, -3, -8, -10, -23, 0,
    -- layer=1 filter=49 channel=80
    2, -9, -1, -9, 3, -3, 0, 0, 3,
    -- layer=1 filter=49 channel=81
    6, -8, -8, -5, 12, 2, -6, 1, -3,
    -- layer=1 filter=49 channel=82
    8, 17, 37, -29, -41, -14, 1, -40, -18,
    -- layer=1 filter=49 channel=83
    -1, -2, 16, -25, 11, 15, -5, -40, -26,
    -- layer=1 filter=49 channel=84
    6, 4, -4, 27, 12, -7, -4, 24, 35,
    -- layer=1 filter=49 channel=85
    19, -17, 23, -6, 5, -7, 26, -1, -21,
    -- layer=1 filter=49 channel=86
    0, -2, -9, 12, 13, 26, 7, 3, 14,
    -- layer=1 filter=49 channel=87
    -23, 31, 7, -30, 14, -23, 28, 18, -29,
    -- layer=1 filter=49 channel=88
    20, 4, 23, 10, 13, 12, 21, 24, 41,
    -- layer=1 filter=49 channel=89
    -19, 17, 29, -12, -42, -6, -8, -2, -34,
    -- layer=1 filter=49 channel=90
    18, 35, -27, -19, 11, 34, 8, -24, -24,
    -- layer=1 filter=49 channel=91
    -11, -9, -8, -38, -78, -76, -19, -80, -58,
    -- layer=1 filter=49 channel=92
    68, 18, 13, 22, 31, -4, 30, 0, -30,
    -- layer=1 filter=49 channel=93
    -33, -26, -25, -50, -46, -20, -32, -47, -38,
    -- layer=1 filter=49 channel=94
    -15, -31, -23, -5, -22, -6, -26, -2, 0,
    -- layer=1 filter=49 channel=95
    -5, 11, -8, 4, -17, -11, -24, 22, 21,
    -- layer=1 filter=49 channel=96
    10, 4, 16, 13, 18, 3, 4, 29, 19,
    -- layer=1 filter=49 channel=97
    -27, -27, -24, -25, -24, -7, -23, -16, -21,
    -- layer=1 filter=49 channel=98
    9, -21, -51, -5, 2, 22, -29, -40, -15,
    -- layer=1 filter=49 channel=99
    21, -18, 37, 30, -47, 15, -31, -15, 37,
    -- layer=1 filter=49 channel=100
    7, 22, 19, 37, 27, 34, 7, 26, 31,
    -- layer=1 filter=49 channel=101
    -34, -4, -8, -75, -110, -88, -54, -67, -58,
    -- layer=1 filter=49 channel=102
    -1, -21, -20, -41, -55, -43, -35, -49, -35,
    -- layer=1 filter=49 channel=103
    11, 22, 21, 10, 50, 38, 18, 29, 26,
    -- layer=1 filter=49 channel=104
    -23, -11, 42, -32, -5, -20, 22, -25, 2,
    -- layer=1 filter=49 channel=105
    -18, -33, -30, -3, -1, -11, -24, -27, -3,
    -- layer=1 filter=49 channel=106
    -3, 0, -10, -29, -59, -40, -21, -45, -64,
    -- layer=1 filter=49 channel=107
    0, 17, 10, 1, 4, 2, 9, -4, 0,
    -- layer=1 filter=49 channel=108
    45, 35, 29, 7, 35, 27, 37, -16, -1,
    -- layer=1 filter=49 channel=109
    0, -2, 5, 0, 0, -11, -6, 1, 8,
    -- layer=1 filter=49 channel=110
    6, -10, 0, 0, -13, -7, -20, -23, -7,
    -- layer=1 filter=49 channel=111
    5, -1, 5, 1, -12, -20, -38, -13, 12,
    -- layer=1 filter=49 channel=112
    11, 23, 22, 14, -8, 2, -16, 5, 22,
    -- layer=1 filter=49 channel=113
    -29, -37, -5, -23, -22, -5, -33, -10, -18,
    -- layer=1 filter=49 channel=114
    4, 18, 6, -6, 41, 47, 50, 26, 20,
    -- layer=1 filter=49 channel=115
    -23, -33, -14, -13, 4, 1, -30, 7, 5,
    -- layer=1 filter=49 channel=116
    2, -7, -10, -10, 2, -4, -2, 0, 0,
    -- layer=1 filter=49 channel=117
    3, 0, 25, 5, -6, -47, -9, -18, 47,
    -- layer=1 filter=49 channel=118
    11, 10, -1, -34, -23, -37, -32, 2, -1,
    -- layer=1 filter=49 channel=119
    49, 43, 0, 6, 12, 15, 27, -29, -8,
    -- layer=1 filter=49 channel=120
    49, 21, -15, -7, -26, -33, -16, -27, 0,
    -- layer=1 filter=49 channel=121
    16, 65, 43, 10, 32, 32, 20, 49, 42,
    -- layer=1 filter=49 channel=122
    4, 8, -9, 2, 4, -9, 0, 0, -3,
    -- layer=1 filter=49 channel=123
    3, 20, 21, 24, 54, 37, 14, 43, 35,
    -- layer=1 filter=49 channel=124
    6, 19, 9, 10, 5, 6, 2, 7, 3,
    -- layer=1 filter=49 channel=125
    70, 92, 104, 25, 11, -22, 10, -38, 39,
    -- layer=1 filter=49 channel=126
    21, 55, -11, 25, 29, 29, -19, -43, -13,
    -- layer=1 filter=49 channel=127
    13, 9, 6, -18, -25, -20, -20, -3, -9,
    -- layer=1 filter=50 channel=0
    -2, 0, 4, -7, -14, -7, -6, 0, -9,
    -- layer=1 filter=50 channel=1
    -10, 2, 1, -2, 3, -11, 8, -7, 8,
    -- layer=1 filter=50 channel=2
    -27, -18, -18, -10, -21, -14, -2, -4, -11,
    -- layer=1 filter=50 channel=3
    -10, -1, -7, -1, 8, -6, -3, -10, 0,
    -- layer=1 filter=50 channel=4
    1, -9, -7, -4, -5, -4, 5, 4, 3,
    -- layer=1 filter=50 channel=5
    -7, -6, -7, 3, -17, -3, -19, -9, -11,
    -- layer=1 filter=50 channel=6
    2, -7, -2, 2, -8, 0, 4, -13, -4,
    -- layer=1 filter=50 channel=7
    -6, 1, 1, 1, -8, -7, -18, 1, 13,
    -- layer=1 filter=50 channel=8
    -2, -4, -11, -5, -17, -8, -4, 4, 5,
    -- layer=1 filter=50 channel=9
    0, 6, 0, -12, -13, 4, 0, -5, -2,
    -- layer=1 filter=50 channel=10
    -6, 4, -14, -17, -4, -9, -11, -2, -3,
    -- layer=1 filter=50 channel=11
    -6, -16, -1, -1, 0, -17, -5, -2, 0,
    -- layer=1 filter=50 channel=12
    3, -6, 7, -3, 7, 4, 9, 0, 4,
    -- layer=1 filter=50 channel=13
    3, -16, -2, -15, -16, -8, -19, -3, -13,
    -- layer=1 filter=50 channel=14
    -18, 4, -21, -14, -5, -3, -7, -3, -8,
    -- layer=1 filter=50 channel=15
    -13, 5, -2, -7, 0, -15, 0, -8, -1,
    -- layer=1 filter=50 channel=16
    -11, -13, -12, -8, -9, 0, 0, 4, -7,
    -- layer=1 filter=50 channel=17
    7, 5, -1, 0, 6, 6, -12, -10, -6,
    -- layer=1 filter=50 channel=18
    0, -5, -19, 1, -13, -9, 1, 0, -13,
    -- layer=1 filter=50 channel=19
    -6, -1, 4, -3, -6, 5, -6, -8, -8,
    -- layer=1 filter=50 channel=20
    -4, -12, 2, -8, -1, -8, 0, 0, -1,
    -- layer=1 filter=50 channel=21
    -7, -3, -14, -8, 4, -1, -12, -8, -1,
    -- layer=1 filter=50 channel=22
    -3, -10, -6, 2, -9, -11, 2, -7, 2,
    -- layer=1 filter=50 channel=23
    -3, 10, 2, 8, 0, -4, 0, -9, -9,
    -- layer=1 filter=50 channel=24
    -7, -5, -15, -26, -11, -2, -18, -11, -23,
    -- layer=1 filter=50 channel=25
    3, -8, -4, -5, -7, -10, -12, -10, -16,
    -- layer=1 filter=50 channel=26
    -12, -1, 0, -4, -10, -13, -22, -16, 0,
    -- layer=1 filter=50 channel=27
    5, 8, 0, -1, 8, -2, 5, 0, 1,
    -- layer=1 filter=50 channel=28
    1, -9, 6, 4, 3, 1, -2, -6, 6,
    -- layer=1 filter=50 channel=29
    -4, -6, 0, -12, 4, -3, 0, -9, -3,
    -- layer=1 filter=50 channel=30
    -10, -13, -20, -20, -23, -5, 15, 0, -12,
    -- layer=1 filter=50 channel=31
    -17, -20, -9, -13, -20, -15, -10, -23, -3,
    -- layer=1 filter=50 channel=32
    -14, -10, -12, -9, -3, -8, 7, -7, 2,
    -- layer=1 filter=50 channel=33
    -6, -15, -2, -9, -8, 0, -5, 3, 4,
    -- layer=1 filter=50 channel=34
    5, -9, 1, 1, 5, -10, 8, 5, -7,
    -- layer=1 filter=50 channel=35
    3, -7, -9, -8, -1, 1, 3, 4, 5,
    -- layer=1 filter=50 channel=36
    -7, 0, -16, -7, -17, -8, -4, -6, 2,
    -- layer=1 filter=50 channel=37
    -3, 11, 5, -8, 1, -1, -15, -11, 0,
    -- layer=1 filter=50 channel=38
    -10, 2, -9, -3, -16, -1, -11, -15, -17,
    -- layer=1 filter=50 channel=39
    -5, 3, -3, -8, -14, -15, -15, -13, -2,
    -- layer=1 filter=50 channel=40
    -7, -32, -5, -9, -18, -16, 3, -10, 7,
    -- layer=1 filter=50 channel=41
    -7, -16, -6, -13, -8, -14, -6, -8, -17,
    -- layer=1 filter=50 channel=42
    -6, -20, -18, -3, -4, -19, 5, -6, 0,
    -- layer=1 filter=50 channel=43
    3, 5, -4, 3, -10, -13, -7, -6, -5,
    -- layer=1 filter=50 channel=44
    3, 7, 4, -2, 2, -5, -7, 3, 7,
    -- layer=1 filter=50 channel=45
    0, 8, -7, -8, -9, -11, 0, 1, -11,
    -- layer=1 filter=50 channel=46
    2, -6, -2, 20, 17, -3, 2, -2, -11,
    -- layer=1 filter=50 channel=47
    3, -2, 2, -1, -7, -15, -1, 2, -12,
    -- layer=1 filter=50 channel=48
    -1, -12, -9, -3, -12, 4, -5, -1, 0,
    -- layer=1 filter=50 channel=49
    -8, 4, -5, -11, -5, 3, -13, 0, -4,
    -- layer=1 filter=50 channel=50
    -3, 3, -9, -10, 4, 8, -1, -1, 8,
    -- layer=1 filter=50 channel=51
    -10, -10, 0, -13, -9, -4, -2, 0, -2,
    -- layer=1 filter=50 channel=52
    -8, 3, 5, 9, -1, 3, -10, 8, 6,
    -- layer=1 filter=50 channel=53
    -3, -9, 7, 0, 7, -10, -1, 6, 10,
    -- layer=1 filter=50 channel=54
    3, -6, -8, -7, -3, 0, -20, 0, -10,
    -- layer=1 filter=50 channel=55
    -11, 0, 3, -15, -1, -11, -3, -6, -6,
    -- layer=1 filter=50 channel=56
    0, -2, -6, -5, 0, 3, 1, 7, -2,
    -- layer=1 filter=50 channel=57
    -13, 7, 0, -16, 0, -2, -3, 8, -3,
    -- layer=1 filter=50 channel=58
    -12, -10, -18, -12, -1, -14, -2, 0, 1,
    -- layer=1 filter=50 channel=59
    7, 0, 1, 3, -10, -9, 8, 10, 3,
    -- layer=1 filter=50 channel=60
    -7, 1, -6, 7, 1, -1, 7, -8, -6,
    -- layer=1 filter=50 channel=61
    4, -3, 7, -11, -4, -1, 0, -6, -4,
    -- layer=1 filter=50 channel=62
    12, 9, -2, 5, -3, 4, -2, -4, -9,
    -- layer=1 filter=50 channel=63
    -18, -16, -10, 1, -9, 0, -17, -1, -12,
    -- layer=1 filter=50 channel=64
    -3, -1, -5, 3, -4, -6, 6, 1, -8,
    -- layer=1 filter=50 channel=65
    -11, -2, 3, 1, -12, -3, -3, -6, -3,
    -- layer=1 filter=50 channel=66
    -6, -18, -7, -18, 0, -11, -2, -7, -11,
    -- layer=1 filter=50 channel=67
    3, 1, -13, -2, -2, 5, -12, -7, -16,
    -- layer=1 filter=50 channel=68
    -4, -3, 3, -7, -5, -7, -13, -4, -4,
    -- layer=1 filter=50 channel=69
    -14, -6, 6, -17, -20, 4, -1, -1, -12,
    -- layer=1 filter=50 channel=70
    -10, -6, -17, 7, -10, 0, -9, -4, -19,
    -- layer=1 filter=50 channel=71
    -10, -4, -21, -2, -16, -19, -15, -10, -9,
    -- layer=1 filter=50 channel=72
    -3, -2, 3, -5, -3, 6, -5, -9, -12,
    -- layer=1 filter=50 channel=73
    -9, -3, -3, 7, -1, 8, -10, 5, -4,
    -- layer=1 filter=50 channel=74
    6, 1, 0, 3, 5, 0, -9, 0, 3,
    -- layer=1 filter=50 channel=75
    1, -9, 0, -8, -9, 2, 12, 10, 6,
    -- layer=1 filter=50 channel=76
    -12, -2, -9, -8, 2, -14, 3, -8, -5,
    -- layer=1 filter=50 channel=77
    6, 0, 7, 8, 0, 2, -7, 9, 1,
    -- layer=1 filter=50 channel=78
    8, 1, -8, 0, -1, -5, 2, 7, 3,
    -- layer=1 filter=50 channel=79
    -13, -8, 4, -1, -15, 0, -13, -3, -8,
    -- layer=1 filter=50 channel=80
    -4, -7, 8, 2, 6, 2, 7, 2, -4,
    -- layer=1 filter=50 channel=81
    -3, -5, 0, -3, -7, 1, -1, -11, 3,
    -- layer=1 filter=50 channel=82
    0, -13, -12, 8, 3, 0, 0, 3, -4,
    -- layer=1 filter=50 channel=83
    -3, -7, -4, 4, -10, -3, -2, 6, -3,
    -- layer=1 filter=50 channel=84
    -9, -9, 0, -17, -8, -1, 6, 7, 0,
    -- layer=1 filter=50 channel=85
    -3, -4, 1, -8, -9, -10, 1, -7, -1,
    -- layer=1 filter=50 channel=86
    -11, -11, -6, -17, -3, -12, -21, -20, -14,
    -- layer=1 filter=50 channel=87
    5, -2, 0, 5, -4, -8, -7, -5, 8,
    -- layer=1 filter=50 channel=88
    5, -5, -17, 0, -8, -7, -12, -3, 0,
    -- layer=1 filter=50 channel=89
    1, -12, -7, -3, -12, 6, -1, -9, -7,
    -- layer=1 filter=50 channel=90
    1, 5, -12, -1, 7, 5, 1, -9, -5,
    -- layer=1 filter=50 channel=91
    2, -10, -14, 4, 0, -11, -4, -11, -10,
    -- layer=1 filter=50 channel=92
    -1, -4, 0, 0, -1, 5, -10, 5, -10,
    -- layer=1 filter=50 channel=93
    1, -14, -18, -9, -8, -4, -6, -12, -12,
    -- layer=1 filter=50 channel=94
    -2, -15, -9, -14, -15, -11, -12, -8, 0,
    -- layer=1 filter=50 channel=95
    -6, -17, -5, -17, 0, 2, -2, -2, 4,
    -- layer=1 filter=50 channel=96
    1, -7, 5, -7, -7, 7, -3, 5, 1,
    -- layer=1 filter=50 channel=97
    -6, -4, -13, -17, 1, -11, -5, -10, 1,
    -- layer=1 filter=50 channel=98
    -5, -2, -7, 0, -12, -1, 1, -12, 6,
    -- layer=1 filter=50 channel=99
    -2, -8, -8, 3, -9, -9, -9, 7, 1,
    -- layer=1 filter=50 channel=100
    -18, -15, -1, -1, -2, -18, -16, -9, -2,
    -- layer=1 filter=50 channel=101
    2, -3, -1, 3, 1, 1, -5, -3, 3,
    -- layer=1 filter=50 channel=102
    4, -1, -10, -7, 3, -10, -5, 3, 5,
    -- layer=1 filter=50 channel=103
    0, -15, -17, -3, -5, 0, -5, -6, -12,
    -- layer=1 filter=50 channel=104
    -3, -6, -6, 9, 5, -4, -2, 8, -6,
    -- layer=1 filter=50 channel=105
    -2, 0, -18, -11, -14, -3, -3, 2, 1,
    -- layer=1 filter=50 channel=106
    -14, -7, 6, -10, -13, 4, -15, -21, 1,
    -- layer=1 filter=50 channel=107
    -3, 1, 0, 2, 6, 0, 6, 0, 2,
    -- layer=1 filter=50 channel=108
    -7, -3, -2, -15, -4, 4, -25, -8, 0,
    -- layer=1 filter=50 channel=109
    -4, -5, 6, 3, 2, -11, 0, 0, 9,
    -- layer=1 filter=50 channel=110
    -4, -2, 7, 2, -8, -11, 8, -8, 5,
    -- layer=1 filter=50 channel=111
    -11, -17, -4, -8, -15, -21, -12, -11, 0,
    -- layer=1 filter=50 channel=112
    -3, 6, 7, 4, -2, 0, 0, 0, 2,
    -- layer=1 filter=50 channel=113
    5, -1, -7, -8, -7, 5, -5, -4, -13,
    -- layer=1 filter=50 channel=114
    5, 11, -5, 5, 0, -1, -3, -8, -1,
    -- layer=1 filter=50 channel=115
    1, -1, -6, -9, 2, -18, -19, -8, -3,
    -- layer=1 filter=50 channel=116
    -1, 4, -9, 1, 8, 7, -6, -8, 2,
    -- layer=1 filter=50 channel=117
    11, 3, -3, 0, -5, -7, -5, 4, -8,
    -- layer=1 filter=50 channel=118
    3, 7, -6, -9, 0, -12, 8, -10, -4,
    -- layer=1 filter=50 channel=119
    -5, -11, -10, -24, -14, -7, -22, -17, -5,
    -- layer=1 filter=50 channel=120
    -12, -2, -7, -2, -3, -12, -13, -10, -1,
    -- layer=1 filter=50 channel=121
    -2, -14, -15, -7, -1, -9, -1, -8, -17,
    -- layer=1 filter=50 channel=122
    -3, -7, -7, -4, -6, 10, 10, -1, -3,
    -- layer=1 filter=50 channel=123
    -4, -3, -7, -17, -4, 3, -5, -18, -20,
    -- layer=1 filter=50 channel=124
    -12, -14, 6, 0, 0, -7, -5, -10, 1,
    -- layer=1 filter=50 channel=125
    -1, -5, -5, -15, -4, -6, -10, -6, -8,
    -- layer=1 filter=50 channel=126
    -1, -6, -4, -6, 4, -8, -10, 0, 6,
    -- layer=1 filter=50 channel=127
    -2, -5, -17, -9, -4, -4, 16, 8, -1,
    -- layer=1 filter=51 channel=0
    0, 0, -25, 7, -6, -25, 14, 19, -9,
    -- layer=1 filter=51 channel=1
    -34, -8, -11, -25, -16, -4, 23, -19, 10,
    -- layer=1 filter=51 channel=2
    -5, -3, 11, 0, -1, 12, 28, 31, 49,
    -- layer=1 filter=51 channel=3
    5, 9, 10, 2, 5, 2, -5, 0, -7,
    -- layer=1 filter=51 channel=4
    -5, -4, 3, 0, 7, 6, 0, 4, 0,
    -- layer=1 filter=51 channel=5
    -12, 14, -8, -37, 3, 0, -4, -27, 2,
    -- layer=1 filter=51 channel=6
    12, 5, 39, -9, -49, 1, 33, -12, 42,
    -- layer=1 filter=51 channel=7
    29, -9, 5, 51, 15, 6, 56, 42, -10,
    -- layer=1 filter=51 channel=8
    -41, -11, -2, -32, 18, -5, -1, -6, 7,
    -- layer=1 filter=51 channel=9
    -15, 9, -18, -43, 1, -14, -9, 49, 17,
    -- layer=1 filter=51 channel=10
    22, 14, -3, 34, 38, -21, 42, 43, -27,
    -- layer=1 filter=51 channel=11
    4, 10, 0, 14, 23, 6, -2, 18, 1,
    -- layer=1 filter=51 channel=12
    -22, -37, 0, -20, -2, -27, 17, 45, 70,
    -- layer=1 filter=51 channel=13
    2, 2, 11, -24, -2, 10, 0, 0, 13,
    -- layer=1 filter=51 channel=14
    2, -39, 19, 5, 9, 0, -5, 37, 32,
    -- layer=1 filter=51 channel=15
    -29, 30, 28, -35, 21, 60, -26, 8, 22,
    -- layer=1 filter=51 channel=16
    -17, 10, -27, -13, -2, -15, 7, -22, 2,
    -- layer=1 filter=51 channel=17
    -18, -16, -11, -6, -5, -28, -10, 7, 36,
    -- layer=1 filter=51 channel=18
    23, -12, -7, -23, -23, -27, 5, -1, -17,
    -- layer=1 filter=51 channel=19
    -15, -61, -41, -60, -71, -114, -24, -69, -64,
    -- layer=1 filter=51 channel=20
    -16, -8, -9, -14, -44, -28, -3, -5, -6,
    -- layer=1 filter=51 channel=21
    -40, -34, -16, -13, -24, -11, 13, 11, 0,
    -- layer=1 filter=51 channel=22
    -30, -25, 7, 4, 8, -12, -4, 7, 22,
    -- layer=1 filter=51 channel=23
    15, 13, 28, 83, 18, 22, 53, 20, 31,
    -- layer=1 filter=51 channel=24
    -4, 19, 40, -20, 36, 7, -18, 20, 32,
    -- layer=1 filter=51 channel=25
    -8, -29, -74, 11, -45, -60, 47, 19, -45,
    -- layer=1 filter=51 channel=26
    0, 25, 18, -18, 41, 29, -40, 21, 35,
    -- layer=1 filter=51 channel=27
    26, 37, 31, 27, 25, 11, 25, 0, 10,
    -- layer=1 filter=51 channel=28
    3, -28, -24, 34, 29, -51, 55, 68, -37,
    -- layer=1 filter=51 channel=29
    0, 0, -2, -12, -1, -11, 1, -29, -1,
    -- layer=1 filter=51 channel=30
    15, -50, -29, -60, -64, -61, -35, -66, -28,
    -- layer=1 filter=51 channel=31
    20, -28, 10, -4, -38, -20, -22, -21, 11,
    -- layer=1 filter=51 channel=32
    -19, 50, 25, -25, 33, 30, -29, 44, 38,
    -- layer=1 filter=51 channel=33
    -3, 23, 30, 0, 15, 26, 10, 10, 11,
    -- layer=1 filter=51 channel=34
    26, 5, 52, 15, 10, 60, 9, 21, 25,
    -- layer=1 filter=51 channel=35
    0, 8, -4, 5, -8, 7, 5, 0, 4,
    -- layer=1 filter=51 channel=36
    24, 27, -1, 7, 27, 2, 4, 13, 12,
    -- layer=1 filter=51 channel=37
    -2, 6, -32, -19, -16, -23, 9, -37, -26,
    -- layer=1 filter=51 channel=38
    2, 2, 2, -16, -9, -10, 15, -11, -6,
    -- layer=1 filter=51 channel=39
    -17, 8, -12, 3, 7, -4, -18, -19, 3,
    -- layer=1 filter=51 channel=40
    17, -40, 10, -54, -43, -10, -17, -23, 26,
    -- layer=1 filter=51 channel=41
    -8, 17, -13, -32, 20, 20, 3, 35, 23,
    -- layer=1 filter=51 channel=42
    15, 11, 32, 29, -9, 25, 22, 31, 51,
    -- layer=1 filter=51 channel=43
    -34, -3, -45, -14, -6, -47, 25, -25, -21,
    -- layer=1 filter=51 channel=44
    8, 65, 30, 7, 55, 54, -16, 59, 38,
    -- layer=1 filter=51 channel=45
    -23, 2, -6, -16, 23, 13, -11, -3, 26,
    -- layer=1 filter=51 channel=46
    7, -36, -13, -27, -54, 5, -13, -47, -32,
    -- layer=1 filter=51 channel=47
    19, 39, 8, 40, 12, 7, 24, 22, 18,
    -- layer=1 filter=51 channel=48
    -5, -36, -28, 0, -47, -41, 2, -20, -20,
    -- layer=1 filter=51 channel=49
    9, 15, 31, -11, -4, 23, 21, 23, 24,
    -- layer=1 filter=51 channel=50
    0, 15, 12, -1, -16, 15, -4, -8, 12,
    -- layer=1 filter=51 channel=51
    -10, -42, -17, -10, -27, -10, 6, 0, -27,
    -- layer=1 filter=51 channel=52
    -17, -3, -6, -11, 0, 1, 0, 7, -16,
    -- layer=1 filter=51 channel=53
    -4, -14, -8, -1, -12, -4, -21, -4, 13,
    -- layer=1 filter=51 channel=54
    -10, -18, -58, 24, -28, -37, 50, 25, -51,
    -- layer=1 filter=51 channel=55
    10, 24, 18, 3, 31, 13, 7, 13, 14,
    -- layer=1 filter=51 channel=56
    5, -11, 6, -10, -10, 5, -8, 0, -2,
    -- layer=1 filter=51 channel=57
    9, -9, -11, 12, 9, -22, 26, 29, -19,
    -- layer=1 filter=51 channel=58
    42, 10, 27, 73, -23, -35, 62, 18, 10,
    -- layer=1 filter=51 channel=59
    -2, 5, -15, 10, 8, -6, 1, 3, -14,
    -- layer=1 filter=51 channel=60
    0, -3, 0, 12, -13, -15, 8, -10, -8,
    -- layer=1 filter=51 channel=61
    -2, -2, -2, -6, 6, -7, -10, -4, -4,
    -- layer=1 filter=51 channel=62
    -28, -3, -31, -36, -3, -47, -5, -27, -6,
    -- layer=1 filter=51 channel=63
    17, 8, 3, 9, 6, 1, 9, 11, 7,
    -- layer=1 filter=51 channel=64
    -18, -18, -10, -13, -14, -22, 4, 0, -3,
    -- layer=1 filter=51 channel=65
    -23, -29, -30, 1, -34, -40, 18, 5, -28,
    -- layer=1 filter=51 channel=66
    12, 2, -5, 15, 7, -10, 9, 0, -2,
    -- layer=1 filter=51 channel=67
    13, 15, 7, 1, -11, 11, 58, 27, 6,
    -- layer=1 filter=51 channel=68
    22, 45, 28, 19, 61, 44, 0, 73, 49,
    -- layer=1 filter=51 channel=69
    -22, 20, 7, -37, 23, 26, -32, 0, 34,
    -- layer=1 filter=51 channel=70
    22, 50, 37, -4, 8, 36, -8, -13, 41,
    -- layer=1 filter=51 channel=71
    -30, -8, 5, -15, 7, 7, 20, -3, -3,
    -- layer=1 filter=51 channel=72
    14, -33, -18, -29, -53, -58, 9, -40, -11,
    -- layer=1 filter=51 channel=73
    -1, 9, 17, 0, 6, 15, 3, 20, 14,
    -- layer=1 filter=51 channel=74
    24, 28, 0, -28, -11, -21, -2, 31, -16,
    -- layer=1 filter=51 channel=75
    1, -43, 8, -9, -10, -27, -19, -13, 19,
    -- layer=1 filter=51 channel=76
    3, 14, -25, -28, -2, 4, -9, 32, -4,
    -- layer=1 filter=51 channel=77
    -6, -6, -16, 10, 0, -33, 24, 12, -14,
    -- layer=1 filter=51 channel=78
    0, -3, -11, 6, 4, -24, -5, 13, -11,
    -- layer=1 filter=51 channel=79
    -23, -10, -10, -18, -2, -17, -1, -14, 0,
    -- layer=1 filter=51 channel=80
    -14, -14, 0, -2, -15, -7, 15, 0, -22,
    -- layer=1 filter=51 channel=81
    -19, -7, -5, 18, 7, 2, 12, 2, 27,
    -- layer=1 filter=51 channel=82
    -29, -41, -25, -19, -45, -11, 1, -21, -5,
    -- layer=1 filter=51 channel=83
    6, -2, 7, 5, 34, 27, 2, -5, 32,
    -- layer=1 filter=51 channel=84
    -9, -8, -21, -55, -35, -14, -12, 23, -10,
    -- layer=1 filter=51 channel=85
    11, -20, 11, 42, -22, -39, 30, -18, 18,
    -- layer=1 filter=51 channel=86
    -6, 9, -10, 6, 8, -6, -10, -7, -21,
    -- layer=1 filter=51 channel=87
    35, 10, 19, -16, -29, -25, 35, 4, -14,
    -- layer=1 filter=51 channel=88
    6, -4, 17, 3, -2, 16, 30, 10, 14,
    -- layer=1 filter=51 channel=89
    -36, -15, -29, -5, -32, -12, -9, 11, -26,
    -- layer=1 filter=51 channel=90
    33, 49, 24, 20, 72, 44, -9, 55, 63,
    -- layer=1 filter=51 channel=91
    1, -28, -33, -7, -57, -46, 13, -30, -38,
    -- layer=1 filter=51 channel=92
    -5, 35, -17, -17, 30, 4, -30, 30, -9,
    -- layer=1 filter=51 channel=93
    -18, -25, -20, -1, -5, -22, 3, -2, -21,
    -- layer=1 filter=51 channel=94
    -11, -19, -26, -6, 3, -32, 9, 8, -31,
    -- layer=1 filter=51 channel=95
    6, -5, -35, -61, -55, -27, -42, 12, -35,
    -- layer=1 filter=51 channel=96
    -5, 3, 1, 10, 0, 15, -1, 8, 4,
    -- layer=1 filter=51 channel=97
    0, -2, -25, 5, 11, -19, -2, 6, -12,
    -- layer=1 filter=51 channel=98
    -51, -11, -50, 7, 22, -32, 9, 0, 16,
    -- layer=1 filter=51 channel=99
    5, 31, -22, 25, 92, -45, 39, 85, -45,
    -- layer=1 filter=51 channel=100
    5, 19, 8, -9, 0, 6, -17, 18, 0,
    -- layer=1 filter=51 channel=101
    -10, -25, -18, -31, -49, -23, -20, -3, -19,
    -- layer=1 filter=51 channel=102
    -1, -14, -19, -1, -16, -33, 13, -10, -34,
    -- layer=1 filter=51 channel=103
    25, 13, 7, 0, -1, -4, -1, 1, -10,
    -- layer=1 filter=51 channel=104
    3, 20, 20, 25, 13, -6, 4, 5, 22,
    -- layer=1 filter=51 channel=105
    7, -1, -37, 13, 9, -21, 10, 5, -13,
    -- layer=1 filter=51 channel=106
    -4, 8, 10, -17, -3, 25, -22, 24, 17,
    -- layer=1 filter=51 channel=107
    5, 8, -1, 7, -9, 7, 1, -4, 13,
    -- layer=1 filter=51 channel=108
    13, 72, 33, 10, 63, 73, -1, 71, 53,
    -- layer=1 filter=51 channel=109
    2, 0, 0, 1, 0, -1, -8, 6, 4,
    -- layer=1 filter=51 channel=110
    -12, -16, -15, 0, 4, -20, -4, 3, -19,
    -- layer=1 filter=51 channel=111
    47, -15, -17, -46, -39, -34, -17, -14, -12,
    -- layer=1 filter=51 channel=112
    -12, -20, -16, -4, -28, -30, -12, 19, -26,
    -- layer=1 filter=51 channel=113
    42, 10, 65, 25, -17, 34, 2, 23, 68,
    -- layer=1 filter=51 channel=114
    6, 51, 16, 3, 45, 30, 39, -3, 20,
    -- layer=1 filter=51 channel=115
    -4, -15, -36, 3, -5, -36, 13, -1, -27,
    -- layer=1 filter=51 channel=116
    -3, 8, -8, -4, 3, -3, 3, -2, -4,
    -- layer=1 filter=51 channel=117
    -18, -19, -23, -47, -5, -68, -15, -6, 7,
    -- layer=1 filter=51 channel=118
    6, 2, -15, -63, -47, -22, -5, -15, -21,
    -- layer=1 filter=51 channel=119
    8, 64, 32, -12, 71, 52, -13, 67, 63,
    -- layer=1 filter=51 channel=120
    -15, -60, -31, 5, -38, -41, 31, -1, -2,
    -- layer=1 filter=51 channel=121
    16, 23, 8, -7, -1, -7, 19, 4, 32,
    -- layer=1 filter=51 channel=122
    3, 6, 5, 9, 10, 5, 1, -10, 5,
    -- layer=1 filter=51 channel=123
    31, 8, 8, 15, 7, 15, 27, 4, 5,
    -- layer=1 filter=51 channel=124
    3, -8, -1, -1, -1, -6, 16, 3, -10,
    -- layer=1 filter=51 channel=125
    5, 37, 30, -23, 14, 58, 16, 6, 43,
    -- layer=1 filter=51 channel=126
    -63, -35, -50, -4, 16, -52, -35, -26, 30,
    -- layer=1 filter=51 channel=127
    5, -22, -31, -65, -59, -30, -27, -23, -35,
    -- layer=1 filter=52 channel=0
    0, 8, -11, 7, 2, -1, 0, 6, -2,
    -- layer=1 filter=52 channel=1
    -6, 1, 2, -8, 1, 1, -7, 1, 3,
    -- layer=1 filter=52 channel=2
    10, -4, -1, 9, -7, 1, 9, 8, -10,
    -- layer=1 filter=52 channel=3
    -1, 5, 1, 0, 3, 3, 2, -2, 10,
    -- layer=1 filter=52 channel=4
    -10, -6, 5, 5, -9, 8, 5, 0, 7,
    -- layer=1 filter=52 channel=5
    -8, -12, -9, 2, 2, 1, -1, -4, 10,
    -- layer=1 filter=52 channel=6
    1, 3, -1, -2, -5, 10, -8, 1, 0,
    -- layer=1 filter=52 channel=7
    1, -6, 0, 6, -4, 0, 7, 5, -9,
    -- layer=1 filter=52 channel=8
    0, 1, -8, 2, -10, -3, -7, -8, 0,
    -- layer=1 filter=52 channel=9
    -7, 7, 9, 0, 5, 10, -7, 5, 3,
    -- layer=1 filter=52 channel=10
    -2, -4, 2, -8, -4, 7, -5, 7, -1,
    -- layer=1 filter=52 channel=11
    2, -2, 0, 7, -9, 7, -4, 2, 6,
    -- layer=1 filter=52 channel=12
    -7, -7, 8, 2, -8, 10, 8, 4, 7,
    -- layer=1 filter=52 channel=13
    -3, 7, -10, -2, 6, 4, 1, -7, 2,
    -- layer=1 filter=52 channel=14
    1, 3, -6, 9, -8, -6, -6, 6, 0,
    -- layer=1 filter=52 channel=15
    -5, -10, -2, 1, -8, -9, -8, 1, -9,
    -- layer=1 filter=52 channel=16
    -4, 4, -4, -4, -9, 4, -4, 3, -7,
    -- layer=1 filter=52 channel=17
    5, -7, 4, 0, 8, 6, 7, -6, -5,
    -- layer=1 filter=52 channel=18
    0, -11, 0, 0, 5, 6, -8, 0, -5,
    -- layer=1 filter=52 channel=19
    8, 2, 2, -11, 7, -11, -12, -3, -12,
    -- layer=1 filter=52 channel=20
    -11, 0, 4, 1, 3, -3, 1, 5, -6,
    -- layer=1 filter=52 channel=21
    -12, 5, -10, -10, -10, -6, 0, -2, -12,
    -- layer=1 filter=52 channel=22
    7, -12, -3, 8, 0, -10, -10, -1, 4,
    -- layer=1 filter=52 channel=23
    0, -11, 0, -4, 3, -7, 2, 5, 2,
    -- layer=1 filter=52 channel=24
    -5, -12, -6, 0, 8, -1, 2, -7, -3,
    -- layer=1 filter=52 channel=25
    -8, 0, 8, -11, -3, 3, -9, 6, 2,
    -- layer=1 filter=52 channel=26
    -3, -7, -5, -5, 5, 3, -3, 3, 6,
    -- layer=1 filter=52 channel=27
    -6, -3, 4, -10, -6, -10, -5, 2, -13,
    -- layer=1 filter=52 channel=28
    -8, -4, -7, 4, 1, -6, 0, 7, -11,
    -- layer=1 filter=52 channel=29
    3, -3, 6, 1, -2, 9, -6, -1, 6,
    -- layer=1 filter=52 channel=30
    -5, 6, 4, 1, -9, 11, 4, 0, -3,
    -- layer=1 filter=52 channel=31
    -7, -9, 0, -6, -8, -1, -5, -4, 6,
    -- layer=1 filter=52 channel=32
    -9, -9, -2, -10, 5, -1, -5, -8, 8,
    -- layer=1 filter=52 channel=33
    7, 6, 5, 1, -5, -8, -5, -2, -9,
    -- layer=1 filter=52 channel=34
    -1, 7, 1, -8, -2, -6, -12, 8, 7,
    -- layer=1 filter=52 channel=35
    -5, 7, 2, 1, 0, -8, 1, -8, 4,
    -- layer=1 filter=52 channel=36
    4, 1, 8, -3, -2, 6, -6, -11, 3,
    -- layer=1 filter=52 channel=37
    -14, 1, 1, 2, -5, -7, 10, 0, 1,
    -- layer=1 filter=52 channel=38
    -6, -7, -4, 2, -9, 6, -12, 3, 6,
    -- layer=1 filter=52 channel=39
    2, 7, 7, 4, 4, -9, 5, 1, -7,
    -- layer=1 filter=52 channel=40
    -6, 0, 9, -1, -10, 3, -8, 1, -4,
    -- layer=1 filter=52 channel=41
    -2, -8, 0, -5, 5, -3, 4, 1, -10,
    -- layer=1 filter=52 channel=42
    0, 0, 0, -5, -2, 3, -9, -6, -4,
    -- layer=1 filter=52 channel=43
    4, -2, -11, -12, 8, 3, -5, -12, -6,
    -- layer=1 filter=52 channel=44
    -6, -10, 7, 7, 7, 4, 6, 0, -6,
    -- layer=1 filter=52 channel=45
    2, 0, 1, 1, 4, -5, -12, 7, -4,
    -- layer=1 filter=52 channel=46
    -7, -7, -6, 0, -1, 10, -8, 0, 7,
    -- layer=1 filter=52 channel=47
    -10, -8, 8, -2, -6, -7, -8, -4, 9,
    -- layer=1 filter=52 channel=48
    0, 1, -8, 7, -12, -4, 4, 5, -3,
    -- layer=1 filter=52 channel=49
    5, -3, -8, -3, 8, -9, -3, -5, -5,
    -- layer=1 filter=52 channel=50
    -9, -7, -1, -1, -5, -5, -12, 1, -2,
    -- layer=1 filter=52 channel=51
    -7, 0, 6, 3, -6, 1, -4, 7, -11,
    -- layer=1 filter=52 channel=52
    -2, 1, 0, 8, -5, 0, -2, 3, -1,
    -- layer=1 filter=52 channel=53
    1, -9, -5, 0, -3, -2, -6, -5, 1,
    -- layer=1 filter=52 channel=54
    5, 1, 4, 0, -10, -1, 2, -1, 2,
    -- layer=1 filter=52 channel=55
    -4, -5, 0, 4, -7, 6, 0, -5, 3,
    -- layer=1 filter=52 channel=56
    -6, 2, -5, -11, 0, -2, -4, 0, -7,
    -- layer=1 filter=52 channel=57
    -7, -7, -6, -1, 0, 1, -3, -4, -1,
    -- layer=1 filter=52 channel=58
    7, 9, -6, -8, -10, 0, 6, -2, 8,
    -- layer=1 filter=52 channel=59
    4, -11, 2, 7, -6, -6, 5, -5, -11,
    -- layer=1 filter=52 channel=60
    10, 0, 2, -2, -1, 3, 8, 1, -2,
    -- layer=1 filter=52 channel=61
    9, 0, 2, 6, 1, -3, -8, -9, 7,
    -- layer=1 filter=52 channel=62
    6, -2, 1, 5, -12, 8, -3, 0, 0,
    -- layer=1 filter=52 channel=63
    0, 6, 7, -3, -1, 0, 1, -1, 2,
    -- layer=1 filter=52 channel=64
    -4, -12, 0, -10, 1, -2, 3, 5, -11,
    -- layer=1 filter=52 channel=65
    -12, -12, 2, -7, 1, 2, -2, -10, 1,
    -- layer=1 filter=52 channel=66
    -8, 0, -8, 2, 4, 0, -7, 3, 5,
    -- layer=1 filter=52 channel=67
    7, -7, 6, 1, 0, 1, 0, 7, 1,
    -- layer=1 filter=52 channel=68
    -11, -6, 5, 7, -2, -10, -1, 4, -6,
    -- layer=1 filter=52 channel=69
    -6, -4, 3, -12, 5, 1, -8, 1, -5,
    -- layer=1 filter=52 channel=70
    0, 7, -2, -10, -3, 7, -2, -6, -4,
    -- layer=1 filter=52 channel=71
    -7, -12, 6, -2, -1, -11, 2, 5, -8,
    -- layer=1 filter=52 channel=72
    8, -10, 0, 3, -11, -2, 2, -1, -6,
    -- layer=1 filter=52 channel=73
    5, 0, -1, -7, 3, 6, -12, 5, 4,
    -- layer=1 filter=52 channel=74
    4, 2, -5, 2, -2, 2, -12, 7, -10,
    -- layer=1 filter=52 channel=75
    5, 5, -5, -2, -3, 0, 10, -8, 6,
    -- layer=1 filter=52 channel=76
    0, -11, -9, -5, -2, 2, -3, -6, -3,
    -- layer=1 filter=52 channel=77
    4, 2, 1, -7, 0, -9, 3, -5, -6,
    -- layer=1 filter=52 channel=78
    -10, 0, -3, -5, 8, 7, -9, 6, -6,
    -- layer=1 filter=52 channel=79
    -11, 4, -7, -1, 4, -4, -7, -2, -3,
    -- layer=1 filter=52 channel=80
    -2, 10, 0, 8, 3, 7, -3, 1, 7,
    -- layer=1 filter=52 channel=81
    -2, 3, 8, 6, -9, -7, 7, 4, 6,
    -- layer=1 filter=52 channel=82
    10, 0, -2, 3, -8, -4, -12, -5, -6,
    -- layer=1 filter=52 channel=83
    -3, -12, -11, 1, 0, -11, 3, 2, -8,
    -- layer=1 filter=52 channel=84
    6, 1, -10, -12, -7, -5, -5, -8, 0,
    -- layer=1 filter=52 channel=85
    -5, -9, -6, 7, 7, -6, -5, 5, 2,
    -- layer=1 filter=52 channel=86
    -5, -6, -6, -6, 2, 4, -10, -11, 0,
    -- layer=1 filter=52 channel=87
    -10, -4, -6, 5, -5, 5, 0, -12, -9,
    -- layer=1 filter=52 channel=88
    0, -7, -9, 3, 1, 1, -7, 4, 8,
    -- layer=1 filter=52 channel=89
    5, 2, 4, 0, -10, -7, 4, -5, 2,
    -- layer=1 filter=52 channel=90
    -8, 2, 7, 1, 2, -12, 5, -4, 4,
    -- layer=1 filter=52 channel=91
    8, 3, -6, 0, -4, -8, 0, 7, 5,
    -- layer=1 filter=52 channel=92
    5, -2, -6, -7, -8, -5, -11, -3, -9,
    -- layer=1 filter=52 channel=93
    -3, -3, 0, -8, 4, 6, 6, -2, 6,
    -- layer=1 filter=52 channel=94
    6, 0, 4, -4, -10, -9, 0, 3, -7,
    -- layer=1 filter=52 channel=95
    7, -7, 3, 6, -1, -2, -5, -6, -4,
    -- layer=1 filter=52 channel=96
    -6, -8, -4, -8, -2, -11, -8, -11, 8,
    -- layer=1 filter=52 channel=97
    -2, 2, -1, 8, -10, -10, 0, 4, -9,
    -- layer=1 filter=52 channel=98
    -6, 4, 1, 3, 8, -7, 7, -2, 7,
    -- layer=1 filter=52 channel=99
    -11, 5, -11, 8, -4, -5, -8, -2, 4,
    -- layer=1 filter=52 channel=100
    2, -9, -2, -11, -7, -2, -3, 4, -10,
    -- layer=1 filter=52 channel=101
    1, 7, -6, -7, -5, -5, 0, -8, -12,
    -- layer=1 filter=52 channel=102
    7, -3, 3, 0, -5, -11, -12, 1, 5,
    -- layer=1 filter=52 channel=103
    -1, -7, 4, 2, 5, 5, 7, -11, -10,
    -- layer=1 filter=52 channel=104
    -3, -7, 6, -6, -7, -3, -1, -6, -11,
    -- layer=1 filter=52 channel=105
    -11, -10, -6, -7, 0, -10, 6, 0, -3,
    -- layer=1 filter=52 channel=106
    2, 0, -9, 1, -2, 0, 0, -9, -11,
    -- layer=1 filter=52 channel=107
    6, -1, 2, 8, 5, -1, 2, -3, -9,
    -- layer=1 filter=52 channel=108
    2, -1, 0, 1, -7, 3, -11, -8, 4,
    -- layer=1 filter=52 channel=109
    1, 8, -4, 2, 2, -6, -10, -11, 8,
    -- layer=1 filter=52 channel=110
    2, -10, -5, 2, 0, 0, 7, 0, -9,
    -- layer=1 filter=52 channel=111
    6, 0, 8, -2, -7, 6, 0, -9, 4,
    -- layer=1 filter=52 channel=112
    -1, 4, -5, 4, 5, 4, 2, -7, 5,
    -- layer=1 filter=52 channel=113
    -6, 4, -4, -3, 5, -12, 6, -10, -10,
    -- layer=1 filter=52 channel=114
    1, -3, -10, -12, -2, 1, 4, 0, 8,
    -- layer=1 filter=52 channel=115
    6, -3, -6, -9, 0, 1, 7, -7, 0,
    -- layer=1 filter=52 channel=116
    -3, 2, 6, -9, 4, -8, 0, 0, -5,
    -- layer=1 filter=52 channel=117
    -2, -6, 0, 1, 0, 6, 1, 3, -9,
    -- layer=1 filter=52 channel=118
    3, 8, 0, -9, 2, 6, -4, 2, -10,
    -- layer=1 filter=52 channel=119
    8, -8, -1, -9, -2, 5, 3, 6, 7,
    -- layer=1 filter=52 channel=120
    0, 0, 9, -7, -11, 3, 1, -4, 3,
    -- layer=1 filter=52 channel=121
    -7, 0, -8, -7, 9, -9, -8, 1, -11,
    -- layer=1 filter=52 channel=122
    9, 0, 0, -9, 4, 3, 1, 6, 8,
    -- layer=1 filter=52 channel=123
    -9, -12, 4, 5, 7, 0, -10, -10, -1,
    -- layer=1 filter=52 channel=124
    11, 0, 6, -9, 7, 1, 1, 0, -6,
    -- layer=1 filter=52 channel=125
    -2, 3, 8, -9, -1, -9, -8, 8, 9,
    -- layer=1 filter=52 channel=126
    -9, 3, 10, -10, 4, 7, 5, 1, -5,
    -- layer=1 filter=52 channel=127
    8, 0, -11, -8, -9, -9, 8, 3, 1,
    -- layer=1 filter=53 channel=0
    -38, -1, 24, -43, 3, 14, 4, 22, 24,
    -- layer=1 filter=53 channel=1
    -33, -16, 33, 20, 45, 31, 33, 14, -25,
    -- layer=1 filter=53 channel=2
    5, 47, 16, 16, -8, -36, 26, -5, -37,
    -- layer=1 filter=53 channel=3
    3, -2, 3, 1, 4, -1, 5, 0, 1,
    -- layer=1 filter=53 channel=4
    -19, -13, -18, -4, -5, 12, -14, -19, -4,
    -- layer=1 filter=53 channel=5
    -56, 3, 28, 21, 65, 42, 43, 24, -5,
    -- layer=1 filter=53 channel=6
    57, -5, -22, 78, -17, -27, -1, -67, -41,
    -- layer=1 filter=53 channel=7
    -43, 44, 56, 45, 61, 28, 54, 54, -18,
    -- layer=1 filter=53 channel=8
    -54, -15, 48, 17, 52, 27, 25, 10, -14,
    -- layer=1 filter=53 channel=9
    36, 28, 5, -2, -76, -75, -52, -26, -58,
    -- layer=1 filter=53 channel=10
    -33, 51, 45, 43, 64, 0, 59, 32, -35,
    -- layer=1 filter=53 channel=11
    -38, -68, 9, -97, -37, 40, -44, 6, 54,
    -- layer=1 filter=53 channel=12
    -42, 34, -49, -15, 16, 1, 23, 1, 23,
    -- layer=1 filter=53 channel=13
    44, -7, -29, 20, -38, -27, -11, -47, -25,
    -- layer=1 filter=53 channel=14
    -115, -5, 14, -52, 1, -16, -10, -8, -31,
    -- layer=1 filter=53 channel=15
    13, 1, -31, 1, -73, 16, -55, -6, -26,
    -- layer=1 filter=53 channel=16
    -47, 33, 53, 35, 62, 22, 36, 2, -13,
    -- layer=1 filter=53 channel=17
    -26, -22, 33, -40, -1, 18, -6, 0, 15,
    -- layer=1 filter=53 channel=18
    13, -11, -46, -25, -2, 20, -50, 1, 5,
    -- layer=1 filter=53 channel=19
    42, 36, 34, 58, 6, -20, -6, -40, -82,
    -- layer=1 filter=53 channel=20
    26, 8, 1, 20, -1, -8, 4, -32, -30,
    -- layer=1 filter=53 channel=21
    16, 3, -10, 17, 15, -8, -5, 4, -46,
    -- layer=1 filter=53 channel=22
    26, -11, 4, 15, -4, -15, -1, -2, -23,
    -- layer=1 filter=53 channel=23
    -64, -74, -41, -43, -73, -70, -18, -33, -28,
    -- layer=1 filter=53 channel=24
    4, -5, -28, -4, -9, -56, -2, -50, -21,
    -- layer=1 filter=53 channel=25
    -21, 63, 62, 56, 82, 19, 77, 49, -32,
    -- layer=1 filter=53 channel=26
    15, -48, -40, -54, -116, -32, -58, -63, 0,
    -- layer=1 filter=53 channel=27
    -65, 6, 27, -31, 20, 13, 25, 33, 42,
    -- layer=1 filter=53 channel=28
    -57, 44, 47, 18, 74, 22, 42, 41, -23,
    -- layer=1 filter=53 channel=29
    -13, 10, 7, 20, -6, 6, 43, 44, 20,
    -- layer=1 filter=53 channel=30
    48, -44, -62, -17, -50, -16, -85, -29, -8,
    -- layer=1 filter=53 channel=31
    12, -9, -26, 16, -26, -20, -5, -40, -36,
    -- layer=1 filter=53 channel=32
    3, -57, -52, -9, -150, -26, -44, -55, 6,
    -- layer=1 filter=53 channel=33
    11, 8, 28, 11, 7, 17, -1, -7, 11,
    -- layer=1 filter=53 channel=34
    20, 14, -2, -18, -34, -22, -19, -56, -66,
    -- layer=1 filter=53 channel=35
    -18, -28, -36, -23, -19, 9, -20, -25, -18,
    -- layer=1 filter=53 channel=36
    -59, -33, 17, -105, -16, 44, -40, 29, 64,
    -- layer=1 filter=53 channel=37
    -23, 43, 47, 48, 64, 32, 42, 28, -23,
    -- layer=1 filter=53 channel=38
    48, 16, -3, 26, 1, -22, -17, -41, -33,
    -- layer=1 filter=53 channel=39
    -63, -1, 1, -38, -8, 17, -13, 19, 6,
    -- layer=1 filter=53 channel=40
    37, 0, -18, 41, 0, -20, -23, -23, -56,
    -- layer=1 filter=53 channel=41
    43, -8, -25, 23, -36, -16, 13, -32, -13,
    -- layer=1 filter=53 channel=42
    14, 41, 37, 7, 10, -10, 21, -11, -19,
    -- layer=1 filter=53 channel=43
    -36, 9, 29, 13, 61, 16, 53, 13, -27,
    -- layer=1 filter=53 channel=44
    -9, -86, -55, -42, -105, -12, -64, -34, 6,
    -- layer=1 filter=53 channel=45
    5, -26, -5, 12, -24, 1, -11, -22, -25,
    -- layer=1 filter=53 channel=46
    27, 19, 58, 46, 37, 14, 18, -29, -15,
    -- layer=1 filter=53 channel=47
    39, -6, -31, 37, -12, -47, 44, -33, -98,
    -- layer=1 filter=53 channel=48
    38, 8, -28, 30, 0, -31, 23, -15, -20,
    -- layer=1 filter=53 channel=49
    62, 44, -10, 63, 3, -44, 26, -27, -65,
    -- layer=1 filter=53 channel=50
    4, 2, 15, 0, 6, 6, 6, 5, -4,
    -- layer=1 filter=53 channel=51
    8, 22, 11, 24, 29, -21, 9, 0, -28,
    -- layer=1 filter=53 channel=52
    2, -23, 0, 7, -2, -17, 30, 21, 10,
    -- layer=1 filter=53 channel=53
    24, 12, 21, 3, 7, 10, 9, 4, 15,
    -- layer=1 filter=53 channel=54
    -30, 39, 54, 56, 91, 4, 50, 20, -42,
    -- layer=1 filter=53 channel=55
    -62, -36, -11, -37, -2, 25, -11, 29, 73,
    -- layer=1 filter=53 channel=56
    7, -10, 3, -5, -3, -5, 3, 9, 6,
    -- layer=1 filter=53 channel=57
    -20, 42, 32, 42, 50, -4, 34, 36, -39,
    -- layer=1 filter=53 channel=58
    -1, 25, 16, 52, 13, -37, 36, 6, -45,
    -- layer=1 filter=53 channel=59
    -4, -1, 14, 13, 1, 23, 1, 12, -7,
    -- layer=1 filter=53 channel=60
    -17, -31, 27, 13, 11, 27, 3, 43, 7,
    -- layer=1 filter=53 channel=61
    -8, -8, 6, -6, 4, 7, -9, 3, -7,
    -- layer=1 filter=53 channel=62
    -38, 26, 43, 32, 67, 20, 39, 15, -11,
    -- layer=1 filter=53 channel=63
    -46, -42, 1, -91, -21, 48, -34, 29, 49,
    -- layer=1 filter=53 channel=64
    5, -3, -11, 2, 12, -14, -3, 13, -19,
    -- layer=1 filter=53 channel=65
    29, 9, -5, 17, -7, -22, -14, -14, -19,
    -- layer=1 filter=53 channel=66
    -79, -16, 23, -57, 6, 39, 3, 38, 37,
    -- layer=1 filter=53 channel=67
    38, 9, -4, 22, 3, -25, 22, -2, -10,
    -- layer=1 filter=53 channel=68
    -29, -101, -32, -62, -112, 24, -87, -2, 36,
    -- layer=1 filter=53 channel=69
    -54, -14, -18, -6, -18, -7, -6, -19, -19,
    -- layer=1 filter=53 channel=70
    -10, -9, -15, 52, 19, 0, 26, -3, -11,
    -- layer=1 filter=53 channel=71
    -29, -3, -6, -1, 20, -6, -1, 3, -18,
    -- layer=1 filter=53 channel=72
    45, -18, -22, -10, -56, 32, -56, -42, -48,
    -- layer=1 filter=53 channel=73
    -2, -2, 11, 0, -18, 2, 5, -4, -3,
    -- layer=1 filter=53 channel=74
    -30, -50, -20, -7, -24, 32, -62, 36, 37,
    -- layer=1 filter=53 channel=75
    -28, -43, -23, -79, -41, -23, -34, -68, -22,
    -- layer=1 filter=53 channel=76
    -19, -67, -28, -69, -15, 7, -59, -2, 39,
    -- layer=1 filter=53 channel=77
    11, 21, -17, 8, 37, -27, 17, 0, -34,
    -- layer=1 filter=53 channel=78
    -43, 12, 15, 0, 35, 9, 14, 10, -4,
    -- layer=1 filter=53 channel=79
    -20, 10, 36, 35, 46, 8, 29, -5, -23,
    -- layer=1 filter=53 channel=80
    -37, 0, 33, -4, -21, 26, 39, 22, -1,
    -- layer=1 filter=53 channel=81
    -10, 13, 0, 0, 13, -22, 23, 8, -11,
    -- layer=1 filter=53 channel=82
    39, 19, -24, 36, 13, -44, 15, -27, -52,
    -- layer=1 filter=53 channel=83
    0, -58, -12, 6, -8, 35, -8, 5, 6,
    -- layer=1 filter=53 channel=84
    45, -42, -61, -39, -1, 0, -71, -19, 39,
    -- layer=1 filter=53 channel=85
    15, -8, 6, 45, -22, -34, 33, -13, -35,
    -- layer=1 filter=53 channel=86
    -79, -20, 39, -41, 11, 30, 9, 39, 35,
    -- layer=1 filter=53 channel=87
    45, 44, 55, 41, -26, -14, -3, -5, -55,
    -- layer=1 filter=53 channel=88
    28, 12, 2, 22, 2, -24, -9, -15, -15,
    -- layer=1 filter=53 channel=89
    36, 2, -43, 30, -19, -31, -17, -37, -24,
    -- layer=1 filter=53 channel=90
    -29, -83, -64, -50, -93, -24, -51, -42, 3,
    -- layer=1 filter=53 channel=91
    51, 22, -5, 32, 24, -15, 18, -7, -27,
    -- layer=1 filter=53 channel=92
    26, 45, -41, 42, -28, 13, -20, -1, -4,
    -- layer=1 filter=53 channel=93
    4, -4, 10, 7, 1, -1, 6, 10, 0,
    -- layer=1 filter=53 channel=94
    -47, 14, 34, -30, 16, 22, -8, 37, 13,
    -- layer=1 filter=53 channel=95
    21, -48, -73, -79, -22, -2, -80, -23, 24,
    -- layer=1 filter=53 channel=96
    -2, -15, -5, -19, -1, 8, -9, 5, 11,
    -- layer=1 filter=53 channel=97
    -28, -3, 13, -29, 16, 14, 0, 24, 25,
    -- layer=1 filter=53 channel=98
    -32, -6, 28, 3, 67, 2, 33, 11, -27,
    -- layer=1 filter=53 channel=99
    -121, -11, 7, -78, -5, -18, -16, 34, -39,
    -- layer=1 filter=53 channel=100
    -49, -60, 0, -60, -18, 70, -42, 3, 49,
    -- layer=1 filter=53 channel=101
    41, -10, -13, 23, -12, -10, 7, -18, -26,
    -- layer=1 filter=53 channel=102
    -21, -6, 14, 2, 10, 13, -8, 13, 6,
    -- layer=1 filter=53 channel=103
    -41, -41, -1, -50, -47, 34, -20, 19, 58,
    -- layer=1 filter=53 channel=104
    7, -34, -45, -13, -44, -28, -21, 5, 11,
    -- layer=1 filter=53 channel=105
    -40, -9, 15, -42, 9, 32, 6, 37, 12,
    -- layer=1 filter=53 channel=106
    33, -36, -44, 30, -71, -29, -36, -61, -6,
    -- layer=1 filter=53 channel=107
    26, 13, 16, 23, 5, 18, 13, 17, 1,
    -- layer=1 filter=53 channel=108
    -19, -55, -53, -43, -108, -13, -50, -48, -7,
    -- layer=1 filter=53 channel=109
    0, 1, 4, -3, 0, 1, 2, -4, -10,
    -- layer=1 filter=53 channel=110
    -12, 0, 2, 2, 17, 2, 0, -1, 17,
    -- layer=1 filter=53 channel=111
    12, -36, -67, -25, -43, 0, -77, -3, 8,
    -- layer=1 filter=53 channel=112
    22, -27, -37, -12, -7, -26, -42, -13, 43,
    -- layer=1 filter=53 channel=113
    59, 53, 34, 31, 6, -15, 9, -7, -41,
    -- layer=1 filter=53 channel=114
    -46, -21, 8, -2, 1, 20, 0, 16, 1,
    -- layer=1 filter=53 channel=115
    -51, 11, 32, -20, 22, 11, 24, 30, -15,
    -- layer=1 filter=53 channel=116
    -4, -2, 5, 10, -8, 0, -1, -9, -9,
    -- layer=1 filter=53 channel=117
    -7, -58, -61, -36, -70, -29, -23, -14, -12,
    -- layer=1 filter=53 channel=118
    21, -49, -47, -30, -45, 23, -75, 6, 35,
    -- layer=1 filter=53 channel=119
    0, -74, -47, -50, -86, -18, -34, -22, 23,
    -- layer=1 filter=53 channel=120
    13, 38, 8, 34, 46, -16, 22, 2, -62,
    -- layer=1 filter=53 channel=121
    -32, -57, -28, -53, -50, -32, -57, -43, -33,
    -- layer=1 filter=53 channel=122
    8, 0, -3, 9, 8, -2, 8, 1, 10,
    -- layer=1 filter=53 channel=123
    -36, -58, -17, -58, -48, -14, -36, -10, 0,
    -- layer=1 filter=53 channel=124
    -14, 3, 3, -3, 17, 3, -1, -14, 0,
    -- layer=1 filter=53 channel=125
    2, 37, -23, 64, 13, -3, 26, 22, -38,
    -- layer=1 filter=53 channel=126
    -64, -22, 14, 10, 61, 14, 55, 19, -4,
    -- layer=1 filter=53 channel=127
    8, -48, -66, -67, -1, 26, -51, -15, 19,
    -- layer=1 filter=54 channel=0
    -10, -16, 13, -23, -10, 12, -15, 1, 14,
    -- layer=1 filter=54 channel=1
    -15, -29, 14, -34, 8, -10, -7, 8, -28,
    -- layer=1 filter=54 channel=2
    13, 16, -6, 37, 7, -13, 13, 11, -13,
    -- layer=1 filter=54 channel=3
    1, 2, 5, -3, 4, -9, 1, 10, -2,
    -- layer=1 filter=54 channel=4
    -9, -10, -3, -14, -4, -14, 1, -13, -17,
    -- layer=1 filter=54 channel=5
    -14, -17, 32, -7, 9, -6, -7, -11, -33,
    -- layer=1 filter=54 channel=6
    16, 16, -8, 12, 10, -15, 14, 0, -1,
    -- layer=1 filter=54 channel=7
    -35, 51, 55, 12, 74, 44, 68, 64, 36,
    -- layer=1 filter=54 channel=8
    -23, -41, 17, -40, -15, -17, -2, -17, -46,
    -- layer=1 filter=54 channel=9
    -23, -20, -35, 0, -32, -15, 0, 5, -62,
    -- layer=1 filter=54 channel=10
    -27, 51, 33, 13, 62, 38, 46, 60, 27,
    -- layer=1 filter=54 channel=11
    -8, -31, -3, -12, -18, 11, 2, 0, 21,
    -- layer=1 filter=54 channel=12
    -15, -15, -29, -49, -42, -46, -46, -76, -49,
    -- layer=1 filter=54 channel=13
    17, -13, -18, 14, -32, -39, 0, -8, -20,
    -- layer=1 filter=54 channel=14
    -55, 6, 25, -33, 16, -19, 7, 7, 11,
    -- layer=1 filter=54 channel=15
    0, -3, -13, 30, 2, -36, -13, 12, -5,
    -- layer=1 filter=54 channel=16
    -61, -14, 34, -6, -4, -13, 0, -27, -20,
    -- layer=1 filter=54 channel=17
    -8, -29, -2, -23, -13, 7, -16, -6, -10,
    -- layer=1 filter=54 channel=18
    4, 2, -9, -3, -41, -29, -21, -22, -6,
    -- layer=1 filter=54 channel=19
    -43, 46, 25, 46, 12, -41, 24, -16, -41,
    -- layer=1 filter=54 channel=20
    0, -5, -5, -1, -2, -8, -14, -10, -10,
    -- layer=1 filter=54 channel=21
    -14, -5, -12, -15, 10, 12, -11, 1, 9,
    -- layer=1 filter=54 channel=22
    15, -19, -1, -20, -6, 3, 8, 14, -5,
    -- layer=1 filter=54 channel=23
    -59, 17, -14, -13, 21, -18, 38, 23, 12,
    -- layer=1 filter=54 channel=24
    6, 0, -4, 9, -21, -40, 8, -21, -30,
    -- layer=1 filter=54 channel=25
    -49, 40, 37, 6, 55, 36, 55, 25, 18,
    -- layer=1 filter=54 channel=26
    21, 5, -37, 26, -27, -60, 26, -21, -44,
    -- layer=1 filter=54 channel=27
    -65, -55, 0, -69, -30, 0, -28, -29, 27,
    -- layer=1 filter=54 channel=28
    -71, 9, 32, -28, 54, 35, 22, 37, 20,
    -- layer=1 filter=54 channel=29
    -12, 2, 36, -3, 14, 33, 2, 5, 8,
    -- layer=1 filter=54 channel=30
    -17, -8, -10, 14, -40, -48, -35, -53, -44,
    -- layer=1 filter=54 channel=31
    19, 24, -12, 0, -5, -28, 3, -24, -16,
    -- layer=1 filter=54 channel=32
    -4, 37, -47, 24, 1, -39, 16, 13, -34,
    -- layer=1 filter=54 channel=33
    -14, -31, -24, -16, -18, 0, 14, 0, -7,
    -- layer=1 filter=54 channel=34
    10, -39, -47, -28, -22, -43, 11, -17, -6,
    -- layer=1 filter=54 channel=35
    -9, -11, 25, -1, 4, 2, -14, -9, 10,
    -- layer=1 filter=54 channel=36
    -14, -19, -10, -1, -8, 29, 10, 5, 27,
    -- layer=1 filter=54 channel=37
    -55, 40, 32, 18, 30, -3, 1, 0, -23,
    -- layer=1 filter=54 channel=38
    0, -7, 4, 13, -13, -6, -9, 1, 4,
    -- layer=1 filter=54 channel=39
    -11, -6, 15, -41, -31, 7, -2, 2, 0,
    -- layer=1 filter=54 channel=40
    34, 21, 22, 2, -5, -2, 6, 10, 16,
    -- layer=1 filter=54 channel=41
    -24, 56, -2, 18, 14, -14, 20, 22, -25,
    -- layer=1 filter=54 channel=42
    18, 33, 20, 31, 44, 11, 43, 22, -3,
    -- layer=1 filter=54 channel=43
    -41, -7, 33, -9, 25, 2, 12, 13, -13,
    -- layer=1 filter=54 channel=44
    17, -10, -50, 21, -28, -69, 21, -25, -40,
    -- layer=1 filter=54 channel=45
    0, -33, -12, -1, -33, -30, -12, -25, -26,
    -- layer=1 filter=54 channel=46
    -22, -5, 0, 47, 8, -14, 9, -17, -6,
    -- layer=1 filter=54 channel=47
    11, 70, -52, 44, 47, -58, 42, 27, -37,
    -- layer=1 filter=54 channel=48
    -13, -12, -18, -2, 6, 14, -20, 0, 17,
    -- layer=1 filter=54 channel=49
    20, 0, -19, 20, 2, -5, 15, 4, -10,
    -- layer=1 filter=54 channel=50
    -29, -14, -34, -8, -26, -42, -18, -15, -14,
    -- layer=1 filter=54 channel=51
    -11, 4, 3, -13, 15, 8, 9, 13, 3,
    -- layer=1 filter=54 channel=52
    11, 17, 11, -5, 0, -11, 4, 7, 1,
    -- layer=1 filter=54 channel=53
    4, 14, 7, -3, 5, 6, 9, 21, 21,
    -- layer=1 filter=54 channel=54
    -47, 53, 39, 44, 61, 22, 55, 34, 10,
    -- layer=1 filter=54 channel=55
    -3, 3, 16, 5, 0, 30, 10, 23, 12,
    -- layer=1 filter=54 channel=56
    -5, 11, 4, -8, -1, 5, 10, 1, 2,
    -- layer=1 filter=54 channel=57
    -14, 45, 28, 18, 60, 36, 23, 36, 40,
    -- layer=1 filter=54 channel=58
    -25, 68, 21, 56, 64, 21, 64, 46, 16,
    -- layer=1 filter=54 channel=59
    -18, -32, 7, -4, -1, -11, -15, -18, 0,
    -- layer=1 filter=54 channel=60
    -14, 25, 7, -1, 16, 14, -1, 20, -2,
    -- layer=1 filter=54 channel=61
    -2, -11, -12, -10, -17, -3, -8, -9, -8,
    -- layer=1 filter=54 channel=62
    -48, 7, 43, -17, 4, -7, 15, -8, -35,
    -- layer=1 filter=54 channel=63
    -18, -36, -22, -3, -19, 22, -9, 4, 23,
    -- layer=1 filter=54 channel=64
    -2, -8, 4, -15, -15, -4, -6, -1, 5,
    -- layer=1 filter=54 channel=65
    -12, -24, -13, -31, -16, 11, -22, -8, 8,
    -- layer=1 filter=54 channel=66
    -19, -24, 5, -21, -1, 33, 1, 9, 22,
    -- layer=1 filter=54 channel=67
    15, -29, -9, -10, 9, 4, 2, 8, 15,
    -- layer=1 filter=54 channel=68
    32, -4, 3, 36, -36, -32, 12, -19, -21,
    -- layer=1 filter=54 channel=69
    -14, -12, -5, 2, -13, -56, -4, -29, -53,
    -- layer=1 filter=54 channel=70
    -5, -19, -15, 2, -5, -5, -22, -11, 0,
    -- layer=1 filter=54 channel=71
    -42, -11, 12, 0, 23, 24, 6, 9, 16,
    -- layer=1 filter=54 channel=72
    0, 10, -14, 38, -14, -18, -5, -18, -23,
    -- layer=1 filter=54 channel=73
    5, -15, 0, 4, 6, 4, 12, -7, -10,
    -- layer=1 filter=54 channel=74
    16, -27, 10, 24, -43, -45, 13, -1, -10,
    -- layer=1 filter=54 channel=75
    -41, -22, -27, -47, -59, -70, -51, -93, -62,
    -- layer=1 filter=54 channel=76
    -3, -35, -24, 18, -70, 2, -6, -15, -4,
    -- layer=1 filter=54 channel=77
    -20, -18, 1, -9, -2, 18, -20, 5, 5,
    -- layer=1 filter=54 channel=78
    -65, -15, -6, -20, 3, 2, 0, 0, 9,
    -- layer=1 filter=54 channel=79
    -39, 5, 18, -6, 2, -24, 6, 0, -31,
    -- layer=1 filter=54 channel=80
    -4, -15, 21, -1, -2, 17, 23, 5, 18,
    -- layer=1 filter=54 channel=81
    -33, -5, -2, -25, -8, 17, 9, 4, 13,
    -- layer=1 filter=54 channel=82
    -6, 2, -9, -1, -9, -5, -11, -4, -2,
    -- layer=1 filter=54 channel=83
    -8, -33, -23, -14, -42, -28, -12, -6, -22,
    -- layer=1 filter=54 channel=84
    13, -4, -24, 27, -77, -55, 14, -47, -30,
    -- layer=1 filter=54 channel=85
    -3, 59, -14, 1, 29, -28, 43, 14, -9,
    -- layer=1 filter=54 channel=86
    -14, -21, 18, -9, 10, 28, 3, 2, 17,
    -- layer=1 filter=54 channel=87
    -12, 34, 5, 50, -15, -7, 23, -2, -24,
    -- layer=1 filter=54 channel=88
    0, -8, -17, -4, -8, -6, -6, -10, 0,
    -- layer=1 filter=54 channel=89
    -3, -25, -31, 0, -34, -7, -17, -10, 8,
    -- layer=1 filter=54 channel=90
    1, -28, -22, 7, -38, -62, 6, -36, -53,
    -- layer=1 filter=54 channel=91
    12, 11, 6, 4, -4, 11, -15, 3, 9,
    -- layer=1 filter=54 channel=92
    18, -7, -36, 22, 1, -24, 15, -3, -4,
    -- layer=1 filter=54 channel=93
    -12, -14, 0, -28, -8, 13, -15, 0, 14,
    -- layer=1 filter=54 channel=94
    -22, -28, 2, -28, 1, 12, -26, 2, 12,
    -- layer=1 filter=54 channel=95
    0, -51, -41, 5, -77, -66, -28, -97, -34,
    -- layer=1 filter=54 channel=96
    2, -34, -17, 19, -9, -22, 9, -15, -7,
    -- layer=1 filter=54 channel=97
    -25, -17, 4, -34, 0, 20, -4, -4, 16,
    -- layer=1 filter=54 channel=98
    -37, -10, 35, -21, 8, 26, 11, 14, -21,
    -- layer=1 filter=54 channel=99
    -31, -24, 19, -15, 23, 14, 0, 42, -3,
    -- layer=1 filter=54 channel=100
    -7, -12, -3, -15, -30, 4, -10, 13, 14,
    -- layer=1 filter=54 channel=101
    10, 0, -18, 4, -18, -9, -12, 0, -1,
    -- layer=1 filter=54 channel=102
    -5, -17, 0, -38, -3, 15, -53, -11, 8,
    -- layer=1 filter=54 channel=103
    -13, -39, -8, -19, -43, 12, -15, 2, 17,
    -- layer=1 filter=54 channel=104
    -31, 32, -30, -13, 6, -29, 14, 1, -11,
    -- layer=1 filter=54 channel=105
    -26, -3, 7, -32, -3, 19, -16, 9, 20,
    -- layer=1 filter=54 channel=106
    34, -7, -36, 12, -40, -38, -2, -20, -36,
    -- layer=1 filter=54 channel=107
    8, 6, 4, 12, 14, 9, 8, 13, 17,
    -- layer=1 filter=54 channel=108
    -8, 4, -41, 22, 0, -50, 10, -5, -44,
    -- layer=1 filter=54 channel=109
    -2, -9, -8, 0, 3, -1, -4, -9, -7,
    -- layer=1 filter=54 channel=110
    -19, -11, 0, -21, -10, 21, -1, 1, 18,
    -- layer=1 filter=54 channel=111
    1, -13, -26, 11, -69, -44, -54, -48, -26,
    -- layer=1 filter=54 channel=112
    -9, -45, -35, -19, -73, -69, -33, -81, 0,
    -- layer=1 filter=54 channel=113
    1, 5, -9, 16, 3, 1, 28, 8, 6,
    -- layer=1 filter=54 channel=114
    -6, -64, 25, -11, -5, -25, 0, -12, -15,
    -- layer=1 filter=54 channel=115
    -44, 16, 23, -10, 23, 34, 17, 36, 26,
    -- layer=1 filter=54 channel=116
    -8, -4, -11, -9, -10, -6, -6, -9, 7,
    -- layer=1 filter=54 channel=117
    -5, -87, -17, -68, -72, -50, -52, -58, -21,
    -- layer=1 filter=54 channel=118
    10, -8, -21, 32, -75, -57, 0, -55, -37,
    -- layer=1 filter=54 channel=119
    16, 15, -27, 39, 5, -24, 14, 5, -40,
    -- layer=1 filter=54 channel=120
    -22, 26, 9, -7, 26, 20, 9, -4, 8,
    -- layer=1 filter=54 channel=121
    -46, -17, 13, 13, 23, -10, 11, -16, 7,
    -- layer=1 filter=54 channel=122
    -7, -4, 10, 5, 1, 4, 5, 6, -2,
    -- layer=1 filter=54 channel=123
    -17, -3, 19, 4, 1, 14, 14, 16, 27,
    -- layer=1 filter=54 channel=124
    -1, 8, 13, 10, -4, 11, 1, -3, 8,
    -- layer=1 filter=54 channel=125
    13, 15, 1, 29, 18, 15, 17, 30, 34,
    -- layer=1 filter=54 channel=126
    -30, -41, 16, -49, -25, 4, -4, -1, -53,
    -- layer=1 filter=54 channel=127
    14, -2, -22, 16, -60, -75, -31, -69, -33,
    -- layer=1 filter=55 channel=0
    0, 0, 8, 8, -8, -2, -9, -5, 4,
    -- layer=1 filter=55 channel=1
    -10, -11, 8, -10, -2, 3, 6, -2, -10,
    -- layer=1 filter=55 channel=2
    5, -3, 2, 3, -1, -6, -4, -9, 7,
    -- layer=1 filter=55 channel=3
    11, -5, -1, 1, -8, 0, -1, 4, 2,
    -- layer=1 filter=55 channel=4
    -7, 5, 7, -4, -5, 4, 8, 6, 6,
    -- layer=1 filter=55 channel=5
    10, -8, -3, 6, -2, -8, 11, -2, 0,
    -- layer=1 filter=55 channel=6
    -4, 9, 7, 6, -8, 2, 3, 5, -9,
    -- layer=1 filter=55 channel=7
    -7, 6, -9, 9, 4, 2, 3, 4, -5,
    -- layer=1 filter=55 channel=8
    -1, -6, 0, 1, 0, 0, 5, -10, -6,
    -- layer=1 filter=55 channel=9
    3, -6, -5, 2, 0, 0, -9, 8, 7,
    -- layer=1 filter=55 channel=10
    -9, -11, -1, -1, 8, -8, 10, 9, -3,
    -- layer=1 filter=55 channel=11
    -10, -5, -6, -8, 6, 8, 7, -11, -12,
    -- layer=1 filter=55 channel=12
    1, -9, -4, 1, -10, -2, 4, 4, 9,
    -- layer=1 filter=55 channel=13
    -5, 4, 7, 4, 8, 2, -9, 4, 7,
    -- layer=1 filter=55 channel=14
    -1, 7, 3, 6, 8, -8, 10, -7, 6,
    -- layer=1 filter=55 channel=15
    -6, 0, -3, 2, -7, -8, 1, -7, 0,
    -- layer=1 filter=55 channel=16
    8, 5, 0, -6, -9, -1, 8, -11, 3,
    -- layer=1 filter=55 channel=17
    -1, 0, -4, 0, -10, -8, -2, 3, 3,
    -- layer=1 filter=55 channel=18
    5, 1, 1, 3, -4, 1, 7, -4, 0,
    -- layer=1 filter=55 channel=19
    8, -7, -5, -5, -6, 2, 7, -2, -4,
    -- layer=1 filter=55 channel=20
    -10, -4, -8, 2, -3, -4, 4, 3, 9,
    -- layer=1 filter=55 channel=21
    -8, -2, -8, -1, 8, -3, 3, -11, -1,
    -- layer=1 filter=55 channel=22
    -8, 7, -4, 7, -1, 4, -8, -9, -5,
    -- layer=1 filter=55 channel=23
    -5, -6, -5, 5, -6, 5, -4, 0, -7,
    -- layer=1 filter=55 channel=24
    5, 4, -9, -5, -1, -10, -10, -8, 7,
    -- layer=1 filter=55 channel=25
    7, -1, -4, -1, -7, -8, -11, 6, -9,
    -- layer=1 filter=55 channel=26
    -5, 6, -1, -11, -1, -5, -6, -11, 2,
    -- layer=1 filter=55 channel=27
    0, 5, 0, 7, 2, 2, -6, 9, 0,
    -- layer=1 filter=55 channel=28
    5, -4, -1, -8, -9, -4, 0, 0, 7,
    -- layer=1 filter=55 channel=29
    6, -9, -7, 5, -7, -2, 4, -8, -7,
    -- layer=1 filter=55 channel=30
    8, 8, -8, -5, 5, 0, -4, -7, 1,
    -- layer=1 filter=55 channel=31
    1, -10, -10, -11, -8, -10, 0, 9, 6,
    -- layer=1 filter=55 channel=32
    -3, 2, 2, -9, 0, -10, -11, -9, -7,
    -- layer=1 filter=55 channel=33
    -6, 9, 0, 0, -4, 4, 4, 6, -1,
    -- layer=1 filter=55 channel=34
    -11, 0, 2, -5, 5, -6, -1, 2, 2,
    -- layer=1 filter=55 channel=35
    -3, -8, 5, -7, 5, 3, 1, 2, 5,
    -- layer=1 filter=55 channel=36
    -6, -4, 2, -9, -5, -2, 7, 6, -10,
    -- layer=1 filter=55 channel=37
    -4, 0, -10, -1, 4, 10, -10, -7, 6,
    -- layer=1 filter=55 channel=38
    -1, -1, 4, 9, -8, -3, 8, 6, -2,
    -- layer=1 filter=55 channel=39
    -1, -11, -10, -5, 1, 1, -8, 5, -3,
    -- layer=1 filter=55 channel=40
    4, 6, -4, -4, 0, 5, -1, -7, 0,
    -- layer=1 filter=55 channel=41
    8, -5, -8, 6, 0, -11, 0, 0, -1,
    -- layer=1 filter=55 channel=42
    1, 0, -5, -9, 0, 3, 9, 2, -8,
    -- layer=1 filter=55 channel=43
    0, -1, 0, -6, -6, -9, -10, 2, 6,
    -- layer=1 filter=55 channel=44
    -10, 6, -3, -11, -10, 0, -2, 5, 1,
    -- layer=1 filter=55 channel=45
    8, -9, -5, 7, -8, -5, 4, 4, -11,
    -- layer=1 filter=55 channel=46
    -10, 5, -9, 1, 0, 10, 3, -5, 0,
    -- layer=1 filter=55 channel=47
    8, -1, -7, -5, -12, -2, 5, -6, -6,
    -- layer=1 filter=55 channel=48
    6, -7, 5, -2, 3, -7, -7, 7, 0,
    -- layer=1 filter=55 channel=49
    -2, -9, 7, -1, 6, 4, -7, 6, -3,
    -- layer=1 filter=55 channel=50
    8, -7, -9, 9, -9, -1, -3, -1, 6,
    -- layer=1 filter=55 channel=51
    8, -5, -1, -4, -6, -1, -4, 0, -4,
    -- layer=1 filter=55 channel=52
    -7, -4, 7, 4, 7, -8, 0, -8, 4,
    -- layer=1 filter=55 channel=53
    -8, 4, -9, -4, 0, -1, -9, -4, 4,
    -- layer=1 filter=55 channel=54
    -2, -5, -13, -7, -12, -3, -3, -8, -3,
    -- layer=1 filter=55 channel=55
    -4, -9, -2, -6, -2, 8, 3, 7, 2,
    -- layer=1 filter=55 channel=56
    -3, 8, -2, 3, 6, -4, 6, -8, -11,
    -- layer=1 filter=55 channel=57
    1, -5, 4, -6, 6, 4, -6, 4, 5,
    -- layer=1 filter=55 channel=58
    -7, 5, -9, -11, -2, -7, -1, -7, -4,
    -- layer=1 filter=55 channel=59
    2, -8, 3, 8, -6, 3, -3, -9, -4,
    -- layer=1 filter=55 channel=60
    -5, -2, 4, 9, -1, 6, -10, -6, 0,
    -- layer=1 filter=55 channel=61
    6, 7, -5, -1, 9, 6, -8, -5, 7,
    -- layer=1 filter=55 channel=62
    8, 3, 0, 5, 0, 6, -1, 6, -11,
    -- layer=1 filter=55 channel=63
    5, -3, -2, 6, 7, -10, 0, -9, -8,
    -- layer=1 filter=55 channel=64
    -12, 6, -2, 5, -11, -5, -9, -9, 0,
    -- layer=1 filter=55 channel=65
    -3, -1, -6, -7, -5, 0, 0, -11, 7,
    -- layer=1 filter=55 channel=66
    6, 8, 0, -11, -4, -9, -9, 4, -5,
    -- layer=1 filter=55 channel=67
    7, 9, -4, -3, 2, 2, -6, 8, -2,
    -- layer=1 filter=55 channel=68
    0, -6, -2, -4, 6, 1, -10, -3, 5,
    -- layer=1 filter=55 channel=69
    -7, -7, 1, -6, -10, 1, 3, 3, 4,
    -- layer=1 filter=55 channel=70
    -3, 2, 4, 7, 5, 6, -9, -7, -3,
    -- layer=1 filter=55 channel=71
    7, 5, 6, 4, 5, -11, 0, -7, 1,
    -- layer=1 filter=55 channel=72
    -4, -5, -5, -11, 7, -8, -10, 0, 7,
    -- layer=1 filter=55 channel=73
    -4, -5, -4, 1, 2, -1, -1, 5, 2,
    -- layer=1 filter=55 channel=74
    -11, -9, 6, 3, 4, -8, 9, 4, 1,
    -- layer=1 filter=55 channel=75
    8, 6, -3, -4, -1, -9, 11, 8, 7,
    -- layer=1 filter=55 channel=76
    1, -4, 3, 5, 0, 2, 0, 1, -8,
    -- layer=1 filter=55 channel=77
    6, 6, 2, -8, 4, -7, 5, -2, -7,
    -- layer=1 filter=55 channel=78
    6, 7, -9, 0, -11, -4, -11, -2, 3,
    -- layer=1 filter=55 channel=79
    -8, -9, -12, -7, 5, 3, 6, -3, 8,
    -- layer=1 filter=55 channel=80
    -4, 9, 6, -9, 3, -8, -11, 3, -6,
    -- layer=1 filter=55 channel=81
    -11, -10, -7, 1, 0, -5, -7, 6, -3,
    -- layer=1 filter=55 channel=82
    -2, -9, 2, 4, 2, -1, 3, -7, 0,
    -- layer=1 filter=55 channel=83
    0, 8, 5, -4, 5, -3, -5, -11, -3,
    -- layer=1 filter=55 channel=84
    6, 0, -10, -6, 3, 0, 4, -9, 0,
    -- layer=1 filter=55 channel=85
    0, 2, -10, -12, -5, -3, -8, -8, -11,
    -- layer=1 filter=55 channel=86
    1, 2, -3, 4, 3, 0, -5, -3, 6,
    -- layer=1 filter=55 channel=87
    1, 3, 8, 6, -8, -5, -2, -7, 0,
    -- layer=1 filter=55 channel=88
    -4, -8, 2, -9, -6, -2, 2, 0, 3,
    -- layer=1 filter=55 channel=89
    -4, -7, 8, -5, 8, 6, 0, -6, -5,
    -- layer=1 filter=55 channel=90
    7, -11, 2, 0, 5, -1, -4, 3, -3,
    -- layer=1 filter=55 channel=91
    -6, -5, -11, -4, -6, 0, 9, 2, -9,
    -- layer=1 filter=55 channel=92
    -9, 0, 2, -5, -5, 0, 8, 3, -8,
    -- layer=1 filter=55 channel=93
    0, -10, 1, -2, -9, 1, 0, 5, 3,
    -- layer=1 filter=55 channel=94
    3, 1, -1, -6, -8, -8, 1, 8, 5,
    -- layer=1 filter=55 channel=95
    -9, -10, -3, -6, -3, 2, -10, -7, 7,
    -- layer=1 filter=55 channel=96
    -7, -5, 4, 5, 2, -2, 6, -11, 2,
    -- layer=1 filter=55 channel=97
    -2, -1, 1, 1, -6, 7, 8, -7, -9,
    -- layer=1 filter=55 channel=98
    -7, 2, 1, -6, 5, 4, 1, 1, -5,
    -- layer=1 filter=55 channel=99
    8, 5, 3, -4, -5, -10, -4, 0, 2,
    -- layer=1 filter=55 channel=100
    -11, -10, 9, 4, 5, 8, 1, -6, -3,
    -- layer=1 filter=55 channel=101
    -11, 1, -11, 8, 0, -8, 7, -2, -11,
    -- layer=1 filter=55 channel=102
    3, -6, 2, 0, 0, -9, -4, -11, -1,
    -- layer=1 filter=55 channel=103
    3, -4, 3, -7, 6, 0, -3, 5, -2,
    -- layer=1 filter=55 channel=104
    -8, -10, -3, -7, 0, -10, 2, -6, -1,
    -- layer=1 filter=55 channel=105
    0, 3, -6, 0, -1, -1, 2, 3, 8,
    -- layer=1 filter=55 channel=106
    -2, -1, 7, 7, 3, 0, -2, 2, 7,
    -- layer=1 filter=55 channel=107
    -11, -4, 0, -2, 0, -11, -7, -6, 2,
    -- layer=1 filter=55 channel=108
    -4, -8, -4, -3, -6, -4, 5, 5, -9,
    -- layer=1 filter=55 channel=109
    -6, -2, 4, 6, -3, 2, -8, 1, 8,
    -- layer=1 filter=55 channel=110
    -7, -1, 8, -1, 6, 4, 2, -10, -2,
    -- layer=1 filter=55 channel=111
    -4, 1, -1, 3, -11, -3, -6, 4, -4,
    -- layer=1 filter=55 channel=112
    -9, -11, 0, 8, -8, -6, -8, 1, 2,
    -- layer=1 filter=55 channel=113
    4, 0, -4, -1, -1, 6, 1, -5, 3,
    -- layer=1 filter=55 channel=114
    0, 3, 6, -8, 4, 10, 8, 6, -5,
    -- layer=1 filter=55 channel=115
    -2, -6, -11, 1, -2, 2, 3, 3, -5,
    -- layer=1 filter=55 channel=116
    10, 3, 0, -1, -1, -5, -1, 2, -10,
    -- layer=1 filter=55 channel=117
    -4, 3, -2, -3, 3, -6, -7, -3, -5,
    -- layer=1 filter=55 channel=118
    -1, 3, 2, -1, 0, -1, 4, -8, -1,
    -- layer=1 filter=55 channel=119
    -10, -3, 0, 6, 2, -11, -1, -7, -2,
    -- layer=1 filter=55 channel=120
    -2, -12, 6, 5, -2, -3, 2, 8, -6,
    -- layer=1 filter=55 channel=121
    -5, 4, -9, 0, -8, 10, -11, -7, 1,
    -- layer=1 filter=55 channel=122
    -6, -6, 8, 1, -5, 10, 6, 8, -6,
    -- layer=1 filter=55 channel=123
    -10, 5, 3, -5, -4, 6, -8, 0, 4,
    -- layer=1 filter=55 channel=124
    -6, 3, -11, -6, -9, -7, 9, 6, -7,
    -- layer=1 filter=55 channel=125
    -3, 1, -2, -1, 4, 2, 2, 5, 4,
    -- layer=1 filter=55 channel=126
    3, -11, -10, -4, 4, -7, -3, 3, 4,
    -- layer=1 filter=55 channel=127
    8, 10, 8, 0, 8, 7, -2, 3, -8,
    -- layer=1 filter=56 channel=0
    3, 15, -13, 15, -3, -6, 22, 5, -4,
    -- layer=1 filter=56 channel=1
    -6, -2, 4, 23, -19, 2, 16, 3, 7,
    -- layer=1 filter=56 channel=2
    -20, -8, -3, 3, -10, -2, -23, -7, -11,
    -- layer=1 filter=56 channel=3
    -3, -7, 0, -12, 12, -9, 0, 7, 6,
    -- layer=1 filter=56 channel=4
    0, -7, -2, 0, -1, 1, -7, 2, 1,
    -- layer=1 filter=56 channel=5
    9, 3, 7, 8, -19, 15, 17, -5, -7,
    -- layer=1 filter=56 channel=6
    -19, 3, 13, 2, 13, 7, -9, -22, -4,
    -- layer=1 filter=56 channel=7
    4, -34, -12, -24, -28, -17, -17, -27, -15,
    -- layer=1 filter=56 channel=8
    -7, -1, -8, 11, -26, 12, 19, 1, -2,
    -- layer=1 filter=56 channel=9
    5, -12, -14, 4, 4, 20, 45, 13, 0,
    -- layer=1 filter=56 channel=10
    0, 0, -27, 5, -20, -14, -22, 4, -27,
    -- layer=1 filter=56 channel=11
    -3, -15, -20, -17, -31, -19, -20, -10, -2,
    -- layer=1 filter=56 channel=12
    -41, -15, -19, -36, -40, -27, 17, -2, -26,
    -- layer=1 filter=56 channel=13
    -21, -19, -14, -8, -29, -20, -2, -19, -8,
    -- layer=1 filter=56 channel=14
    -13, -13, -24, -8, -42, -37, 10, -8, -20,
    -- layer=1 filter=56 channel=15
    1, -31, -3, -21, -5, -27, -11, -36, -45,
    -- layer=1 filter=56 channel=16
    8, 2, 2, 1, -9, 33, 4, 8, -9,
    -- layer=1 filter=56 channel=17
    -24, -37, -38, -38, -61, -48, -32, -44, -51,
    -- layer=1 filter=56 channel=18
    0, -7, -7, -36, -24, -23, -18, -28, -20,
    -- layer=1 filter=56 channel=19
    27, -2, 25, 16, 60, 57, 52, 20, 35,
    -- layer=1 filter=56 channel=20
    -13, -24, -18, -21, -20, -21, -35, -28, -28,
    -- layer=1 filter=56 channel=21
    4, 19, 11, 18, 44, 14, 11, 23, 27,
    -- layer=1 filter=56 channel=22
    -40, -48, -20, -40, -71, -32, -35, -59, -25,
    -- layer=1 filter=56 channel=23
    46, -6, 24, -8, -1, -30, 6, -3, -1,
    -- layer=1 filter=56 channel=24
    19, 24, 12, 18, 27, 52, 35, 19, 27,
    -- layer=1 filter=56 channel=25
    -6, 4, -1, -17, -8, 5, -16, 12, 0,
    -- layer=1 filter=56 channel=26
    9, -22, -29, 3, -29, -7, -8, -34, -12,
    -- layer=1 filter=56 channel=27
    21, 13, 13, 36, 16, 14, 28, 16, 22,
    -- layer=1 filter=56 channel=28
    -23, -7, -24, 12, 1, 1, 18, 29, 15,
    -- layer=1 filter=56 channel=29
    -7, -25, -34, -4, -18, -25, -26, -34, -30,
    -- layer=1 filter=56 channel=30
    27, 18, 2, 23, 17, 28, 52, 18, 11,
    -- layer=1 filter=56 channel=31
    -55, -48, -25, -74, -70, -90, -29, -52, -56,
    -- layer=1 filter=56 channel=32
    6, 3, 0, 9, 1, -14, 13, -17, -18,
    -- layer=1 filter=56 channel=33
    2, -11, -10, -15, -11, -18, 0, -9, 7,
    -- layer=1 filter=56 channel=34
    -25, -32, -11, -23, -27, -16, -21, -25, -14,
    -- layer=1 filter=56 channel=35
    5, 5, 14, 5, 6, 3, 3, 7, 12,
    -- layer=1 filter=56 channel=36
    -21, -5, 1, -6, -25, 0, -9, -5, 10,
    -- layer=1 filter=56 channel=37
    17, 6, 32, 4, 10, 24, 4, -8, -10,
    -- layer=1 filter=56 channel=38
    -3, 5, -2, 5, -5, -8, -7, 9, -5,
    -- layer=1 filter=56 channel=39
    3, 8, -2, 8, 1, -1, 15, 9, 15,
    -- layer=1 filter=56 channel=40
    -29, -40, -6, -37, -45, -26, -50, -64, -42,
    -- layer=1 filter=56 channel=41
    3, -2, -24, 6, 15, 3, 3, 2, 24,
    -- layer=1 filter=56 channel=42
    -33, -29, -20, -12, -18, -8, -29, -35, -36,
    -- layer=1 filter=56 channel=43
    27, 16, 0, 18, -9, 15, 23, -4, 16,
    -- layer=1 filter=56 channel=44
    6, -19, -21, 11, -18, 4, 5, -21, -22,
    -- layer=1 filter=56 channel=45
    13, 21, -5, 13, 11, 15, 2, 14, 9,
    -- layer=1 filter=56 channel=46
    16, 1, -15, -4, 21, 0, 6, -6, -12,
    -- layer=1 filter=56 channel=47
    12, 10, 19, -23, 16, -27, 3, 5, -24,
    -- layer=1 filter=56 channel=48
    19, 9, 8, 9, 19, 19, 13, 22, 16,
    -- layer=1 filter=56 channel=49
    19, 21, 9, 9, 18, 20, 8, 16, 11,
    -- layer=1 filter=56 channel=50
    6, -1, 0, 0, -11, 12, -4, 1, -1,
    -- layer=1 filter=56 channel=51
    11, 5, 8, 11, 21, 1, 14, 19, 15,
    -- layer=1 filter=56 channel=52
    1, -1, 4, 17, 10, 16, -14, -31, 6,
    -- layer=1 filter=56 channel=53
    -11, 0, -14, 1, -10, -10, -7, -17, -13,
    -- layer=1 filter=56 channel=54
    28, 8, 23, 5, 1, 27, -1, 24, 10,
    -- layer=1 filter=56 channel=55
    -12, -14, 5, 1, -24, 1, -6, 0, 10,
    -- layer=1 filter=56 channel=56
    -6, 4, -2, 6, 1, -14, -14, -14, 0,
    -- layer=1 filter=56 channel=57
    -35, -62, -50, -21, -73, -42, -50, -46, -49,
    -- layer=1 filter=56 channel=58
    32, -6, -5, -15, -15, 12, -11, -2, -13,
    -- layer=1 filter=56 channel=59
    7, 5, 2, -3, -9, 11, 4, 4, 6,
    -- layer=1 filter=56 channel=60
    -1, -17, -16, -14, -6, -8, -2, -15, -4,
    -- layer=1 filter=56 channel=61
    5, 3, 9, 2, 0, 1, -4, -2, -3,
    -- layer=1 filter=56 channel=62
    0, 0, -18, 8, -16, 27, 8, -1, 0,
    -- layer=1 filter=56 channel=63
    2, -1, 16, 6, 22, 12, 18, 20, 37,
    -- layer=1 filter=56 channel=64
    -15, -5, -3, 1, -13, -10, -4, 8, 11,
    -- layer=1 filter=56 channel=65
    19, 10, -8, 22, 28, 12, 12, 16, -2,
    -- layer=1 filter=56 channel=66
    9, 11, 24, 14, 4, 10, 15, 20, 19,
    -- layer=1 filter=56 channel=67
    6, 12, -9, 1, 2, 7, -17, -4, -9,
    -- layer=1 filter=56 channel=68
    1, 4, -8, 4, 1, 26, -5, 3, 11,
    -- layer=1 filter=56 channel=69
    13, -28, -4, 5, -24, 18, -11, -17, -16,
    -- layer=1 filter=56 channel=70
    0, 13, 26, 18, 3, 8, -12, -25, 0,
    -- layer=1 filter=56 channel=71
    16, 16, 7, 46, 45, 24, 35, 34, 23,
    -- layer=1 filter=56 channel=72
    -8, -13, -3, 27, -2, 31, 25, -25, 2,
    -- layer=1 filter=56 channel=73
    6, -1, 7, 8, 3, 5, -1, 8, 16,
    -- layer=1 filter=56 channel=74
    7, 6, -3, -3, 3, 10, 7, -12, 8,
    -- layer=1 filter=56 channel=75
    14, -2, 20, -30, 14, -9, 11, -1, -1,
    -- layer=1 filter=56 channel=76
    7, 2, 9, 6, 0, 0, 12, 3, 3,
    -- layer=1 filter=56 channel=77
    7, 23, 0, 29, 35, 24, 19, 24, 20,
    -- layer=1 filter=56 channel=78
    -17, -9, -14, -8, -7, -2, -21, -6, -24,
    -- layer=1 filter=56 channel=79
    4, -9, 1, 2, -9, 8, 0, 0, 6,
    -- layer=1 filter=56 channel=80
    -5, 0, -23, -3, -13, -4, -5, -11, -6,
    -- layer=1 filter=56 channel=81
    2, 16, 0, 32, 50, 28, 17, 35, 21,
    -- layer=1 filter=56 channel=82
    8, 17, 2, 42, 49, 31, 23, 42, 20,
    -- layer=1 filter=56 channel=83
    3, -11, 3, 10, -6, 0, 11, 2, -8,
    -- layer=1 filter=56 channel=84
    4, 24, 13, 11, 21, 5, -8, 2, 9,
    -- layer=1 filter=56 channel=85
    25, -5, 12, -18, 16, 3, -9, -3, 5,
    -- layer=1 filter=56 channel=86
    -27, -36, -22, -30, -58, -47, -22, -50, -22,
    -- layer=1 filter=56 channel=87
    -22, -18, -8, -39, 9, -5, 4, 7, -3,
    -- layer=1 filter=56 channel=88
    4, 10, -8, 5, 6, -1, -9, -1, 2,
    -- layer=1 filter=56 channel=89
    22, 19, 26, 36, 38, 25, 4, 30, 9,
    -- layer=1 filter=56 channel=90
    -13, -33, -42, 13, -32, 17, 8, -16, -4,
    -- layer=1 filter=56 channel=91
    -2, -9, 4, -13, -8, -11, -21, -7, -16,
    -- layer=1 filter=56 channel=92
    32, 9, -16, -14, 2, -26, -22, 23, -21,
    -- layer=1 filter=56 channel=93
    21, 18, 23, 39, 34, 28, 31, 34, 24,
    -- layer=1 filter=56 channel=94
    -19, -12, -3, -17, -16, -21, -15, -16, -17,
    -- layer=1 filter=56 channel=95
    21, 14, 29, 15, 21, 29, 23, 32, 24,
    -- layer=1 filter=56 channel=96
    -9, -4, 5, -2, -3, -5, 0, -12, -3,
    -- layer=1 filter=56 channel=97
    8, 8, -2, 19, 4, 15, 15, 4, 15,
    -- layer=1 filter=56 channel=98
    5, 7, 1, 5, -3, 3, 18, 7, 0,
    -- layer=1 filter=56 channel=99
    -5, 20, -13, 20, 4, 7, 30, 25, 12,
    -- layer=1 filter=56 channel=100
    -2, -15, -2, -11, 13, -1, 12, 1, 12,
    -- layer=1 filter=56 channel=101
    0, 1, -1, 4, 3, 2, 11, 1, 5,
    -- layer=1 filter=56 channel=102
    -8, -27, -27, -20, -26, -27, -14, -19, -14,
    -- layer=1 filter=56 channel=103
    1, -3, -6, 17, 3, 10, -20, -11, -1,
    -- layer=1 filter=56 channel=104
    21, 9, -9, -17, -27, -56, 0, 5, -31,
    -- layer=1 filter=56 channel=105
    -5, 8, 2, 9, -1, 1, 17, 9, 16,
    -- layer=1 filter=56 channel=106
    -13, -4, -3, 12, -9, 0, -14, 7, -7,
    -- layer=1 filter=56 channel=107
    2, 9, -8, 8, 0, 12, -9, -15, -1,
    -- layer=1 filter=56 channel=108
    17, -6, -10, 6, -3, 7, 9, -1, -6,
    -- layer=1 filter=56 channel=109
    -7, 9, 5, -4, 0, 1, -7, -11, 4,
    -- layer=1 filter=56 channel=110
    8, 3, 3, -4, 3, -7, -5, 7, -8,
    -- layer=1 filter=56 channel=111
    13, 13, 0, 12, 12, 22, 26, 8, 18,
    -- layer=1 filter=56 channel=112
    27, 14, 37, 19, 5, -5, -8, 19, 9,
    -- layer=1 filter=56 channel=113
    -5, -14, -19, 7, -13, 3, 0, -38, -8,
    -- layer=1 filter=56 channel=114
    -6, -6, -1, -9, -27, -6, -7, -15, -17,
    -- layer=1 filter=56 channel=115
    -19, -32, -31, -36, -53, -50, -44, -39, -52,
    -- layer=1 filter=56 channel=116
    -4, 3, -2, 1, 0, -3, -9, 7, -11,
    -- layer=1 filter=56 channel=117
    26, 11, -5, 40, -15, 2, -11, 0, -31,
    -- layer=1 filter=56 channel=118
    4, 25, 1, 3, 12, 22, 21, 5, 4,
    -- layer=1 filter=56 channel=119
    -1, 6, -17, 8, -5, 20, 14, 15, 16,
    -- layer=1 filter=56 channel=120
    14, 6, 0, 14, 23, 18, -4, 15, 16,
    -- layer=1 filter=56 channel=121
    -9, -11, -21, 2, -15, 5, 46, 30, -4,
    -- layer=1 filter=56 channel=122
    -1, 4, -8, 9, -2, 2, 2, -3, 5,
    -- layer=1 filter=56 channel=123
    7, -4, 4, -12, -2, 13, 12, 13, 1,
    -- layer=1 filter=56 channel=124
    -10, -3, -22, -15, -14, -3, -13, -5, -17,
    -- layer=1 filter=56 channel=125
    16, 32, 22, 38, 22, 2, 18, -5, 15,
    -- layer=1 filter=56 channel=126
    -1, 10, 17, 26, -10, -4, 16, 23, 18,
    -- layer=1 filter=56 channel=127
    15, 11, 23, 5, 16, 9, 21, 10, 3,
    -- layer=1 filter=57 channel=0
    -16, -9, -3, -18, -13, -10, -38, -18, 45,
    -- layer=1 filter=57 channel=1
    -66, -35, -41, -13, -7, -9, 0, -18, 54,
    -- layer=1 filter=57 channel=2
    -27, 3, -17, 4, 15, -95, -14, -32, -96,
    -- layer=1 filter=57 channel=3
    6, -4, -8, -6, 6, -10, 0, -5, 3,
    -- layer=1 filter=57 channel=4
    13, 1, 3, 8, 3, 7, 11, -4, -8,
    -- layer=1 filter=57 channel=5
    -52, -80, -49, 14, -24, -4, -9, -5, 38,
    -- layer=1 filter=57 channel=6
    0, -69, -68, -89, -120, -90, -111, -43, -4,
    -- layer=1 filter=57 channel=7
    -82, -28, 72, -11, -21, 69, -15, 61, 110,
    -- layer=1 filter=57 channel=8
    -69, -74, -15, -8, -4, 0, 5, 2, 55,
    -- layer=1 filter=57 channel=9
    -10, 33, -22, 8, -15, -28, -36, -13, -7,
    -- layer=1 filter=57 channel=10
    -33, -39, 64, -15, -26, 88, -38, 57, 105,
    -- layer=1 filter=57 channel=11
    5, -9, 16, -5, -1, 6, -8, -5, 10,
    -- layer=1 filter=57 channel=12
    14, 6, -66, -28, -64, -67, -36, -52, -58,
    -- layer=1 filter=57 channel=13
    -56, -40, -41, -58, -42, -23, -56, -18, -44,
    -- layer=1 filter=57 channel=14
    -32, -5, 44, -13, -74, 38, -2, -36, 56,
    -- layer=1 filter=57 channel=15
    -39, -75, -25, -12, -42, -32, -7, -11, -57,
    -- layer=1 filter=57 channel=16
    -39, -84, -1, 17, -9, 32, -17, 27, 60,
    -- layer=1 filter=57 channel=17
    -65, -55, -68, -100, -44, -28, -57, -40, 5,
    -- layer=1 filter=57 channel=18
    33, 22, 12, 15, -76, -111, -46, -46, -82,
    -- layer=1 filter=57 channel=19
    48, 35, 5, 10, -27, 30, -67, 24, -17,
    -- layer=1 filter=57 channel=20
    -72, -34, -7, -44, -28, -12, -33, 5, 37,
    -- layer=1 filter=57 channel=21
    -7, -2, -9, 0, -1, 7, 39, 12, 70,
    -- layer=1 filter=57 channel=22
    -89, -34, -7, -15, -28, 0, -23, -3, 48,
    -- layer=1 filter=57 channel=23
    -66, -94, 65, -21, -5, 78, -10, 64, 51,
    -- layer=1 filter=57 channel=24
    -6, -2, -26, 1, 13, -24, 10, 20, -66,
    -- layer=1 filter=57 channel=25
    -46, -52, 54, 10, 5, 92, -17, 49, 117,
    -- layer=1 filter=57 channel=26
    -101, -44, -72, -95, -69, -45, -99, -30, -72,
    -- layer=1 filter=57 channel=27
    22, 44, 0, 54, 59, 11, 41, 25, -11,
    -- layer=1 filter=57 channel=28
    -81, -36, 34, -23, -23, 64, -28, 29, 97,
    -- layer=1 filter=57 channel=29
    -10, 12, -25, 29, 21, -11, -1, 0, -2,
    -- layer=1 filter=57 channel=30
    61, 36, -1, 14, -43, -69, -61, -39, -38,
    -- layer=1 filter=57 channel=31
    37, 13, -31, -27, -72, -42, -92, -104, -85,
    -- layer=1 filter=57 channel=32
    -58, -42, -73, -95, -70, -25, -140, -11, -46,
    -- layer=1 filter=57 channel=33
    -4, 0, 18, 3, -48, 7, 4, 28, 43,
    -- layer=1 filter=57 channel=34
    16, -24, -37, 0, -37, 1, -13, -24, 6,
    -- layer=1 filter=57 channel=35
    -8, -16, -24, -16, -31, -15, -11, -3, -17,
    -- layer=1 filter=57 channel=36
    11, -1, 5, 5, 0, 26, -20, -28, 3,
    -- layer=1 filter=57 channel=37
    -11, -90, -2, 14, -13, 37, -11, 44, 29,
    -- layer=1 filter=57 channel=38
    -17, -9, -10, -34, -15, -1, -20, 4, 5,
    -- layer=1 filter=57 channel=39
    -5, -2, 21, 15, 35, 65, -3, 20, 35,
    -- layer=1 filter=57 channel=40
    29, -33, -31, -57, -117, -62, -60, -77, -28,
    -- layer=1 filter=57 channel=41
    12, -7, 1, -5, -16, 36, -77, 9, 21,
    -- layer=1 filter=57 channel=42
    -20, -29, 2, 5, 20, -27, -29, -23, -48,
    -- layer=1 filter=57 channel=43
    -64, -86, 52, 22, 12, 56, 17, 37, 75,
    -- layer=1 filter=57 channel=44
    -102, -50, -82, -134, -89, -17, -99, -34, -44,
    -- layer=1 filter=57 channel=45
    -51, -39, -16, -27, -26, -60, -13, -10, -34,
    -- layer=1 filter=57 channel=46
    48, -5, 35, 9, 0, -15, -43, 28, -57,
    -- layer=1 filter=57 channel=47
    -17, -46, 51, -41, 32, -18, -48, 37, -43,
    -- layer=1 filter=57 channel=48
    -17, -29, 2, -34, -34, 39, 9, 5, 30,
    -- layer=1 filter=57 channel=49
    -13, -30, -15, -51, -7, -3, -32, -23, -10,
    -- layer=1 filter=57 channel=50
    -43, 27, -15, 17, 29, 0, 14, 26, -6,
    -- layer=1 filter=57 channel=51
    -28, -23, 36, -4, -47, 50, 6, 11, 79,
    -- layer=1 filter=57 channel=52
    -43, -43, 12, 7, -2, 11, 22, 47, 20,
    -- layer=1 filter=57 channel=53
    -19, -14, -18, -3, -7, -22, -19, -16, -7,
    -- layer=1 filter=57 channel=54
    0, -52, 82, 21, 29, 96, -16, 85, 111,
    -- layer=1 filter=57 channel=55
    9, 10, 3, 16, 26, -3, 32, 16, -21,
    -- layer=1 filter=57 channel=56
    -11, -12, -6, 7, 5, 2, -12, -6, 0,
    -- layer=1 filter=57 channel=57
    -27, -45, 38, -32, -31, 73, -29, 38, 82,
    -- layer=1 filter=57 channel=58
    -33, -47, 109, -33, 29, 114, -7, 121, 91,
    -- layer=1 filter=57 channel=59
    -12, 7, -2, -9, -16, 2, -20, -10, 4,
    -- layer=1 filter=57 channel=60
    8, 24, 21, 34, 6, 3, 26, 22, 5,
    -- layer=1 filter=57 channel=61
    2, 1, 1, 1, -10, 1, -8, -3, 6,
    -- layer=1 filter=57 channel=62
    -62, -91, 12, 4, -19, 40, -7, 36, 58,
    -- layer=1 filter=57 channel=63
    23, 5, 17, 17, -2, -13, -27, -14, -34,
    -- layer=1 filter=57 channel=64
    -50, -41, -19, -42, -10, 0, -49, -34, 35,
    -- layer=1 filter=57 channel=65
    -53, -32, -20, -33, -31, 0, -9, 5, 32,
    -- layer=1 filter=57 channel=66
    7, 15, 33, -6, 2, 22, -13, -25, 28,
    -- layer=1 filter=57 channel=67
    -52, -45, -45, -98, -27, -22, -36, -31, -9,
    -- layer=1 filter=57 channel=68
    -76, -61, -33, -124, -56, 26, -119, -35, -31,
    -- layer=1 filter=57 channel=69
    -55, -66, -42, -2, -40, -31, -16, 7, -39,
    -- layer=1 filter=57 channel=70
    -31, -45, -67, -117, -66, -35, -87, -60, 42,
    -- layer=1 filter=57 channel=71
    1, 27, 19, 47, 23, 47, 46, 43, 46,
    -- layer=1 filter=57 channel=72
    52, 31, 19, 19, -37, -28, -38, 9, -9,
    -- layer=1 filter=57 channel=73
    -9, -4, -1, -8, -9, -6, 6, -7, 0,
    -- layer=1 filter=57 channel=74
    54, -12, -3, -71, -7, 68, -123, -2, -1,
    -- layer=1 filter=57 channel=75
    38, 36, -1, 20, -39, -59, -19, -45, -71,
    -- layer=1 filter=57 channel=76
    -42, -33, -23, -77, -42, -10, -52, -31, -3,
    -- layer=1 filter=57 channel=77
    -23, -7, -23, -15, -6, -4, 8, -6, 35,
    -- layer=1 filter=57 channel=78
    -30, -10, -8, -42, -15, -3, -35, -6, 27,
    -- layer=1 filter=57 channel=79
    -54, -96, 8, 0, -11, 46, -20, 49, 37,
    -- layer=1 filter=57 channel=80
    -6, -39, -18, -20, -40, 27, 22, -4, 10,
    -- layer=1 filter=57 channel=81
    5, -17, -10, 20, 25, 39, 24, 35, 7,
    -- layer=1 filter=57 channel=82
    4, 3, -2, -9, 0, 5, 20, 8, 17,
    -- layer=1 filter=57 channel=83
    -81, -61, 31, -58, -62, -45, 0, -49, -24,
    -- layer=1 filter=57 channel=84
    14, 7, -4, -26, -60, -46, -86, 6, -45,
    -- layer=1 filter=57 channel=85
    -39, -25, 78, -70, 59, 95, -13, 115, 57,
    -- layer=1 filter=57 channel=86
    -39, -7, 15, -25, -13, 22, -27, -23, 32,
    -- layer=1 filter=57 channel=87
    48, 58, 28, -4, -3, 3, -42, 5, 10,
    -- layer=1 filter=57 channel=88
    -30, -48, -18, -37, -38, 13, -25, -12, -16,
    -- layer=1 filter=57 channel=89
    -15, -5, -31, -34, -16, -44, 2, 0, 10,
    -- layer=1 filter=57 channel=90
    -104, -72, -58, -116, -60, -17, -94, -40, -37,
    -- layer=1 filter=57 channel=91
    -31, -22, 3, -38, -32, 5, -29, -5, 28,
    -- layer=1 filter=57 channel=92
    -64, -45, -10, -79, -92, -63, -62, -3, -62,
    -- layer=1 filter=57 channel=93
    -8, -9, -12, -12, 0, 5, 1, -2, 37,
    -- layer=1 filter=57 channel=94
    -31, -25, 18, -37, -27, 2, -58, -23, 18,
    -- layer=1 filter=57 channel=95
    30, -1, 6, -13, -28, -62, -74, -8, -50,
    -- layer=1 filter=57 channel=96
    11, 24, 16, -7, 10, -36, 5, -15, -8,
    -- layer=1 filter=57 channel=97
    -50, -16, 4, -34, -29, 13, -30, -3, 39,
    -- layer=1 filter=57 channel=98
    -66, -85, 28, 7, 3, 64, -8, 38, 76,
    -- layer=1 filter=57 channel=99
    -20, -68, -10, -20, -73, 42, -21, -25, 90,
    -- layer=1 filter=57 channel=100
    11, 6, 18, 4, -2, -15, -11, -15, -10,
    -- layer=1 filter=57 channel=101
    -30, -22, -19, -47, -29, -8, -18, -15, 21,
    -- layer=1 filter=57 channel=102
    -19, -29, -23, -89, -55, -55, -88, -42, -18,
    -- layer=1 filter=57 channel=103
    28, -4, 11, 6, -6, -9, -13, 4, 10,
    -- layer=1 filter=57 channel=104
    -2, -32, -7, -32, -2, 76, -28, 18, 6,
    -- layer=1 filter=57 channel=105
    -4, -11, 22, -33, -18, 32, -23, -13, 45,
    -- layer=1 filter=57 channel=106
    -36, -33, -41, -102, -50, -53, -100, 2, -14,
    -- layer=1 filter=57 channel=107
    4, 1, 10, 12, 12, 5, 15, 6, 8,
    -- layer=1 filter=57 channel=108
    -94, -75, -69, -94, -75, -48, -76, -26, -50,
    -- layer=1 filter=57 channel=109
    2, 4, 0, 1, 3, 3, 7, -8, -6,
    -- layer=1 filter=57 channel=110
    -9, -14, -12, -12, -15, 3, -11, 0, 16,
    -- layer=1 filter=57 channel=111
    39, 25, 6, 12, -55, -97, -52, -24, -51,
    -- layer=1 filter=57 channel=112
    29, 12, -5, 26, -25, -39, -38, -3, -25,
    -- layer=1 filter=57 channel=113
    -31, -39, 31, -18, -16, 32, -65, -20, 16,
    -- layer=1 filter=57 channel=114
    -31, -41, -65, 24, -12, 2, 11, 0, -11,
    -- layer=1 filter=57 channel=115
    -50, -37, 39, -9, -22, 52, -43, 17, 73,
    -- layer=1 filter=57 channel=116
    -7, -8, -9, -3, -9, 9, -3, 1, 8,
    -- layer=1 filter=57 channel=117
    45, 16, 7, 13, -88, -53, -6, -33, -21,
    -- layer=1 filter=57 channel=118
    34, 12, 0, -22, -29, -58, -124, -1, -57,
    -- layer=1 filter=57 channel=119
    -74, -46, -62, -89, -52, -23, -103, -3, -45,
    -- layer=1 filter=57 channel=120
    -18, -40, 26, -3, -2, 54, 19, 44, 85,
    -- layer=1 filter=57 channel=121
    62, 51, 13, 51, 11, -36, 1, -32, -58,
    -- layer=1 filter=57 channel=122
    1, -9, -4, -9, 4, 3, -10, 9, -6,
    -- layer=1 filter=57 channel=123
    33, 39, 42, 45, 31, 7, 18, 10, -3,
    -- layer=1 filter=57 channel=124
    -1, 25, 7, 16, 11, 1, 2, 0, -16,
    -- layer=1 filter=57 channel=125
    -15, -66, -58, -144, -128, -38, -74, -54, 9,
    -- layer=1 filter=57 channel=126
    -93, -44, 15, -46, -23, -24, -8, -7, 36,
    -- layer=1 filter=57 channel=127
    39, 18, 7, -4, -40, -84, -90, -28, -69,
    -- layer=1 filter=58 channel=0
    -22, -47, -4, -26, -29, -7, -52, -57, -32,
    -- layer=1 filter=58 channel=1
    12, -18, 9, -27, -30, 0, -15, -28, -25,
    -- layer=1 filter=58 channel=2
    -10, 51, 51, 7, 42, 58, 46, 57, 75,
    -- layer=1 filter=58 channel=3
    3, 9, 10, -4, -2, 3, 3, -5, 14,
    -- layer=1 filter=58 channel=4
    0, 5, -7, -1, 7, 9, 5, 5, 6,
    -- layer=1 filter=58 channel=5
    -20, -59, -15, -74, -72, -16, -34, -30, -30,
    -- layer=1 filter=58 channel=6
    7, -62, -73, 2, -67, -77, -36, -59, -80,
    -- layer=1 filter=58 channel=7
    -53, -55, 29, -94, 2, 32, -43, 21, 23,
    -- layer=1 filter=58 channel=8
    -50, -70, -41, -117, -80, 0, -49, -75, -74,
    -- layer=1 filter=58 channel=9
    80, 88, 42, 155, 110, 74, 81, 14, 96,
    -- layer=1 filter=58 channel=10
    -63, -56, 36, -87, 1, 45, -32, 5, -2,
    -- layer=1 filter=58 channel=11
    17, -51, -60, -1, -49, -51, -11, -59, -11,
    -- layer=1 filter=58 channel=12
    -34, -66, 22, 82, 7, 30, -3, 24, 25,
    -- layer=1 filter=58 channel=13
    8, -5, -39, 3, -31, -45, -32, -79, -45,
    -- layer=1 filter=58 channel=14
    -12, -80, 42, -53, 0, 23, -31, -23, 19,
    -- layer=1 filter=58 channel=15
    -39, -9, -49, -24, -37, -41, -7, -7, 0,
    -- layer=1 filter=58 channel=16
    -51, -56, -11, -97, -60, 7, -52, -44, -65,
    -- layer=1 filter=58 channel=17
    19, -11, -13, -63, -43, 1, -79, -80, -33,
    -- layer=1 filter=58 channel=18
    29, -30, -35, 65, 2, -28, -31, -54, 42,
    -- layer=1 filter=58 channel=19
    -6, 28, -23, 58, 35, -27, -2, 24, 18,
    -- layer=1 filter=58 channel=20
    -18, -46, -49, -61, -67, -67, -52, -62, -63,
    -- layer=1 filter=58 channel=21
    34, 31, 25, 25, 35, 38, 20, 23, 11,
    -- layer=1 filter=58 channel=22
    -2, -72, -44, -23, -93, -60, -41, -51, -56,
    -- layer=1 filter=58 channel=23
    12, 62, 3, -10, 6, -15, -27, 40, 23,
    -- layer=1 filter=58 channel=24
    41, 68, 43, 60, 55, 47, 37, 27, 30,
    -- layer=1 filter=58 channel=25
    -57, -38, 20, -50, -11, 53, -37, 9, 0,
    -- layer=1 filter=58 channel=26
    48, 40, -33, 39, -20, -57, -10, -102, -19,
    -- layer=1 filter=58 channel=27
    10, 24, 31, 50, 24, 31, 38, 23, 10,
    -- layer=1 filter=58 channel=28
    -28, -53, 30, -42, 5, 61, -13, 13, 15,
    -- layer=1 filter=58 channel=29
    27, 17, 20, 22, 23, 25, 22, 8, 13,
    -- layer=1 filter=58 channel=30
    60, 26, -19, 108, 31, -16, 18, -42, 9,
    -- layer=1 filter=58 channel=31
    -4, -50, -39, 35, -12, -18, 12, 13, 38,
    -- layer=1 filter=58 channel=32
    57, 63, -39, 55, -3, -20, 9, -71, 8,
    -- layer=1 filter=58 channel=33
    -4, -16, -43, 16, 6, -55, 6, 7, -27,
    -- layer=1 filter=58 channel=34
    31, 4, -10, 28, -20, -32, 40, -35, -3,
    -- layer=1 filter=58 channel=35
    10, 0, 0, 0, -8, -2, 10, 3, 8,
    -- layer=1 filter=58 channel=36
    0, -51, -53, -23, -63, -29, -36, -79, -17,
    -- layer=1 filter=58 channel=37
    -54, -56, 2, -61, -24, 12, -44, -20, -45,
    -- layer=1 filter=58 channel=38
    0, -16, -18, 11, 0, -20, -1, -21, -31,
    -- layer=1 filter=58 channel=39
    -21, -43, -24, -47, -69, -22, -9, -34, -21,
    -- layer=1 filter=58 channel=40
    -13, -70, -56, 24, -40, -35, -57, -57, -26,
    -- layer=1 filter=58 channel=41
    75, 78, -44, 92, 42, 9, 36, -53, 28,
    -- layer=1 filter=58 channel=42
    -18, 12, 54, 6, 20, 49, 41, 47, 59,
    -- layer=1 filter=58 channel=43
    -4, -7, 18, -8, -6, 45, -22, 4, -26,
    -- layer=1 filter=58 channel=44
    42, 36, -22, 27, -41, -16, -12, -99, -7,
    -- layer=1 filter=58 channel=45
    11, 15, 10, 0, 18, 19, 9, -19, -3,
    -- layer=1 filter=58 channel=46
    -40, -41, -51, -14, 15, -1, 3, 30, 52,
    -- layer=1 filter=58 channel=47
    7, 52, 1, 17, 10, -5, 1, -2, 6,
    -- layer=1 filter=58 channel=48
    -7, 5, -1, 8, 20, 8, 13, 10, 8,
    -- layer=1 filter=58 channel=49
    15, 33, 19, 31, 27, 17, 19, 15, 27,
    -- layer=1 filter=58 channel=50
    -17, 11, -5, 38, 24, -16, -7, -16, 1,
    -- layer=1 filter=58 channel=51
    -19, 9, 15, -8, 28, 13, 5, 19, -4,
    -- layer=1 filter=58 channel=52
    -33, -10, 1, -6, 9, 7, -8, -17, -13,
    -- layer=1 filter=58 channel=53
    4, 1, 14, 1, 0, 19, 5, 9, -3,
    -- layer=1 filter=58 channel=54
    -45, 6, 35, -2, 23, 51, -12, 39, -11,
    -- layer=1 filter=58 channel=55
    -26, -30, -46, -21, -20, -9, -4, -24, -23,
    -- layer=1 filter=58 channel=56
    -6, 4, -1, 3, 0, 15, 0, 0, -10,
    -- layer=1 filter=58 channel=57
    -61, -88, 27, -72, -31, 35, -49, -8, -15,
    -- layer=1 filter=58 channel=58
    -43, 20, 16, -16, 44, 40, -9, 60, 32,
    -- layer=1 filter=58 channel=59
    -2, -10, -15, -18, -2, 8, -10, -13, 5,
    -- layer=1 filter=58 channel=60
    -14, -3, -10, 1, -1, 26, -29, 34, -2,
    -- layer=1 filter=58 channel=61
    15, 0, -1, -11, 3, 0, -8, -3, 8,
    -- layer=1 filter=58 channel=62
    -64, -24, -20, -102, -64, -3, -60, -19, -62,
    -- layer=1 filter=58 channel=63
    -1, -38, -38, 30, -49, -13, -33, -51, -20,
    -- layer=1 filter=58 channel=64
    6, -26, -11, -8, 6, -1, -20, -9, -26,
    -- layer=1 filter=58 channel=65
    9, 20, 8, 2, 21, 3, 10, 12, -2,
    -- layer=1 filter=58 channel=66
    -12, -27, -11, -29, -17, 2, -22, -12, 0,
    -- layer=1 filter=58 channel=67
    61, 9, 8, 45, 37, 0, 35, 33, 14,
    -- layer=1 filter=58 channel=68
    48, 30, -11, 45, -42, 25, -14, -98, 4,
    -- layer=1 filter=58 channel=69
    -37, 0, -24, -49, -59, -42, -23, -43, -40,
    -- layer=1 filter=58 channel=70
    -3, -79, -38, -24, -38, -63, -3, -41, -46,
    -- layer=1 filter=58 channel=71
    28, 43, 30, 24, 50, 22, 30, 50, 19,
    -- layer=1 filter=58 channel=72
    11, -10, -56, 91, 31, -39, -5, -47, 12,
    -- layer=1 filter=58 channel=73
    -1, -11, -9, 4, 7, 6, 12, -2, 6,
    -- layer=1 filter=58 channel=74
    42, -6, -33, 69, -43, 21, -59, -55, -5,
    -- layer=1 filter=58 channel=75
    22, -16, 22, 52, 18, 8, 1, 57, 88,
    -- layer=1 filter=58 channel=76
    32, 19, -19, 55, -19, 22, -8, -76, -9,
    -- layer=1 filter=58 channel=77
    24, 12, 11, 10, 31, 31, 18, 16, 8,
    -- layer=1 filter=58 channel=78
    14, -9, -4, -12, -10, 28, 0, -36, -9,
    -- layer=1 filter=58 channel=79
    -63, -22, -29, -54, -40, -9, -48, -11, -70,
    -- layer=1 filter=58 channel=80
    -16, -5, 1, -28, -40, -18, -26, -20, -30,
    -- layer=1 filter=58 channel=81
    11, 40, 33, 31, 49, 43, 21, 39, 24,
    -- layer=1 filter=58 channel=82
    23, 21, 25, 18, 39, 14, 34, 34, 14,
    -- layer=1 filter=58 channel=83
    -7, -37, -44, -38, -48, -58, -51, -66, -50,
    -- layer=1 filter=58 channel=84
    52, 16, -50, 98, -26, -33, -15, -123, -29,
    -- layer=1 filter=58 channel=85
    28, 64, 50, 31, 53, 6, 5, 54, 61,
    -- layer=1 filter=58 channel=86
    -9, -75, -54, -49, -82, -17, -42, -34, 10,
    -- layer=1 filter=58 channel=87
    9, 18, -56, 89, 67, -15, 9, 4, 30,
    -- layer=1 filter=58 channel=88
    30, 42, 25, 35, 22, 22, 12, 22, 18,
    -- layer=1 filter=58 channel=89
    32, 25, 12, 38, 38, 12, 12, 11, 10,
    -- layer=1 filter=58 channel=90
    44, 9, -6, 13, -44, -19, -6, -105, -15,
    -- layer=1 filter=58 channel=91
    -14, -34, -35, -12, -23, -41, -31, -46, -48,
    -- layer=1 filter=58 channel=92
    -8, 19, -19, -17, 1, -7, 7, -26, 32,
    -- layer=1 filter=58 channel=93
    13, 13, 22, 24, 23, 18, 9, 22, 7,
    -- layer=1 filter=58 channel=94
    -8, -55, 13, -27, -39, 15, -94, -68, 21,
    -- layer=1 filter=58 channel=95
    65, 15, -19, 88, -4, -4, 1, -34, 5,
    -- layer=1 filter=58 channel=96
    20, 52, 34, 41, 40, 40, 13, 38, 31,
    -- layer=1 filter=58 channel=97
    3, -27, -10, -15, -22, 0, -25, -17, -13,
    -- layer=1 filter=58 channel=98
    -50, -38, -17, -49, -46, 32, -71, -17, -57,
    -- layer=1 filter=58 channel=99
    2, -26, 36, 0, -19, 41, -15, -16, -13,
    -- layer=1 filter=58 channel=100
    21, -41, -59, 32, -59, -56, -10, -69, -41,
    -- layer=1 filter=58 channel=101
    13, 3, -26, 0, -1, -20, -12, -28, -17,
    -- layer=1 filter=58 channel=102
    -23, -67, -46, -34, -53, -27, -65, -60, -5,
    -- layer=1 filter=58 channel=103
    -17, -33, -68, 37, -24, -59, 32, -38, -34,
    -- layer=1 filter=58 channel=104
    20, 42, -17, 38, 30, -59, 0, 16, 1,
    -- layer=1 filter=58 channel=105
    -23, -19, -6, -32, -25, -5, -20, -4, -2,
    -- layer=1 filter=58 channel=106
    31, -3, -44, 20, -27, -27, -22, -63, -22,
    -- layer=1 filter=58 channel=107
    -2, 15, 3, 8, 16, 5, -4, 17, 8,
    -- layer=1 filter=58 channel=108
    57, 65, -1, 43, 11, 9, 0, -45, 14,
    -- layer=1 filter=58 channel=109
    -7, -4, 9, 0, -5, -9, 3, -6, -7,
    -- layer=1 filter=58 channel=110
    0, 2, -9, -1, -2, -12, -6, -10, -6,
    -- layer=1 filter=58 channel=111
    40, -6, -25, 81, 8, -8, -4, -59, 0,
    -- layer=1 filter=58 channel=112
    6, 4, -38, 36, -25, -19, -44, -45, 24,
    -- layer=1 filter=58 channel=113
    -21, -30, 4, -16, -15, -5, 27, 31, 22,
    -- layer=1 filter=58 channel=114
    -70, -96, -52, -52, -94, -48, -14, -69, -36,
    -- layer=1 filter=58 channel=115
    -38, -77, -2, -108, -41, 8, -84, -16, 10,
    -- layer=1 filter=58 channel=116
    -7, -3, -6, -1, -9, 4, -4, 2, -8,
    -- layer=1 filter=58 channel=117
    -44, -21, -50, 1, -19, -21, -14, -81, -20,
    -- layer=1 filter=58 channel=118
    48, 15, -36, 104, 3, -5, 7, -84, -28,
    -- layer=1 filter=58 channel=119
    81, 72, 0, 64, 11, 26, 11, -55, 11,
    -- layer=1 filter=58 channel=120
    -2, 4, 34, 9, 28, 38, 22, 39, -2,
    -- layer=1 filter=58 channel=121
    5, -14, -17, 29, 9, -2, 26, 11, 32,
    -- layer=1 filter=58 channel=122
    -2, -8, 5, 0, -3, -5, 5, 2, 3,
    -- layer=1 filter=58 channel=123
    16, -10, 1, 39, 29, 5, 19, 8, 10,
    -- layer=1 filter=58 channel=124
    22, 33, 34, 27, 39, 41, 19, 26, 18,
    -- layer=1 filter=58 channel=125
    -28, -60, -47, -36, -46, -38, -2, -40, -37,
    -- layer=1 filter=58 channel=126
    0, -10, 6, -5, -9, 40, -20, 14, -16,
    -- layer=1 filter=58 channel=127
    59, -5, -31, 77, -21, -51, -27, -76, -28,
    -- layer=1 filter=59 channel=0
    -3, -2, -10, 4, 3, -5, 0, -8, -12,
    -- layer=1 filter=59 channel=1
    -4, -6, 3, 0, 7, -4, -10, -8, -10,
    -- layer=1 filter=59 channel=2
    -8, -5, 0, 9, 0, -1, 0, -9, -7,
    -- layer=1 filter=59 channel=3
    -10, -2, 5, 4, -6, -7, -7, 3, 5,
    -- layer=1 filter=59 channel=4
    4, 0, 7, -4, -6, -4, -9, -1, -9,
    -- layer=1 filter=59 channel=5
    -7, -3, -4, -4, -8, -2, 0, 0, 3,
    -- layer=1 filter=59 channel=6
    4, 6, 6, 6, -3, -8, -4, -2, -5,
    -- layer=1 filter=59 channel=7
    -4, -5, -4, 8, -4, 0, -13, -5, 1,
    -- layer=1 filter=59 channel=8
    1, -10, -4, -1, 2, 0, -4, 0, -9,
    -- layer=1 filter=59 channel=9
    -1, 6, -8, -9, 0, -5, 7, -5, -7,
    -- layer=1 filter=59 channel=10
    -1, -5, -1, -3, -10, 0, -9, -2, -9,
    -- layer=1 filter=59 channel=11
    0, 7, -3, 0, 0, -2, -7, 8, -10,
    -- layer=1 filter=59 channel=12
    3, -10, 1, 2, 0, -3, 9, 0, 4,
    -- layer=1 filter=59 channel=13
    -9, -3, 0, 6, -10, -6, -9, -2, -6,
    -- layer=1 filter=59 channel=14
    6, 9, -5, -10, 1, -1, 6, 0, 5,
    -- layer=1 filter=59 channel=15
    -6, -4, 6, 6, 2, 2, -7, 0, 6,
    -- layer=1 filter=59 channel=16
    2, -5, -9, -2, 0, -6, -2, -3, 3,
    -- layer=1 filter=59 channel=17
    -11, 6, 0, 1, -13, 0, -13, -9, 0,
    -- layer=1 filter=59 channel=18
    6, 4, -10, -2, -5, -9, -1, 3, 0,
    -- layer=1 filter=59 channel=19
    -5, -11, 4, -1, 7, 7, -9, 7, 5,
    -- layer=1 filter=59 channel=20
    -13, -3, -6, 5, -3, 0, -3, -4, 0,
    -- layer=1 filter=59 channel=21
    2, 0, -4, 3, -8, 7, 5, -9, -3,
    -- layer=1 filter=59 channel=22
    -2, -7, 5, 0, -1, -2, -2, 9, 0,
    -- layer=1 filter=59 channel=23
    6, 3, -2, 2, 0, -2, 5, 3, -11,
    -- layer=1 filter=59 channel=24
    -4, 4, 2, 4, -13, -5, -5, 0, -1,
    -- layer=1 filter=59 channel=25
    -9, 1, -8, -2, -8, -3, -9, -3, 5,
    -- layer=1 filter=59 channel=26
    3, -10, 5, 0, -13, -5, -9, -7, -15,
    -- layer=1 filter=59 channel=27
    -6, 6, -1, 9, 10, 6, -8, 0, 10,
    -- layer=1 filter=59 channel=28
    2, -8, 0, -5, 4, 5, 3, 1, -9,
    -- layer=1 filter=59 channel=29
    -9, -5, -4, 10, 10, 6, -3, 7, -2,
    -- layer=1 filter=59 channel=30
    0, 0, 0, -6, -15, 2, 8, -3, 0,
    -- layer=1 filter=59 channel=31
    -6, 0, -7, -5, -12, 4, 11, -9, 0,
    -- layer=1 filter=59 channel=32
    -1, -4, 4, -4, 4, 0, 3, 5, -10,
    -- layer=1 filter=59 channel=33
    3, -8, 6, 4, 9, 5, -9, 4, -6,
    -- layer=1 filter=59 channel=34
    1, -9, -7, -9, -9, 5, 5, 0, -3,
    -- layer=1 filter=59 channel=35
    7, -10, -9, -8, 2, 0, -3, 4, 2,
    -- layer=1 filter=59 channel=36
    0, 6, -11, -3, -2, -5, -1, -11, 2,
    -- layer=1 filter=59 channel=37
    4, 2, -8, 2, -2, 0, 1, -2, 1,
    -- layer=1 filter=59 channel=38
    0, 5, 2, 0, -8, -9, 3, -5, 8,
    -- layer=1 filter=59 channel=39
    -3, 5, 0, -7, 3, 3, -2, -3, -7,
    -- layer=1 filter=59 channel=40
    2, -7, -14, -2, -2, 7, 4, 3, 6,
    -- layer=1 filter=59 channel=41
    -4, -8, -1, -12, -8, -1, 3, -2, -5,
    -- layer=1 filter=59 channel=42
    7, -4, -9, 9, 4, -13, 9, -5, -12,
    -- layer=1 filter=59 channel=43
    9, -2, -4, -3, 0, 7, 8, -4, -12,
    -- layer=1 filter=59 channel=44
    0, -13, -1, -5, -9, -7, 2, -13, -8,
    -- layer=1 filter=59 channel=45
    0, 5, -5, 0, 6, -5, 7, -8, -5,
    -- layer=1 filter=59 channel=46
    0, -4, 2, 2, -9, -13, -5, -4, 3,
    -- layer=1 filter=59 channel=47
    1, -5, 0, 6, 7, 2, -3, 2, -7,
    -- layer=1 filter=59 channel=48
    5, 3, 0, -2, -9, -1, 6, 9, -4,
    -- layer=1 filter=59 channel=49
    4, -10, -10, 4, -7, 2, -2, -1, -4,
    -- layer=1 filter=59 channel=50
    5, 8, -13, -2, 6, -5, -9, 3, 0,
    -- layer=1 filter=59 channel=51
    0, -11, -5, -1, -3, 1, 0, 1, -3,
    -- layer=1 filter=59 channel=52
    4, 8, 10, 2, -9, 11, 0, 3, -7,
    -- layer=1 filter=59 channel=53
    -6, -10, 5, -1, 0, -1, -10, -9, -11,
    -- layer=1 filter=59 channel=54
    -2, -7, -9, -1, -4, 0, -9, -7, 7,
    -- layer=1 filter=59 channel=55
    -12, -4, -7, -7, -10, 8, 7, 7, 8,
    -- layer=1 filter=59 channel=56
    -9, 1, 0, 3, 0, -5, 6, -10, 2,
    -- layer=1 filter=59 channel=57
    8, -10, 7, -6, 0, 6, -10, -2, -4,
    -- layer=1 filter=59 channel=58
    -6, -1, 0, -4, -8, -10, -5, 10, -8,
    -- layer=1 filter=59 channel=59
    7, -4, -3, -3, 5, 6, 9, 7, -11,
    -- layer=1 filter=59 channel=60
    0, -6, 5, -8, -2, 11, 10, -7, -8,
    -- layer=1 filter=59 channel=61
    -4, 0, -6, 8, 0, -4, 3, -8, 10,
    -- layer=1 filter=59 channel=62
    1, -4, 4, -4, 3, 1, -4, -3, -1,
    -- layer=1 filter=59 channel=63
    -4, 1, 0, 1, -4, 2, 0, -4, -4,
    -- layer=1 filter=59 channel=64
    -7, 5, -2, -3, -5, -10, 0, -5, 5,
    -- layer=1 filter=59 channel=65
    -8, -12, -10, 2, 3, 3, -3, -11, 0,
    -- layer=1 filter=59 channel=66
    6, 1, -10, 5, -7, -3, -3, -8, -5,
    -- layer=1 filter=59 channel=67
    2, -1, -6, -9, 2, 0, -7, -1, -6,
    -- layer=1 filter=59 channel=68
    2, 9, 4, -12, -11, 2, 3, 4, 0,
    -- layer=1 filter=59 channel=69
    -1, -1, -3, 0, 0, -12, 2, 0, -14,
    -- layer=1 filter=59 channel=70
    -1, 0, -8, -4, -10, 3, 4, 11, 0,
    -- layer=1 filter=59 channel=71
    7, -5, 0, 7, 6, -9, -1, 9, 3,
    -- layer=1 filter=59 channel=72
    -7, -12, 2, 4, -9, 1, -8, 9, -10,
    -- layer=1 filter=59 channel=73
    4, -6, -7, 4, 5, -9, 4, 0, -7,
    -- layer=1 filter=59 channel=74
    5, 0, -7, 0, -5, -7, 6, -11, 3,
    -- layer=1 filter=59 channel=75
    7, -6, -10, 0, -4, 3, -1, 6, 1,
    -- layer=1 filter=59 channel=76
    6, 3, -8, 5, 2, 8, 1, 0, 8,
    -- layer=1 filter=59 channel=77
    -1, -9, -12, -5, 1, 7, 5, -10, 8,
    -- layer=1 filter=59 channel=78
    0, 0, -2, 5, -2, 2, 4, 0, 1,
    -- layer=1 filter=59 channel=79
    -7, 7, 7, 8, -7, 0, -9, -10, 6,
    -- layer=1 filter=59 channel=80
    3, 5, -2, 2, 4, -9, 0, -7, 6,
    -- layer=1 filter=59 channel=81
    0, -9, 4, -5, 4, -6, -6, -13, -2,
    -- layer=1 filter=59 channel=82
    3, -6, 5, -1, -2, -4, 3, -7, -5,
    -- layer=1 filter=59 channel=83
    -5, -12, -10, -5, 0, 4, 9, 4, -7,
    -- layer=1 filter=59 channel=84
    -1, 0, -8, -8, -6, 5, -8, 7, 2,
    -- layer=1 filter=59 channel=85
    -7, 1, 0, 2, 3, 6, -1, -5, -9,
    -- layer=1 filter=59 channel=86
    -11, -9, 8, -4, -4, -10, -9, 0, 0,
    -- layer=1 filter=59 channel=87
    2, -7, 6, 8, -2, 2, -11, 11, -2,
    -- layer=1 filter=59 channel=88
    -14, -7, 4, 1, 0, -7, -7, -10, 6,
    -- layer=1 filter=59 channel=89
    0, -11, -11, -5, -7, -6, 6, -6, -4,
    -- layer=1 filter=59 channel=90
    -8, -8, -6, 7, -11, -5, 3, -11, -11,
    -- layer=1 filter=59 channel=91
    0, -10, 0, 0, -6, 5, -6, 4, -4,
    -- layer=1 filter=59 channel=92
    -8, 5, -4, 1, -4, -8, -5, -10, 6,
    -- layer=1 filter=59 channel=93
    -2, -6, -8, 5, 8, -7, -6, -4, 0,
    -- layer=1 filter=59 channel=94
    6, 7, -2, -3, 5, 6, -10, 1, -12,
    -- layer=1 filter=59 channel=95
    -6, -9, -1, -12, -7, 4, 6, -8, 2,
    -- layer=1 filter=59 channel=96
    -8, -10, 0, 1, 4, -3, 10, -11, 0,
    -- layer=1 filter=59 channel=97
    -7, 0, 6, 5, -9, -1, 2, -2, -11,
    -- layer=1 filter=59 channel=98
    -11, -9, -6, -2, -6, 6, 6, 4, -14,
    -- layer=1 filter=59 channel=99
    5, -2, -11, -1, -3, -11, -2, -9, 6,
    -- layer=1 filter=59 channel=100
    1, 0, -7, -3, -4, -5, 5, 2, -11,
    -- layer=1 filter=59 channel=101
    -1, 4, -3, 0, -7, -8, -9, -2, 0,
    -- layer=1 filter=59 channel=102
    0, -12, -6, -13, -2, 2, -11, 6, 3,
    -- layer=1 filter=59 channel=103
    0, 1, -9, -8, -10, 0, 5, -11, 2,
    -- layer=1 filter=59 channel=104
    -12, 5, -5, 0, -2, -10, -9, 8, -9,
    -- layer=1 filter=59 channel=105
    -9, 4, 1, 0, -5, -5, -4, 1, 0,
    -- layer=1 filter=59 channel=106
    1, 8, -13, -13, -1, -5, 0, 9, -5,
    -- layer=1 filter=59 channel=107
    -8, -8, 5, 0, 7, -3, -5, -7, 9,
    -- layer=1 filter=59 channel=108
    -1, 4, -9, 8, -4, 3, -2, -6, -17,
    -- layer=1 filter=59 channel=109
    6, -8, 2, -8, 5, 6, 2, 7, 7,
    -- layer=1 filter=59 channel=110
    3, -3, -8, -6, -4, -7, 9, -12, -9,
    -- layer=1 filter=59 channel=111
    4, 2, 0, 0, -10, -1, -6, 8, 10,
    -- layer=1 filter=59 channel=112
    0, 3, 5, 1, 1, 2, -6, -6, -6,
    -- layer=1 filter=59 channel=113
    -4, -6, 6, -5, 2, -6, 0, -8, -3,
    -- layer=1 filter=59 channel=114
    4, 3, 12, 4, 7, -1, -5, -10, 0,
    -- layer=1 filter=59 channel=115
    -2, -6, -5, -3, -12, -9, 6, -7, 7,
    -- layer=1 filter=59 channel=116
    -9, -2, -1, -1, 0, -10, 7, 1, 9,
    -- layer=1 filter=59 channel=117
    11, 9, 6, 0, -11, 8, 0, -5, -7,
    -- layer=1 filter=59 channel=118
    -2, -10, -2, -11, -7, -4, -5, -4, 6,
    -- layer=1 filter=59 channel=119
    -2, -3, -2, 1, -5, -12, -13, 0, -5,
    -- layer=1 filter=59 channel=120
    0, -10, -3, 3, 4, -10, 1, -9, 8,
    -- layer=1 filter=59 channel=121
    -3, 5, -13, -1, 2, -7, -8, 1, 0,
    -- layer=1 filter=59 channel=122
    4, -6, -8, 1, -5, 0, 5, 6, -6,
    -- layer=1 filter=59 channel=123
    -7, -9, 1, 2, -6, 1, -3, -10, -7,
    -- layer=1 filter=59 channel=124
    4, -3, 8, -10, 0, 2, 2, -8, -6,
    -- layer=1 filter=59 channel=125
    -11, -2, 8, -10, 3, -10, 5, -4, 2,
    -- layer=1 filter=59 channel=126
    6, 1, 6, 5, 0, 5, -1, 9, -3,
    -- layer=1 filter=59 channel=127
    -4, -4, -3, 6, -10, 8, -8, -5, -8,
    -- layer=1 filter=60 channel=0
    -19, -16, -3, -27, -15, -22, -17, -7, -25,
    -- layer=1 filter=60 channel=1
    10, -8, 16, 28, 6, -8, -2, -7, -4,
    -- layer=1 filter=60 channel=2
    -3, 5, -3, 10, 20, 6, 7, 9, 22,
    -- layer=1 filter=60 channel=3
    -8, -6, 0, 2, -7, 8, -10, -5, 8,
    -- layer=1 filter=60 channel=4
    0, 1, 7, 2, 9, 6, -6, -8, 2,
    -- layer=1 filter=60 channel=5
    2, 1, 5, 27, 7, 12, 9, 12, -19,
    -- layer=1 filter=60 channel=6
    3, 13, 3, -48, 14, -20, -37, -26, -70,
    -- layer=1 filter=60 channel=7
    -3, -2, 17, 12, -35, 13, 17, -27, 42,
    -- layer=1 filter=60 channel=8
    -26, -1, -11, 28, -12, -17, -9, 1, -16,
    -- layer=1 filter=60 channel=9
    -13, -16, -37, 12, 14, 4, 17, -2, -7,
    -- layer=1 filter=60 channel=10
    2, 25, 25, 28, -24, 17, 11, -33, 34,
    -- layer=1 filter=60 channel=11
    -1, -20, -13, -5, -1, -21, 10, -12, 1,
    -- layer=1 filter=60 channel=12
    -34, 24, -1, 5, -6, -24, 7, 20, -6,
    -- layer=1 filter=60 channel=13
    -30, -34, -39, -35, -66, -59, -30, -36, -46,
    -- layer=1 filter=60 channel=14
    -17, 8, 48, 8, -17, 10, -8, 11, 61,
    -- layer=1 filter=60 channel=15
    -21, -59, -4, -5, -17, -57, -59, -55, -29,
    -- layer=1 filter=60 channel=16
    -15, -7, -24, 16, 1, 8, 0, 23, -14,
    -- layer=1 filter=60 channel=17
    -37, -35, -39, -43, -60, -59, -46, -57, -55,
    -- layer=1 filter=60 channel=18
    15, 2, 3, -2, 13, -5, 16, -5, 18,
    -- layer=1 filter=60 channel=19
    -47, -18, 22, 19, 1, 59, 27, 5, -26,
    -- layer=1 filter=60 channel=20
    -40, -28, -14, -58, -73, -68, -66, -56, -52,
    -- layer=1 filter=60 channel=21
    11, 16, 0, 0, 1, -10, -12, -8, -5,
    -- layer=1 filter=60 channel=22
    -65, -61, -21, -31, -61, -96, -42, -49, -29,
    -- layer=1 filter=60 channel=23
    -31, -21, 21, -6, -4, 7, 20, 7, 28,
    -- layer=1 filter=60 channel=24
    23, 39, 3, 42, 33, 42, 40, 29, 29,
    -- layer=1 filter=60 channel=25
    -23, -16, -9, 15, -41, 22, -10, -5, 4,
    -- layer=1 filter=60 channel=26
    -36, -42, -21, -21, -39, -24, -2, 0, 4,
    -- layer=1 filter=60 channel=27
    6, -8, -37, 8, 6, -7, 24, 8, -2,
    -- layer=1 filter=60 channel=28
    -6, 5, 6, 38, -15, 19, 37, -12, 39,
    -- layer=1 filter=60 channel=29
    -12, -20, -31, -17, -27, -27, -20, -36, -41,
    -- layer=1 filter=60 channel=30
    13, 22, 21, 13, 5, 19, 30, 15, 0,
    -- layer=1 filter=60 channel=31
    -24, 8, 2, -15, 0, -13, -21, -25, 1,
    -- layer=1 filter=60 channel=32
    0, -24, 18, 0, -19, 3, 12, 33, 58,
    -- layer=1 filter=60 channel=33
    -10, 3, -3, 0, 8, -8, 8, 9, -5,
    -- layer=1 filter=60 channel=34
    -4, -6, -17, -2, 5, -2, -1, -6, 0,
    -- layer=1 filter=60 channel=35
    1, -5, -2, -7, 1, -4, -15, -3, -8,
    -- layer=1 filter=60 channel=36
    -5, -4, -11, 11, 10, 20, 19, 13, 1,
    -- layer=1 filter=60 channel=37
    16, 28, -27, 18, 8, 16, 24, 22, -27,
    -- layer=1 filter=60 channel=38
    -18, -5, -15, -36, -38, -44, -30, -48, -62,
    -- layer=1 filter=60 channel=39
    -25, -29, -33, -8, -20, -11, -12, -12, -27,
    -- layer=1 filter=60 channel=40
    -48, -2, -31, -43, -32, -25, -23, -43, -16,
    -- layer=1 filter=60 channel=41
    17, -35, 0, 46, -13, 51, 57, 34, 37,
    -- layer=1 filter=60 channel=42
    -26, -12, 5, -10, -1, -5, -11, -3, -10,
    -- layer=1 filter=60 channel=43
    7, -8, -14, 17, -2, 5, 9, 15, 10,
    -- layer=1 filter=60 channel=44
    -12, -33, 0, 12, -8, -10, 0, 13, 34,
    -- layer=1 filter=60 channel=45
    -21, -15, -10, 12, -10, -12, -13, -22, -42,
    -- layer=1 filter=60 channel=46
    -44, -39, 11, -16, -4, 11, -5, -15, -78,
    -- layer=1 filter=60 channel=47
    -27, -16, 24, 7, -6, -20, 9, -8, 0,
    -- layer=1 filter=60 channel=48
    22, -1, -8, -12, -16, -13, -9, -34, -21,
    -- layer=1 filter=60 channel=49
    3, 14, -16, -10, -7, -4, -19, -28, -10,
    -- layer=1 filter=60 channel=50
    -5, -9, -24, 4, 13, 12, -13, -41, 0,
    -- layer=1 filter=60 channel=51
    17, 4, -5, 3, -29, -27, -5, -56, -19,
    -- layer=1 filter=60 channel=52
    -3, -6, 8, 6, 7, 15, 6, 2, 24,
    -- layer=1 filter=60 channel=53
    5, 3, 3, 16, 2, 0, -3, 3, 0,
    -- layer=1 filter=60 channel=54
    14, 23, -15, 35, -17, 37, 25, 3, -10,
    -- layer=1 filter=60 channel=55
    27, -1, -6, 48, 21, 19, 50, 40, 40,
    -- layer=1 filter=60 channel=56
    -1, 3, 7, 5, -8, 8, 0, 7, 0,
    -- layer=1 filter=60 channel=57
    -22, -37, -3, -20, -78, -6, -42, -69, 9,
    -- layer=1 filter=60 channel=58
    -23, -6, 32, 11, -21, 21, 28, -30, 32,
    -- layer=1 filter=60 channel=59
    -9, -7, -18, -6, -11, 0, -23, -24, -26,
    -- layer=1 filter=60 channel=60
    0, -3, -11, 10, 0, 11, -2, -4, -13,
    -- layer=1 filter=60 channel=61
    2, -2, 6, 3, -6, 2, 4, 10, -1,
    -- layer=1 filter=60 channel=62
    -25, -9, -43, 5, 9, 10, 8, 11, -23,
    -- layer=1 filter=60 channel=63
    19, 12, 18, 0, 2, 13, 23, 16, 24,
    -- layer=1 filter=60 channel=64
    -12, -21, 0, -6, -12, -18, -10, -8, -24,
    -- layer=1 filter=60 channel=65
    -1, -5, -1, -5, -10, -22, -25, -11, -33,
    -- layer=1 filter=60 channel=66
    0, -8, 10, 0, 14, 11, 9, -1, -3,
    -- layer=1 filter=60 channel=67
    12, -4, -18, -5, -23, -20, -33, -44, -45,
    -- layer=1 filter=60 channel=68
    -20, -33, -7, 16, 0, 7, 29, 0, 14,
    -- layer=1 filter=60 channel=69
    -25, -9, -24, 19, 23, 6, 14, 31, -13,
    -- layer=1 filter=60 channel=70
    32, 49, -2, -12, 25, 27, -23, -15, -39,
    -- layer=1 filter=60 channel=71
    34, 35, 29, 43, 39, 40, 39, 27, 12,
    -- layer=1 filter=60 channel=72
    -8, 8, 18, 15, 17, -10, 32, -2, -16,
    -- layer=1 filter=60 channel=73
    -1, 12, 0, -1, 9, 13, 13, -1, 8,
    -- layer=1 filter=60 channel=74
    6, 3, -20, -20, 4, 0, 16, -17, -23,
    -- layer=1 filter=60 channel=75
    17, 30, 60, -4, 32, -27, 29, 16, 39,
    -- layer=1 filter=60 channel=76
    21, -11, -5, -9, -14, -27, 6, -3, -15,
    -- layer=1 filter=60 channel=77
    14, 17, -1, 1, 23, 0, -15, -1, -18,
    -- layer=1 filter=60 channel=78
    -28, -17, -16, -13, -23, 2, -31, -23, 0,
    -- layer=1 filter=60 channel=79
    -32, -20, -38, -4, 0, -8, 11, 4, -13,
    -- layer=1 filter=60 channel=80
    -8, 6, 3, 0, -9, -4, -4, 0, 0,
    -- layer=1 filter=60 channel=81
    26, 23, 7, 24, 36, 35, 23, 16, 18,
    -- layer=1 filter=60 channel=82
    19, 17, -3, -7, -1, 4, -12, -18, -8,
    -- layer=1 filter=60 channel=83
    -23, 1, -9, 14, -13, -40, -17, -23, -39,
    -- layer=1 filter=60 channel=84
    15, 2, -10, -28, 3, -19, 29, 13, 39,
    -- layer=1 filter=60 channel=85
    -27, 0, 14, -5, -37, 5, 45, -23, -5,
    -- layer=1 filter=60 channel=86
    -14, -19, -1, -13, -7, -16, -1, -11, -10,
    -- layer=1 filter=60 channel=87
    -53, -13, -9, 1, 24, 28, 17, 18, -19,
    -- layer=1 filter=60 channel=88
    0, 0, -16, -20, -3, -29, -18, -33, -17,
    -- layer=1 filter=60 channel=89
    9, 11, 2, -6, 19, -5, -27, 1, -6,
    -- layer=1 filter=60 channel=90
    -28, -51, -25, -2, -15, -24, 7, -1, -8,
    -- layer=1 filter=60 channel=91
    -15, -27, -33, -36, -50, -39, -40, -77, -37,
    -- layer=1 filter=60 channel=92
    15, -34, -26, 30, -16, -42, 17, -6, 17,
    -- layer=1 filter=60 channel=93
    17, 11, 20, 25, 16, 17, 8, 13, 12,
    -- layer=1 filter=60 channel=94
    -32, -15, -18, -21, -33, -25, -38, -23, -15,
    -- layer=1 filter=60 channel=95
    11, 5, 5, -13, 8, -18, 20, 24, 37,
    -- layer=1 filter=60 channel=96
    12, 1, 8, 10, 10, -7, 19, 1, -1,
    -- layer=1 filter=60 channel=97
    -8, 4, 5, 7, 9, -5, 0, 1, 7,
    -- layer=1 filter=60 channel=98
    -32, -13, -31, 4, -20, -27, 0, -8, -10,
    -- layer=1 filter=60 channel=99
    -14, 21, -9, 27, 33, 31, 40, 26, 18,
    -- layer=1 filter=60 channel=100
    3, -16, -9, -2, -4, -17, 9, -11, -11,
    -- layer=1 filter=60 channel=101
    -20, -14, -21, -45, -28, -39, -43, -46, -35,
    -- layer=1 filter=60 channel=102
    -4, 1, 0, -30, -36, -29, -23, -45, -32,
    -- layer=1 filter=60 channel=103
    9, -7, -7, -11, -13, -19, 8, -2, -5,
    -- layer=1 filter=60 channel=104
    -36, 5, 15, -12, -19, 1, 20, 16, 2,
    -- layer=1 filter=60 channel=105
    1, 0, 2, 6, -5, 2, -4, -11, 9,
    -- layer=1 filter=60 channel=106
    -22, -23, -25, -37, -52, -56, -64, -35, -35,
    -- layer=1 filter=60 channel=107
    -15, -9, -5, 6, 2, -4, 18, 15, 5,
    -- layer=1 filter=60 channel=108
    -9, -52, -29, 28, -3, 2, 18, 17, 46,
    -- layer=1 filter=60 channel=109
    7, -4, -2, -4, 8, -6, 2, -4, 10,
    -- layer=1 filter=60 channel=110
    -8, 5, -9, -12, -2, 2, -9, -10, 0,
    -- layer=1 filter=60 channel=111
    24, 0, 5, -8, 11, -6, 32, 11, 31,
    -- layer=1 filter=60 channel=112
    18, -14, -1, -13, 3, -17, -12, -14, 19,
    -- layer=1 filter=60 channel=113
    -47, -31, -13, -40, -45, -19, -43, -48, -28,
    -- layer=1 filter=60 channel=114
    -27, -28, -42, 26, 20, -1, 24, 21, -27,
    -- layer=1 filter=60 channel=115
    -24, -8, -7, -26, -29, -6, -22, -37, -3,
    -- layer=1 filter=60 channel=116
    8, -3, 4, 1, 0, -8, -9, -8, -13,
    -- layer=1 filter=60 channel=117
    26, -15, 6, -24, 7, -16, 14, 2, 34,
    -- layer=1 filter=60 channel=118
    7, 6, 12, -16, -5, 0, 21, -1, 12,
    -- layer=1 filter=60 channel=119
    -11, -28, -12, 12, -18, 17, 28, 34, 51,
    -- layer=1 filter=60 channel=120
    6, 6, -8, -3, -18, -22, -13, -22, -17,
    -- layer=1 filter=60 channel=121
    2, 19, 8, 44, 27, 36, 34, 49, 31,
    -- layer=1 filter=60 channel=122
    -9, -8, 2, 3, -7, 5, -9, -5, -4,
    -- layer=1 filter=60 channel=123
    21, 28, 24, 41, 26, 45, 46, 40, 46,
    -- layer=1 filter=60 channel=124
    -7, -7, -5, -9, -7, -15, -9, -17, -8,
    -- layer=1 filter=60 channel=125
    43, 68, 20, 1, -1, 32, -20, -21, -44,
    -- layer=1 filter=60 channel=126
    -7, 7, -20, 42, -8, -37, -9, -18, -22,
    -- layer=1 filter=60 channel=127
    20, 14, 14, -14, 5, -7, 8, 5, 9,
    -- layer=1 filter=61 channel=0
    -9, -3, 1, -2, -20, -12, -1, -1, -2,
    -- layer=1 filter=61 channel=1
    0, -20, 3, 9, -1, 3, -1, 0, 7,
    -- layer=1 filter=61 channel=2
    -38, -9, -19, -22, -14, -32, -14, 0, -29,
    -- layer=1 filter=61 channel=3
    -8, -2, 1, -8, -2, 3, -17, 9, -2,
    -- layer=1 filter=61 channel=4
    -3, -9, 0, 4, 6, -5, -1, -2, -6,
    -- layer=1 filter=61 channel=5
    3, -25, 12, 4, 14, -4, -2, -18, 6,
    -- layer=1 filter=61 channel=6
    7, 13, 5, 0, 7, -1, -10, 6, -8,
    -- layer=1 filter=61 channel=7
    2, 53, 24, -17, 61, 39, 11, 28, 57,
    -- layer=1 filter=61 channel=8
    2, -16, 7, 8, -14, -17, 9, -7, 22,
    -- layer=1 filter=61 channel=9
    7, -2, 7, -11, 11, -17, -17, -10, -44,
    -- layer=1 filter=61 channel=10
    -7, 36, 32, -20, 36, 16, -8, 22, 40,
    -- layer=1 filter=61 channel=11
    14, -15, -13, 5, 0, 3, 27, 29, 16,
    -- layer=1 filter=61 channel=12
    -20, -41, -15, -48, -73, -34, -27, -26, 11,
    -- layer=1 filter=61 channel=13
    4, 15, 1, 7, 16, 3, 8, 17, 9,
    -- layer=1 filter=61 channel=14
    -14, 16, -10, -30, -8, 19, -22, -9, 15,
    -- layer=1 filter=61 channel=15
    16, -1, 33, -7, 34, 36, 16, 18, -3,
    -- layer=1 filter=61 channel=16
    -8, -22, 1, 10, -15, -1, 0, -9, -5,
    -- layer=1 filter=61 channel=17
    6, 0, -4, 6, 3, 0, 26, 18, 6,
    -- layer=1 filter=61 channel=18
    -8, -14, 0, -12, -19, 15, 1, -22, -15,
    -- layer=1 filter=61 channel=19
    -18, 15, 11, 0, -3, 40, -8, 11, -12,
    -- layer=1 filter=61 channel=20
    1, 12, 4, 8, 6, 1, 0, 15, 7,
    -- layer=1 filter=61 channel=21
    -3, 3, 5, 3, -21, 2, -14, -4, 5,
    -- layer=1 filter=61 channel=22
    0, 2, 8, -6, 6, -4, 3, 17, 13,
    -- layer=1 filter=61 channel=23
    -3, 58, 22, 34, 54, 88, 28, 47, 29,
    -- layer=1 filter=61 channel=24
    2, 5, 5, 1, -2, -6, 6, 9, -8,
    -- layer=1 filter=61 channel=25
    -24, 21, 19, -34, 14, 9, -7, -9, 29,
    -- layer=1 filter=61 channel=26
    -7, 28, 1, -1, 39, 18, 24, 34, 0,
    -- layer=1 filter=61 channel=27
    -10, -30, -7, -11, -52, -19, -26, -49, -36,
    -- layer=1 filter=61 channel=28
    -18, 2, 13, -24, -3, 0, -34, 0, 25,
    -- layer=1 filter=61 channel=29
    2, 1, 29, -8, -29, 7, -15, -25, 2,
    -- layer=1 filter=61 channel=30
    -26, -9, 6, -32, -31, 8, -12, -34, -34,
    -- layer=1 filter=61 channel=31
    -5, 11, 10, -7, -1, -3, -11, -8, -4,
    -- layer=1 filter=61 channel=32
    14, 38, 29, 17, 48, 27, 15, 42, 31,
    -- layer=1 filter=61 channel=33
    13, 11, 12, -2, 0, -16, 3, -4, 3,
    -- layer=1 filter=61 channel=34
    -9, 10, 26, -12, 1, 5, 8, 5, 5,
    -- layer=1 filter=61 channel=35
    -3, 6, 5, 9, 8, 5, 10, 7, 1,
    -- layer=1 filter=61 channel=36
    0, -21, -14, 18, -17, 3, 7, 7, -5,
    -- layer=1 filter=61 channel=37
    -5, -24, 1, 9, -18, -6, -23, -15, -8,
    -- layer=1 filter=61 channel=38
    10, -5, 10, 9, -2, -5, -7, 5, 6,
    -- layer=1 filter=61 channel=39
    -4, -23, -5, 13, -9, -3, 11, -1, -4,
    -- layer=1 filter=61 channel=40
    0, 8, 14, 0, -7, 11, 1, -17, -4,
    -- layer=1 filter=61 channel=41
    21, 29, 6, -31, 40, -3, -7, 6, -14,
    -- layer=1 filter=61 channel=42
    -34, -7, -24, -40, -39, -23, -15, -20, -18,
    -- layer=1 filter=61 channel=43
    -11, -22, 0, -7, -20, -17, -11, -19, 0,
    -- layer=1 filter=61 channel=44
    24, 30, 20, -8, 37, 8, 29, 31, 38,
    -- layer=1 filter=61 channel=45
    16, 6, -11, 22, 12, -1, 25, 9, 18,
    -- layer=1 filter=61 channel=46
    -42, -11, -23, 0, -16, 25, -36, -29, 6,
    -- layer=1 filter=61 channel=47
    -16, 44, 46, -1, 34, 38, 17, 36, -5,
    -- layer=1 filter=61 channel=48
    -1, -16, 1, -7, -4, 5, 0, -10, -6,
    -- layer=1 filter=61 channel=49
    1, 3, -3, 0, 9, -5, -6, 2, -9,
    -- layer=1 filter=61 channel=50
    10, 14, 4, 6, -20, 0, -7, 13, 0,
    -- layer=1 filter=61 channel=51
    4, 12, 0, -27, -11, 18, -13, -3, 3,
    -- layer=1 filter=61 channel=52
    9, 0, -2, -18, -5, -15, 13, -1, -3,
    -- layer=1 filter=61 channel=53
    -1, 6, 9, -2, 15, 12, -3, 10, 0,
    -- layer=1 filter=61 channel=54
    -16, 22, 22, -30, 0, 3, -7, -8, 31,
    -- layer=1 filter=61 channel=55
    0, 3, 8, 8, 2, 11, 16, 10, 5,
    -- layer=1 filter=61 channel=56
    11, 0, 7, 0, 4, 20, 3, 5, 14,
    -- layer=1 filter=61 channel=57
    -16, 34, 25, -30, 25, 7, -17, 5, 27,
    -- layer=1 filter=61 channel=58
    -4, 91, 43, 36, 64, 68, 25, 82, 51,
    -- layer=1 filter=61 channel=59
    -5, 9, 3, 0, 2, -3, -3, 3, 1,
    -- layer=1 filter=61 channel=60
    2, 5, 17, -2, 16, 17, 7, 10, 21,
    -- layer=1 filter=61 channel=61
    4, -13, -9, -12, -2, -16, 1, -13, 1,
    -- layer=1 filter=61 channel=62
    -12, -5, 16, -10, -3, 6, -10, -12, 3,
    -- layer=1 filter=61 channel=63
    12, -7, -11, 6, -17, -2, 7, 4, 0,
    -- layer=1 filter=61 channel=64
    9, 1, 3, 6, 11, -2, -7, -2, 7,
    -- layer=1 filter=61 channel=65
    4, -8, 2, -3, -22, -10, -17, -15, -5,
    -- layer=1 filter=61 channel=66
    12, 0, -12, 6, -14, 1, 5, -10, -13,
    -- layer=1 filter=61 channel=67
    -10, -14, 9, -32, -28, -14, -16, -27, -2,
    -- layer=1 filter=61 channel=68
    39, 48, 15, 25, 56, 24, 42, 46, 32,
    -- layer=1 filter=61 channel=69
    2, 8, 12, 10, 0, 20, 9, -3, 9,
    -- layer=1 filter=61 channel=70
    -37, -16, 13, -20, 0, -18, -38, -19, -9,
    -- layer=1 filter=61 channel=71
    2, 0, 13, -7, -11, -6, -21, -32, 8,
    -- layer=1 filter=61 channel=72
    -12, -7, -9, -21, -21, 15, -2, -30, -37,
    -- layer=1 filter=61 channel=73
    2, -8, -7, 0, 3, -4, 0, -2, -7,
    -- layer=1 filter=61 channel=74
    4, -1, 0, -9, 10, 0, -14, -2, -1,
    -- layer=1 filter=61 channel=75
    -23, 10, -14, -28, -8, -8, -32, -44, -29,
    -- layer=1 filter=61 channel=76
    17, 4, -13, -1, -10, -27, 18, -2, -7,
    -- layer=1 filter=61 channel=77
    14, -3, -9, -11, -15, 2, 0, -26, 0,
    -- layer=1 filter=61 channel=78
    -20, -9, 11, -26, -6, -7, -15, 2, 11,
    -- layer=1 filter=61 channel=79
    -10, 0, 9, 10, -5, 7, -7, -13, 3,
    -- layer=1 filter=61 channel=80
    0, -13, -3, -3, 0, 3, 8, 16, 6,
    -- layer=1 filter=61 channel=81
    4, -17, -3, 1, -30, -14, 7, -21, -12,
    -- layer=1 filter=61 channel=82
    4, -15, -1, -13, -11, -1, -14, -6, 9,
    -- layer=1 filter=61 channel=83
    4, 2, -14, 5, -6, -7, 28, 5, -2,
    -- layer=1 filter=61 channel=84
    -6, -18, 9, -10, 6, -23, 33, -20, -22,
    -- layer=1 filter=61 channel=85
    -13, 51, 26, 21, 40, 46, 22, 47, -6,
    -- layer=1 filter=61 channel=86
    9, -4, -7, 23, 22, -1, 21, 19, 19,
    -- layer=1 filter=61 channel=87
    23, 11, 0, 0, -2, 23, -17, 11, -31,
    -- layer=1 filter=61 channel=88
    2, 21, 9, 9, 1, 13, 22, 15, 10,
    -- layer=1 filter=61 channel=89
    7, -12, -9, -12, 1, -16, 1, -4, -3,
    -- layer=1 filter=61 channel=90
    35, 48, 27, 13, 45, 19, 33, 46, 24,
    -- layer=1 filter=61 channel=91
    4, 0, 11, -9, 11, 9, -4, 5, -1,
    -- layer=1 filter=61 channel=92
    2, -41, -1, -39, -33, -47, -16, -45, 0,
    -- layer=1 filter=61 channel=93
    -1, -4, 0, -7, -15, -4, -7, -6, -11,
    -- layer=1 filter=61 channel=94
    10, -13, -5, -10, -9, -13, 1, -10, -1,
    -- layer=1 filter=61 channel=95
    -3, -8, -12, -18, -1, -6, 11, -43, -31,
    -- layer=1 filter=61 channel=96
    7, 0, -21, 0, -4, -11, 2, 7, -15,
    -- layer=1 filter=61 channel=97
    2, -3, -2, -5, -1, -19, 6, -6, -11,
    -- layer=1 filter=61 channel=98
    -10, 2, 7, -20, -2, -11, -1, -7, 12,
    -- layer=1 filter=61 channel=99
    11, 33, 51, 10, 41, 59, -4, 43, 70,
    -- layer=1 filter=61 channel=100
    2, -10, -17, -8, -6, 0, 0, 4, 5,
    -- layer=1 filter=61 channel=101
    3, 2, 12, 2, 8, -2, -3, 3, 1,
    -- layer=1 filter=61 channel=102
    6, -11, -9, 3, -21, -10, 2, -14, -20,
    -- layer=1 filter=61 channel=103
    -12, -19, -28, 4, -16, -4, -4, 1, -12,
    -- layer=1 filter=61 channel=104
    -15, 16, 11, 13, 1, 40, 17, 18, -16,
    -- layer=1 filter=61 channel=105
    0, -10, -13, 0, -15, -16, 14, -13, -7,
    -- layer=1 filter=61 channel=106
    13, 8, 0, 8, 29, -4, 18, 24, 11,
    -- layer=1 filter=61 channel=107
    -14, -7, 0, -27, -8, -13, 1, 1, 2,
    -- layer=1 filter=61 channel=108
    24, 37, 31, 8, 49, 18, 17, 44, 26,
    -- layer=1 filter=61 channel=109
    -6, 1, 7, -11, -8, -1, -8, -10, 6,
    -- layer=1 filter=61 channel=110
    -1, 5, 7, -9, -2, -12, 0, 0, -10,
    -- layer=1 filter=61 channel=111
    -26, 0, 8, -9, -14, 11, 11, -27, -35,
    -- layer=1 filter=61 channel=112
    -17, -33, -23, -13, -9, -31, 22, -10, 10,
    -- layer=1 filter=61 channel=113
    -15, -1, 14, -40, -3, 21, -27, 4, -9,
    -- layer=1 filter=61 channel=114
    -8, -22, 3, -8, -25, -6, -14, -19, -15,
    -- layer=1 filter=61 channel=115
    5, 5, -9, 2, 6, -5, 14, 11, 12,
    -- layer=1 filter=61 channel=116
    -8, -1, -7, 3, -10, 4, -3, -2, 3,
    -- layer=1 filter=61 channel=117
    -59, -41, -24, -6, -13, -9, 7, -24, 7,
    -- layer=1 filter=61 channel=118
    3, -7, 3, -6, -1, -16, 7, -20, -37,
    -- layer=1 filter=61 channel=119
    38, 39, 25, 21, 65, 24, 22, 65, 22,
    -- layer=1 filter=61 channel=120
    -4, -9, -7, -8, -4, -2, -9, -6, 18,
    -- layer=1 filter=61 channel=121
    -21, 10, 7, -22, -23, 8, -33, -28, 11,
    -- layer=1 filter=61 channel=122
    7, -7, -9, 8, -7, 0, 7, 4, -7,
    -- layer=1 filter=61 channel=123
    -16, -13, -10, -12, -34, -6, -20, -21, 7,
    -- layer=1 filter=61 channel=124
    10, 4, 22, 6, 10, 1, 6, 4, 7,
    -- layer=1 filter=61 channel=125
    -29, -20, 7, -6, -12, 15, -24, -7, 15,
    -- layer=1 filter=61 channel=126
    -16, -21, 18, -37, -30, -14, 0, -4, 8,
    -- layer=1 filter=61 channel=127
    -16, -9, 3, -12, -10, 2, -3, -44, -19,
    -- layer=1 filter=62 channel=0
    -2, -4, -11, 6, -1, -14, -2, -4, -14,
    -- layer=1 filter=62 channel=1
    11, -6, -3, 6, 19, 6, 4, 1, 8,
    -- layer=1 filter=62 channel=2
    -38, -13, -29, -14, -44, -29, -6, 3, -9,
    -- layer=1 filter=62 channel=3
    -4, 10, 8, -1, 2, 0, 6, -7, 10,
    -- layer=1 filter=62 channel=4
    3, 1, 1, 8, 1, 10, 3, 9, -8,
    -- layer=1 filter=62 channel=5
    26, 6, 20, 11, 11, 27, 19, -11, 16,
    -- layer=1 filter=62 channel=6
    -9, -25, -32, -85, -76, -63, -19, 2, 13,
    -- layer=1 filter=62 channel=7
    -20, -52, 21, -12, -58, 10, -27, -26, 6,
    -- layer=1 filter=62 channel=8
    22, -11, 15, 30, 22, 7, 17, 1, 36,
    -- layer=1 filter=62 channel=9
    -10, -84, 30, 39, -15, -9, -49, -25, 6,
    -- layer=1 filter=62 channel=10
    0, -50, 41, -8, -50, -16, -19, -28, 21,
    -- layer=1 filter=62 channel=11
    11, 1, -9, 21, 25, 4, -7, 6, -4,
    -- layer=1 filter=62 channel=12
    -43, -31, -35, -8, -3, -9, -25, 16, 0,
    -- layer=1 filter=62 channel=13
    4, 7, -2, -6, 2, -4, 14, 31, 12,
    -- layer=1 filter=62 channel=14
    -49, -45, 5, -7, -50, -20, -12, 5, 6,
    -- layer=1 filter=62 channel=15
    -30, -40, -4, -31, -39, -41, -6, -45, -11,
    -- layer=1 filter=62 channel=16
    15, -22, -6, 19, 19, 11, 24, 0, 25,
    -- layer=1 filter=62 channel=17
    5, 4, -15, 8, -4, -15, 0, -4, 11,
    -- layer=1 filter=62 channel=18
    30, 10, 11, 22, 11, -4, -2, 36, -3,
    -- layer=1 filter=62 channel=19
    5, -6, 45, 50, 27, 23, 2, 9, 32,
    -- layer=1 filter=62 channel=20
    -6, 1, -5, -10, -14, -7, 16, -1, 0,
    -- layer=1 filter=62 channel=21
    -32, -25, -23, -29, -11, -24, 1, -14, -12,
    -- layer=1 filter=62 channel=22
    -5, -17, -16, -4, 2, -11, 31, 3, 26,
    -- layer=1 filter=62 channel=23
    -14, 4, 15, -23, -37, 5, 17, -31, 4,
    -- layer=1 filter=62 channel=24
    -11, -16, -2, 0, 6, 15, -7, -21, 4,
    -- layer=1 filter=62 channel=25
    -8, -27, 20, 11, -8, 8, -22, -37, 28,
    -- layer=1 filter=62 channel=26
    -9, -6, 3, -27, 12, -8, 1, 20, -9,
    -- layer=1 filter=62 channel=27
    -39, -21, -51, -10, -18, -25, -25, -20, -20,
    -- layer=1 filter=62 channel=28
    -16, -35, 11, -7, -13, -7, -12, -4, 17,
    -- layer=1 filter=62 channel=29
    -40, -28, -41, -17, -24, -32, -19, -1, -15,
    -- layer=1 filter=62 channel=30
    44, 0, 42, 25, -8, -3, 1, 16, 26,
    -- layer=1 filter=62 channel=31
    -44, -25, -28, -15, -22, -43, -25, -6, -21,
    -- layer=1 filter=62 channel=32
    5, 10, 28, -12, -5, -9, -2, -2, -27,
    -- layer=1 filter=62 channel=33
    7, 7, 0, -6, -7, 0, 6, 5, 4,
    -- layer=1 filter=62 channel=34
    -21, -30, -6, -8, -6, 1, -19, 0, -27,
    -- layer=1 filter=62 channel=35
    -10, -14, -2, -8, -13, -7, -11, -15, -4,
    -- layer=1 filter=62 channel=36
    28, 11, 15, 31, 32, 7, 14, 14, 10,
    -- layer=1 filter=62 channel=37
    26, -3, 8, 7, 28, 12, 12, -9, 20,
    -- layer=1 filter=62 channel=38
    -18, -26, -36, -16, -21, -15, -6, 7, 2,
    -- layer=1 filter=62 channel=39
    -14, -2, -20, -7, 9, -4, -2, 1, 23,
    -- layer=1 filter=62 channel=40
    -20, -30, -42, -12, -56, -41, 9, 22, 12,
    -- layer=1 filter=62 channel=41
    44, -24, 29, -2, 2, -25, -31, -7, -14,
    -- layer=1 filter=62 channel=42
    -23, -18, -35, -5, -23, -49, 3, -22, -31,
    -- layer=1 filter=62 channel=43
    -4, -19, -4, 17, 16, 1, 9, -21, 27,
    -- layer=1 filter=62 channel=44
    -2, -15, 13, -40, 16, 6, -2, 16, -11,
    -- layer=1 filter=62 channel=45
    -21, -34, 8, -24, -3, -3, -22, -19, 4,
    -- layer=1 filter=62 channel=46
    7, 4, 25, 27, 28, 13, 23, -3, 4,
    -- layer=1 filter=62 channel=47
    0, -27, 29, -15, -57, -26, -12, -19, 0,
    -- layer=1 filter=62 channel=48
    -1, -13, -1, 0, -6, -11, -6, 0, 13,
    -- layer=1 filter=62 channel=49
    -10, -17, -28, -14, -31, -26, -22, -2, -12,
    -- layer=1 filter=62 channel=50
    -12, -17, 11, -9, -15, -14, -17, -30, -9,
    -- layer=1 filter=62 channel=51
    -9, -14, 5, -21, -40, -17, -14, -30, -7,
    -- layer=1 filter=62 channel=52
    2, 11, 0, 1, -23, -6, 0, 6, 18,
    -- layer=1 filter=62 channel=53
    -14, 4, 0, -18, -10, -9, -17, -6, -14,
    -- layer=1 filter=62 channel=54
    1, -17, 27, 25, -3, -7, -30, -27, 26,
    -- layer=1 filter=62 channel=55
    17, 7, 0, 5, 12, 19, -1, -3, -5,
    -- layer=1 filter=62 channel=56
    -5, 11, -11, -7, 0, -6, 9, -8, -7,
    -- layer=1 filter=62 channel=57
    -26, -52, 12, -4, -49, -20, -14, -25, 3,
    -- layer=1 filter=62 channel=58
    -31, -46, 36, 1, -107, -14, -24, -57, 14,
    -- layer=1 filter=62 channel=59
    6, -8, 5, -7, -6, 0, 3, -9, 2,
    -- layer=1 filter=62 channel=60
    9, 12, 16, 22, 8, 5, 9, 1, 17,
    -- layer=1 filter=62 channel=61
    0, -4, 0, 4, 6, 10, 5, 10, -5,
    -- layer=1 filter=62 channel=62
    15, -21, 27, 31, 33, 23, 16, 3, 42,
    -- layer=1 filter=62 channel=63
    17, 11, 10, 18, 5, 7, 8, 0, -17,
    -- layer=1 filter=62 channel=64
    3, -8, 3, 0, -14, -20, -12, -13, 4,
    -- layer=1 filter=62 channel=65
    -18, -3, -8, -6, -12, 0, 0, -19, -10,
    -- layer=1 filter=62 channel=66
    1, 7, 5, 4, 4, 1, -9, -8, -1,
    -- layer=1 filter=62 channel=67
    -13, -28, -37, -37, -19, -4, -38, -39, -38,
    -- layer=1 filter=62 channel=68
    12, -12, 15, -41, 4, 14, 9, 6, 11,
    -- layer=1 filter=62 channel=69
    -6, -16, -3, -9, 10, 18, 27, -6, 5,
    -- layer=1 filter=62 channel=70
    5, 20, -36, -33, -9, -38, -45, -35, -37,
    -- layer=1 filter=62 channel=71
    -24, -21, -9, -2, -3, 18, -10, -26, -3,
    -- layer=1 filter=62 channel=72
    2, -10, 28, 9, -1, -19, -22, 8, 13,
    -- layer=1 filter=62 channel=73
    -8, 2, 6, -10, 2, -4, -6, 3, -7,
    -- layer=1 filter=62 channel=74
    4, -3, 0, -9, -24, -17, -2, -1, -1,
    -- layer=1 filter=62 channel=75
    -42, -27, -10, -24, -33, -30, -17, 26, 10,
    -- layer=1 filter=62 channel=76
    18, -9, -1, -15, 9, -12, -6, -7, -8,
    -- layer=1 filter=62 channel=77
    -9, 1, 8, 1, -11, -7, -6, 0, 11,
    -- layer=1 filter=62 channel=78
    4, -2, 11, -14, -4, 5, -10, 7, 7,
    -- layer=1 filter=62 channel=79
    0, -28, 20, 28, 20, 7, 18, -9, 17,
    -- layer=1 filter=62 channel=80
    9, -7, 4, 8, 2, -6, 10, 9, -5,
    -- layer=1 filter=62 channel=81
    -19, -34, -25, -5, -6, 0, -13, -6, 3,
    -- layer=1 filter=62 channel=82
    -13, -10, 4, -5, -9, 5, 1, -10, -9,
    -- layer=1 filter=62 channel=83
    -9, -9, 20, -8, -9, -13, -17, -9, 13,
    -- layer=1 filter=62 channel=84
    42, 13, 2, 17, 19, 0, 13, 41, 13,
    -- layer=1 filter=62 channel=85
    -7, -9, 31, -2, -67, -8, -28, -34, 17,
    -- layer=1 filter=62 channel=86
    13, 6, 7, 4, 17, 6, -8, 3, 2,
    -- layer=1 filter=62 channel=87
    -17, -48, 34, 28, -16, -31, -36, -8, 5,
    -- layer=1 filter=62 channel=88
    -5, 0, -8, -17, -4, -10, 0, 6, 0,
    -- layer=1 filter=62 channel=89
    -21, -4, 9, -28, -31, -15, 10, 10, -23,
    -- layer=1 filter=62 channel=90
    -6, -12, 10, -31, 1, 8, -7, 3, -11,
    -- layer=1 filter=62 channel=91
    11, -12, -9, -25, -21, -35, -1, 3, 4,
    -- layer=1 filter=62 channel=92
    7, -58, -14, -53, -43, -8, -27, -29, -14,
    -- layer=1 filter=62 channel=93
    -4, -2, 0, -8, -5, 3, 1, -16, 7,
    -- layer=1 filter=62 channel=94
    -2, 0, -9, 5, -11, -9, 0, 0, -7,
    -- layer=1 filter=62 channel=95
    23, 2, 26, 4, 7, -6, 16, 40, 3,
    -- layer=1 filter=62 channel=96
    -5, 6, -4, -7, -7, -2, -4, 13, 4,
    -- layer=1 filter=62 channel=97
    -3, -3, 4, 0, 9, -6, 0, 6, 3,
    -- layer=1 filter=62 channel=98
    9, -9, -1, 11, 0, -5, 13, 0, 31,
    -- layer=1 filter=62 channel=99
    -21, -64, -1, -8, -54, -49, -17, 0, 25,
    -- layer=1 filter=62 channel=100
    1, 4, -10, 0, -3, -11, 9, -1, -27,
    -- layer=1 filter=62 channel=101
    8, -1, 2, -15, -17, -30, 15, 0, -4,
    -- layer=1 filter=62 channel=102
    19, 4, 1, -10, -27, -19, -9, 0, 1,
    -- layer=1 filter=62 channel=103
    -6, -1, -11, 3, -3, 1, 0, -12, -24,
    -- layer=1 filter=62 channel=104
    -20, 2, -1, 8, -28, -5, -15, -15, -18,
    -- layer=1 filter=62 channel=105
    10, 6, -2, 11, 8, -9, -11, 3, 1,
    -- layer=1 filter=62 channel=106
    -11, 3, -9, -65, -18, -31, -2, 23, -10,
    -- layer=1 filter=62 channel=107
    11, 6, -6, -2, -4, 3, -13, -6, 3,
    -- layer=1 filter=62 channel=108
    -24, -38, -1, -27, -13, -6, -10, -14, -30,
    -- layer=1 filter=62 channel=109
    -8, 0, -7, 9, 8, 3, -1, -8, -4,
    -- layer=1 filter=62 channel=110
    -5, 7, -3, -5, 5, 4, -6, -9, -9,
    -- layer=1 filter=62 channel=111
    54, 7, 38, 25, 6, 6, 11, 29, 11,
    -- layer=1 filter=62 channel=112
    47, 22, 8, 23, 2, 4, 19, 22, 6,
    -- layer=1 filter=62 channel=113
    -2, 0, -33, 3, -24, -48, 21, -40, -27,
    -- layer=1 filter=62 channel=114
    4, -11, -25, -12, 7, -9, 29, -19, 21,
    -- layer=1 filter=62 channel=115
    3, -3, 15, 18, -4, 12, -1, -5, 25,
    -- layer=1 filter=62 channel=116
    -7, 3, 7, 4, -7, 9, 3, -6, 0,
    -- layer=1 filter=62 channel=117
    67, 14, 31, 35, -16, 18, 31, 40, 40,
    -- layer=1 filter=62 channel=118
    23, 4, 8, 3, -2, 0, 15, 33, 5,
    -- layer=1 filter=62 channel=119
    3, -4, 6, -37, 18, -19, -20, -3, -22,
    -- layer=1 filter=62 channel=120
    -1, -8, -1, -5, -30, -21, -7, -30, 2,
    -- layer=1 filter=62 channel=121
    -19, -22, -4, 10, -1, -9, -4, 9, -11,
    -- layer=1 filter=62 channel=122
    -3, 9, 5, 9, -9, -6, -10, 8, -2,
    -- layer=1 filter=62 channel=123
    -24, -11, -9, 0, -3, 0, 13, 11, 1,
    -- layer=1 filter=62 channel=124
    -7, -6, 0, -6, 2, -5, -10, -11, -1,
    -- layer=1 filter=62 channel=125
    -14, 1, 3, -35, -6, -23, -48, -62, -29,
    -- layer=1 filter=62 channel=126
    15, 23, 30, 21, 5, -13, 30, 9, 50,
    -- layer=1 filter=62 channel=127
    28, 21, 28, 14, 12, -9, 9, 22, 4,
    -- layer=1 filter=63 channel=0
    1, -3, -12, 2, -9, 0, -2, -1, -2,
    -- layer=1 filter=63 channel=1
    6, -9, 0, -3, 6, -5, -3, -3, -10,
    -- layer=1 filter=63 channel=2
    6, 2, -16, -5, -7, 8, -5, 1, 9,
    -- layer=1 filter=63 channel=3
    -6, -4, -5, 6, 0, 8, 5, 10, 0,
    -- layer=1 filter=63 channel=4
    4, -3, -4, 1, -11, 3, -8, 6, 4,
    -- layer=1 filter=63 channel=5
    0, -4, 0, -6, -2, -21, -17, -1, -3,
    -- layer=1 filter=63 channel=6
    -5, -13, -14, 8, 0, 8, -7, -2, -7,
    -- layer=1 filter=63 channel=7
    8, 11, -4, 0, 13, -10, -11, -11, -14,
    -- layer=1 filter=63 channel=8
    1, 2, 3, 3, 5, -15, -15, -4, -4,
    -- layer=1 filter=63 channel=9
    -2, -4, -14, -6, -11, 4, -4, 9, 2,
    -- layer=1 filter=63 channel=10
    7, 0, 1, -9, -13, -13, -3, -4, -19,
    -- layer=1 filter=63 channel=11
    7, -9, -5, -8, 0, 2, 4, 4, -2,
    -- layer=1 filter=63 channel=12
    9, 8, 7, 4, 2, 7, 9, 6, 9,
    -- layer=1 filter=63 channel=13
    -7, 4, -11, 2, -16, -7, -4, 5, 2,
    -- layer=1 filter=63 channel=14
    5, 6, -5, 0, 16, 2, 12, 6, 7,
    -- layer=1 filter=63 channel=15
    5, -12, 1, 7, -12, 7, -8, -3, -7,
    -- layer=1 filter=63 channel=16
    1, -14, 4, 8, -3, -2, -6, 5, 3,
    -- layer=1 filter=63 channel=17
    -6, -6, 3, 3, -3, -4, 5, -3, 6,
    -- layer=1 filter=63 channel=18
    -6, -4, 1, -20, -16, 7, -21, -8, -9,
    -- layer=1 filter=63 channel=19
    0, -1, 4, -6, 5, -11, 3, 7, 2,
    -- layer=1 filter=63 channel=20
    -5, -2, -8, 0, 1, 0, 7, -8, -3,
    -- layer=1 filter=63 channel=21
    -15, -5, 1, -3, 3, -5, -4, -16, 6,
    -- layer=1 filter=63 channel=22
    9, 0, -4, -5, -4, -1, -12, -16, 3,
    -- layer=1 filter=63 channel=23
    -9, -15, 1, -11, 1, 6, -4, -1, -10,
    -- layer=1 filter=63 channel=24
    0, 5, -15, -1, -11, -9, 2, -10, 7,
    -- layer=1 filter=63 channel=25
    -12, -2, 0, -8, 1, -5, -6, -13, 0,
    -- layer=1 filter=63 channel=26
    4, -4, 8, -5, -7, -9, -4, 3, 2,
    -- layer=1 filter=63 channel=27
    0, 4, 2, -13, 1, -5, -7, -25, -1,
    -- layer=1 filter=63 channel=28
    7, -5, 0, 4, 0, -6, -8, 5, -10,
    -- layer=1 filter=63 channel=29
    2, 0, 0, -18, -5, 8, -2, -12, -9,
    -- layer=1 filter=63 channel=30
    -9, 0, 7, -1, 3, 9, -9, -1, 6,
    -- layer=1 filter=63 channel=31
    4, -11, -11, -8, 0, 5, -1, -7, -1,
    -- layer=1 filter=63 channel=32
    3, -1, -9, -9, 6, 0, -4, 14, -1,
    -- layer=1 filter=63 channel=33
    -2, -9, 9, 6, -6, 3, 1, 1, -9,
    -- layer=1 filter=63 channel=34
    -4, -6, 8, -8, -2, -6, 0, 1, 0,
    -- layer=1 filter=63 channel=35
    -1, -9, -3, -2, -10, -3, -12, -9, -11,
    -- layer=1 filter=63 channel=36
    -7, -1, 1, -4, -1, -13, -8, 0, -8,
    -- layer=1 filter=63 channel=37
    -5, -4, 5, 11, -15, -13, -11, -1, -16,
    -- layer=1 filter=63 channel=38
    -11, -2, -2, -7, -2, -7, -11, -11, -6,
    -- layer=1 filter=63 channel=39
    6, 6, -13, -11, -4, -4, -12, -11, -7,
    -- layer=1 filter=63 channel=40
    -6, -5, -17, -6, 2, -4, -1, 5, 8,
    -- layer=1 filter=63 channel=41
    -2, -4, -2, -8, 1, 3, -1, -3, 6,
    -- layer=1 filter=63 channel=42
    -5, 3, -8, 2, 3, -4, -3, 6, 3,
    -- layer=1 filter=63 channel=43
    -3, -13, 1, 3, -6, -1, 2, -15, 0,
    -- layer=1 filter=63 channel=44
    -3, 7, 9, -3, -11, -5, 6, -1, -1,
    -- layer=1 filter=63 channel=45
    -5, -15, 7, -4, -5, 0, -8, 1, -10,
    -- layer=1 filter=63 channel=46
    -21, -12, -12, 4, -4, -11, -6, 1, -2,
    -- layer=1 filter=63 channel=47
    -5, -1, -4, -16, 6, -8, 6, -4, -14,
    -- layer=1 filter=63 channel=48
    -9, -12, 3, 7, 2, 1, -8, -10, -5,
    -- layer=1 filter=63 channel=49
    -5, -2, -18, -14, -10, -12, 6, 1, -1,
    -- layer=1 filter=63 channel=50
    0, -2, 0, 8, -9, -2, -3, -3, -6,
    -- layer=1 filter=63 channel=51
    7, -9, -10, 2, -1, 6, -7, -11, -11,
    -- layer=1 filter=63 channel=52
    1, 6, -2, 0, -9, 5, -2, 2, 4,
    -- layer=1 filter=63 channel=53
    -3, 3, -11, -5, -11, -11, -5, 5, 3,
    -- layer=1 filter=63 channel=54
    -8, -4, 11, 3, -14, -1, -11, -1, 1,
    -- layer=1 filter=63 channel=55
    6, -6, 0, 0, 5, -8, -20, 5, -13,
    -- layer=1 filter=63 channel=56
    3, 7, -7, 7, 6, -3, 8, -1, -3,
    -- layer=1 filter=63 channel=57
    3, 6, -12, -16, -3, -10, -12, 8, 3,
    -- layer=1 filter=63 channel=58
    5, -13, 5, -15, -11, -13, -1, -5, -2,
    -- layer=1 filter=63 channel=59
    -6, -9, 0, -1, 0, 0, 5, 5, 2,
    -- layer=1 filter=63 channel=60
    -2, -3, 8, 3, -1, 8, -8, -8, 6,
    -- layer=1 filter=63 channel=61
    -1, -4, -9, 0, -6, 7, 11, 6, 0,
    -- layer=1 filter=63 channel=62
    -4, -14, -10, 15, -10, -5, -4, -13, -9,
    -- layer=1 filter=63 channel=63
    -8, -13, -5, -3, 1, 6, -5, -5, -1,
    -- layer=1 filter=63 channel=64
    -8, -5, 0, -9, -3, 6, 7, -3, 0,
    -- layer=1 filter=63 channel=65
    5, -10, -4, 0, 4, -9, -1, -12, -9,
    -- layer=1 filter=63 channel=66
    -2, -3, -4, -15, 2, -5, -5, 2, -1,
    -- layer=1 filter=63 channel=67
    0, 7, -3, 7, -1, -2, -2, 8, -7,
    -- layer=1 filter=63 channel=68
    -1, 10, 3, 1, -3, 10, 0, 9, -4,
    -- layer=1 filter=63 channel=69
    -8, -4, -1, 13, -7, -9, -3, 9, 3,
    -- layer=1 filter=63 channel=70
    -15, 2, -13, 0, 13, 4, 7, 2, 6,
    -- layer=1 filter=63 channel=71
    -10, -2, -4, 5, -5, -10, -8, -11, -5,
    -- layer=1 filter=63 channel=72
    -14, -5, -2, -2, -2, 7, -3, 0, 3,
    -- layer=1 filter=63 channel=73
    4, -6, 2, 1, -4, -11, -9, -9, 8,
    -- layer=1 filter=63 channel=74
    -9, 3, -7, 0, -7, -8, 7, 3, -4,
    -- layer=1 filter=63 channel=75
    -5, 0, -1, 4, 11, 17, -9, -6, 6,
    -- layer=1 filter=63 channel=76
    -12, 3, -10, -2, -1, -5, 6, -2, -9,
    -- layer=1 filter=63 channel=77
    2, 0, 7, 5, 6, 1, 1, 0, -9,
    -- layer=1 filter=63 channel=78
    0, -8, -7, 1, -10, -9, 6, 5, -1,
    -- layer=1 filter=63 channel=79
    -6, 7, 5, 7, -15, -2, -16, 4, -5,
    -- layer=1 filter=63 channel=80
    -3, -1, -8, -2, 1, 9, -11, -7, -2,
    -- layer=1 filter=63 channel=81
    -3, 2, 3, 3, -6, -8, -1, -9, -6,
    -- layer=1 filter=63 channel=82
    -9, -18, 4, -12, -5, -9, -8, -7, -10,
    -- layer=1 filter=63 channel=83
    -3, 5, 5, -1, -8, 0, -2, -8, -13,
    -- layer=1 filter=63 channel=84
    -10, 0, 2, 0, -14, -5, -11, -6, 0,
    -- layer=1 filter=63 channel=85
    -2, 9, -6, -4, -10, -5, 4, 12, -14,
    -- layer=1 filter=63 channel=86
    -9, -8, -8, 0, 2, -14, 0, -13, -1,
    -- layer=1 filter=63 channel=87
    -10, 0, -5, 0, -8, -9, -4, -1, -8,
    -- layer=1 filter=63 channel=88
    -13, -6, -16, -2, -4, -7, 0, 0, -6,
    -- layer=1 filter=63 channel=89
    -3, -3, 1, -12, -10, -9, 3, -9, -12,
    -- layer=1 filter=63 channel=90
    6, -1, -2, 1, -4, -4, -3, -2, 5,
    -- layer=1 filter=63 channel=91
    2, 0, 4, 0, 6, -14, -9, 5, 2,
    -- layer=1 filter=63 channel=92
    3, 0, -6, -11, -13, 7, -10, 4, -9,
    -- layer=1 filter=63 channel=93
    -7, -4, -7, 4, -10, -12, -9, 5, -5,
    -- layer=1 filter=63 channel=94
    -8, -11, -1, -5, -4, 4, -2, 0, -6,
    -- layer=1 filter=63 channel=95
    -5, 4, 1, -1, -2, 13, 5, 7, 2,
    -- layer=1 filter=63 channel=96
    -1, -8, -7, 7, 4, -1, 1, 2, -11,
    -- layer=1 filter=63 channel=97
    -7, -11, 1, -1, -7, -7, 1, 0, -6,
    -- layer=1 filter=63 channel=98
    6, -9, 3, -4, -20, -15, -13, 6, -18,
    -- layer=1 filter=63 channel=99
    1, 6, 5, -4, 2, -5, -11, 6, -2,
    -- layer=1 filter=63 channel=100
    -1, -9, 0, -7, -3, 6, -12, -12, -9,
    -- layer=1 filter=63 channel=101
    0, -6, -13, -6, -1, -3, 7, 7, 0,
    -- layer=1 filter=63 channel=102
    5, -7, -12, 3, -3, -1, -7, 1, -10,
    -- layer=1 filter=63 channel=103
    2, -12, 3, -9, -1, -2, -1, -8, -8,
    -- layer=1 filter=63 channel=104
    0, -2, 0, -6, -2, -8, 0, -1, 6,
    -- layer=1 filter=63 channel=105
    -11, 4, 0, -3, -9, -9, -4, 0, -5,
    -- layer=1 filter=63 channel=106
    -2, 6, -3, 4, -7, -1, 4, 9, -13,
    -- layer=1 filter=63 channel=107
    2, 3, 2, 4, -1, -11, -8, -3, -1,
    -- layer=1 filter=63 channel=108
    3, 8, -4, 5, -2, -1, -4, 9, 4,
    -- layer=1 filter=63 channel=109
    -6, -2, 0, -9, 0, -2, 2, 9, 3,
    -- layer=1 filter=63 channel=110
    4, -8, -10, -10, -7, 0, -8, -2, -7,
    -- layer=1 filter=63 channel=111
    -8, -1, -4, -2, -5, 0, 0, 2, -3,
    -- layer=1 filter=63 channel=112
    5, 0, -5, -6, 0, 3, 2, 5, -12,
    -- layer=1 filter=63 channel=113
    -14, 1, -13, -7, 2, 1, -8, 8, -7,
    -- layer=1 filter=63 channel=114
    1, -7, 0, 9, 6, -10, -3, 0, -6,
    -- layer=1 filter=63 channel=115
    -13, -4, -6, -12, -8, 4, -8, -4, 5,
    -- layer=1 filter=63 channel=116
    -4, -9, 1, 10, -2, 2, 7, -8, -2,
    -- layer=1 filter=63 channel=117
    6, 2, 4, 3, -7, -9, -3, -9, 1,
    -- layer=1 filter=63 channel=118
    3, -3, 5, 0, -9, 3, -4, 0, 0,
    -- layer=1 filter=63 channel=119
    -7, -7, 6, -11, 7, 5, -4, 0, -10,
    -- layer=1 filter=63 channel=120
    -8, -11, 0, -6, -14, -15, -1, -9, -18,
    -- layer=1 filter=63 channel=121
    -4, 0, -2, -9, 0, 2, -9, -25, -4,
    -- layer=1 filter=63 channel=122
    -3, 10, 1, 0, 6, -6, -6, -10, -5,
    -- layer=1 filter=63 channel=123
    -17, 3, -15, -18, 0, -1, -2, -13, 1,
    -- layer=1 filter=63 channel=124
    -7, 3, -3, 0, -5, -2, -7, -4, -10,
    -- layer=1 filter=63 channel=125
    1, -7, -11, -5, 8, 4, 0, -7, -6,
    -- layer=1 filter=63 channel=126
    0, 8, 5, 3, 2, 2, -6, 4, -10,
    -- layer=1 filter=63 channel=127
    -15, -3, -4, -1, -9, 5, -14, -2, -3,
    -- layer=1 filter=64 channel=0
    -5, 7, 6, 6, -9, -3, 7, -6, 4,
    -- layer=1 filter=64 channel=1
    -42, -11, -9, -64, -29, -33, 3, -41, -8,
    -- layer=1 filter=64 channel=2
    20, 16, -19, 32, 16, 0, 50, 39, 14,
    -- layer=1 filter=64 channel=3
    -2, 4, -1, -10, -3, 3, 0, 10, 3,
    -- layer=1 filter=64 channel=4
    -5, 10, 7, 1, -4, 7, -5, -12, -5,
    -- layer=1 filter=64 channel=5
    -89, -73, -98, -119, -86, -69, -51, -78, -25,
    -- layer=1 filter=64 channel=6
    -15, -8, 0, 7, -5, -2, -1, 8, -8,
    -- layer=1 filter=64 channel=7
    -24, 40, 21, -6, 29, -1, 37, 38, 29,
    -- layer=1 filter=64 channel=8
    -73, -70, -73, -82, -72, -58, -60, -98, -36,
    -- layer=1 filter=64 channel=9
    -41, 20, -14, -16, -2, -6, 7, -9, 34,
    -- layer=1 filter=64 channel=10
    -25, 28, 7, 11, 37, -5, 40, 37, 17,
    -- layer=1 filter=64 channel=11
    20, 1, 5, 11, -9, -4, 11, 11, 8,
    -- layer=1 filter=64 channel=12
    -32, -46, -12, -77, -88, -1, 13, -11, -20,
    -- layer=1 filter=64 channel=13
    2, 4, -3, -5, 7, 0, 5, 8, 13,
    -- layer=1 filter=64 channel=14
    -7, 28, 34, -33, -7, -10, 10, 23, -5,
    -- layer=1 filter=64 channel=15
    -33, -31, -58, -57, -63, -7, 16, -37, -1,
    -- layer=1 filter=64 channel=16
    -97, -79, -96, -72, -68, -31, -49, -90, -35,
    -- layer=1 filter=64 channel=17
    8, 9, 6, 5, -6, -3, -8, -5, 2,
    -- layer=1 filter=64 channel=18
    0, -4, 19, -30, -8, 8, -24, -31, -12,
    -- layer=1 filter=64 channel=19
    -91, -60, -47, -66, -105, -47, -89, -105, 5,
    -- layer=1 filter=64 channel=20
    0, 9, -14, 14, 13, 4, 20, 7, 8,
    -- layer=1 filter=64 channel=21
    -14, -17, -8, 11, 12, 5, 31, 11, 8,
    -- layer=1 filter=64 channel=22
    -11, 5, -23, -9, 0, -11, 29, 1, 10,
    -- layer=1 filter=64 channel=23
    12, -41, -4, 12, -27, 21, 36, 42, 35,
    -- layer=1 filter=64 channel=24
    -12, 0, 0, -22, 5, 10, 22, -5, 9,
    -- layer=1 filter=64 channel=25
    -47, -2, -19, -2, -7, -22, -7, 32, 24,
    -- layer=1 filter=64 channel=26
    -7, 2, -1, -3, 15, -1, 26, 37, 26,
    -- layer=1 filter=64 channel=27
    13, -14, -1, 11, 0, -12, -1, -11, -16,
    -- layer=1 filter=64 channel=28
    -34, 20, 15, 2, 30, 1, 23, 33, 4,
    -- layer=1 filter=64 channel=29
    -7, -25, -37, -13, -25, -25, -36, -46, -46,
    -- layer=1 filter=64 channel=30
    -21, -3, 0, -26, -45, -15, -63, -65, -12,
    -- layer=1 filter=64 channel=31
    6, 13, 34, 18, -2, 15, 4, 17, 34,
    -- layer=1 filter=64 channel=32
    -12, 2, 17, 5, 7, 12, 19, 45, 24,
    -- layer=1 filter=64 channel=33
    -20, -20, -15, 4, 1, -8, 3, 15, 25,
    -- layer=1 filter=64 channel=34
    -46, -44, -30, -45, -37, -16, -36, -41, -26,
    -- layer=1 filter=64 channel=35
    -3, -19, -4, -16, -4, -19, -8, -13, -3,
    -- layer=1 filter=64 channel=36
    11, 15, 17, 21, 5, -4, 11, 10, -4,
    -- layer=1 filter=64 channel=37
    -141, -103, -102, -107, -112, -44, -53, -95, -30,
    -- layer=1 filter=64 channel=38
    3, 10, -6, 18, 12, 3, 20, 18, 1,
    -- layer=1 filter=64 channel=39
    -2, -3, -1, 2, -9, -2, -7, -2, -14,
    -- layer=1 filter=64 channel=40
    20, 27, 17, 23, 19, 31, 19, 20, 23,
    -- layer=1 filter=64 channel=41
    3, -31, 11, -9, -10, 13, 0, 24, 9,
    -- layer=1 filter=64 channel=42
    44, 16, 13, 48, 26, 17, 76, 57, 7,
    -- layer=1 filter=64 channel=43
    -68, -57, -73, -50, -57, -30, -17, -62, -24,
    -- layer=1 filter=64 channel=44
    16, 30, 4, 10, 20, 1, 47, 58, 24,
    -- layer=1 filter=64 channel=45
    -24, 6, -9, -19, -8, 3, 24, -6, -4,
    -- layer=1 filter=64 channel=46
    -42, -35, -27, -40, -80, -10, -20, -38, 19,
    -- layer=1 filter=64 channel=47
    13, -16, -19, 17, -17, 38, 68, 54, 53,
    -- layer=1 filter=64 channel=48
    -1, -8, -2, 11, 3, 15, 12, -5, -4,
    -- layer=1 filter=64 channel=49
    10, 5, -1, 14, 14, 28, 40, 20, 29,
    -- layer=1 filter=64 channel=50
    5, 10, 14, 13, 20, 16, -2, 7, 25,
    -- layer=1 filter=64 channel=51
    6, 15, -10, 5, 17, -5, 26, 18, 16,
    -- layer=1 filter=64 channel=52
    9, 15, -5, 1, -4, -6, -7, -9, 0,
    -- layer=1 filter=64 channel=53
    -3, -12, -1, -4, -21, 1, -16, 1, -21,
    -- layer=1 filter=64 channel=54
    -45, -27, -29, -1, -35, -18, -13, 1, 5,
    -- layer=1 filter=64 channel=55
    4, -6, -3, -2, -4, -5, 1, 2, -12,
    -- layer=1 filter=64 channel=56
    3, 9, 0, 8, 5, 2, 1, -3, 0,
    -- layer=1 filter=64 channel=57
    -11, 32, 4, 10, 36, 0, 24, 40, 26,
    -- layer=1 filter=64 channel=58
    -4, -20, -12, 35, 14, 34, 66, 63, 53,
    -- layer=1 filter=64 channel=59
    6, -13, 5, 13, -3, 4, -7, -5, -2,
    -- layer=1 filter=64 channel=60
    3, 16, 4, -4, 3, -2, 13, -2, 17,
    -- layer=1 filter=64 channel=61
    1, 2, -3, -10, 0, -1, 11, 1, 0,
    -- layer=1 filter=64 channel=62
    -115, -102, -91, -83, -98, -35, -77, -95, -28,
    -- layer=1 filter=64 channel=63
    8, -4, 4, -2, 0, -2, -11, -14, -7,
    -- layer=1 filter=64 channel=64
    -7, 6, -14, -26, 0, 0, 0, -7, -9,
    -- layer=1 filter=64 channel=65
    1, 10, -3, 16, 1, -15, 19, 5, 4,
    -- layer=1 filter=64 channel=66
    -4, -15, -3, -14, -5, -9, 3, -16, -4,
    -- layer=1 filter=64 channel=67
    2, 0, 5, 2, -18, -2, 12, -21, -21,
    -- layer=1 filter=64 channel=68
    0, 19, 20, -7, 27, -9, 39, 59, 16,
    -- layer=1 filter=64 channel=69
    -39, -3, -32, -41, -18, -15, 7, -21, -8,
    -- layer=1 filter=64 channel=70
    -41, -49, -14, -30, -60, -33, -41, -71, -34,
    -- layer=1 filter=64 channel=71
    -15, -21, 0, -3, -5, 9, 3, -15, -6,
    -- layer=1 filter=64 channel=72
    -7, 25, 31, -53, -61, -19, -43, -47, 8,
    -- layer=1 filter=64 channel=73
    4, -4, 4, 4, -9, -7, 1, -4, -2,
    -- layer=1 filter=64 channel=74
    -11, 13, -1, -8, 24, -18, 14, 54, 10,
    -- layer=1 filter=64 channel=75
    -4, -14, 14, -26, -38, 7, -76, -4, -40,
    -- layer=1 filter=64 channel=76
    15, 6, 11, 0, -2, -8, -5, 11, -6,
    -- layer=1 filter=64 channel=77
    4, 3, 6, 12, 7, -2, 22, -6, 4,
    -- layer=1 filter=64 channel=78
    -6, 10, -11, 8, 2, -7, -3, -2, 6,
    -- layer=1 filter=64 channel=79
    -82, -74, -73, -63, -71, -24, -41, -72, -19,
    -- layer=1 filter=64 channel=80
    -7, -10, -7, -3, 3, 10, -5, -1, 5,
    -- layer=1 filter=64 channel=81
    -11, -14, 8, -13, -3, 16, 16, -18, -4,
    -- layer=1 filter=64 channel=82
    1, -10, 11, 0, 1, -3, 7, 12, 14,
    -- layer=1 filter=64 channel=83
    -9, 2, -31, -25, -25, -32, -2, -25, -16,
    -- layer=1 filter=64 channel=84
    3, -9, 17, -20, -12, 13, -16, -15, -6,
    -- layer=1 filter=64 channel=85
    6, -33, -6, 28, -31, 25, 52, 32, 30,
    -- layer=1 filter=64 channel=86
    24, 11, 13, 5, 4, 8, 1, 1, 10,
    -- layer=1 filter=64 channel=87
    -22, 12, -7, -50, -16, -14, 2, -23, 20,
    -- layer=1 filter=64 channel=88
    2, -10, 9, 12, -4, 0, 19, 0, -1,
    -- layer=1 filter=64 channel=89
    4, 7, -1, 11, 6, 19, 17, 17, -3,
    -- layer=1 filter=64 channel=90
    -4, 25, 17, -10, 19, -5, 38, 39, 19,
    -- layer=1 filter=64 channel=91
    19, 12, 8, 13, 4, 11, 18, 12, 10,
    -- layer=1 filter=64 channel=92
    -16, 0, -26, -19, -20, -30, 58, -12, -14,
    -- layer=1 filter=64 channel=93
    -9, 5, -1, 9, -9, -4, 14, -8, -14,
    -- layer=1 filter=64 channel=94
    3, 26, -3, 0, 6, -5, 4, 4, 8,
    -- layer=1 filter=64 channel=95
    -22, -15, -8, -41, -18, -8, -55, -33, -37,
    -- layer=1 filter=64 channel=96
    -9, -10, -6, -1, 6, 11, -5, -6, -1,
    -- layer=1 filter=64 channel=97
    -4, 15, 8, -9, -9, -11, -3, -9, -17,
    -- layer=1 filter=64 channel=98
    -61, -34, -50, -26, -44, -39, -21, -50, -24,
    -- layer=1 filter=64 channel=99
    -11, 39, 3, 36, 47, -22, 33, 50, 32,
    -- layer=1 filter=64 channel=100
    -4, -5, 0, -12, -17, -15, -6, -13, -1,
    -- layer=1 filter=64 channel=101
    6, 19, 12, 0, 7, -3, 5, 19, 12,
    -- layer=1 filter=64 channel=102
    18, 19, 6, 9, 0, -2, 6, 2, 0,
    -- layer=1 filter=64 channel=103
    -6, -8, 17, -9, -10, -2, 0, 5, 1,
    -- layer=1 filter=64 channel=104
    3, -14, -2, 3, -17, 29, 13, 26, 22,
    -- layer=1 filter=64 channel=105
    5, 6, 9, 0, 8, -8, -10, -17, -15,
    -- layer=1 filter=64 channel=106
    15, -3, 18, -4, 18, 11, 20, 15, 6,
    -- layer=1 filter=64 channel=107
    0, 6, 10, 3, -21, -11, 0, 3, 1,
    -- layer=1 filter=64 channel=108
    -9, -14, -12, -6, 0, 11, 35, 39, 0,
    -- layer=1 filter=64 channel=109
    8, 10, 0, -4, 6, 6, -4, 4, -3,
    -- layer=1 filter=64 channel=110
    0, 5, -8, 4, -9, -10, -3, -2, 0,
    -- layer=1 filter=64 channel=111
    -21, -22, -1, -53, -19, 3, -69, -72, -36,
    -- layer=1 filter=64 channel=112
    -58, -27, -23, -46, -36, 4, -51, -68, -58,
    -- layer=1 filter=64 channel=113
    -16, -21, -20, 2, -11, -6, 9, -5, -5,
    -- layer=1 filter=64 channel=114
    -23, -40, -53, -48, -96, -47, -51, -83, -18,
    -- layer=1 filter=64 channel=115
    5, 24, 18, 19, 12, 17, 9, 15, 8,
    -- layer=1 filter=64 channel=116
    3, -3, 2, 0, -11, 10, -10, 6, 7,
    -- layer=1 filter=64 channel=117
    -98, -44, -31, -97, -76, -32, -101, -115, -65,
    -- layer=1 filter=64 channel=118
    13, -5, 26, -9, 18, 18, -20, 4, 14,
    -- layer=1 filter=64 channel=119
    -11, 13, 16, -21, 10, -1, 28, 41, 17,
    -- layer=1 filter=64 channel=120
    -21, 2, -16, 9, 0, 4, 23, 0, 14,
    -- layer=1 filter=64 channel=121
    10, -3, 3, -1, -20, -6, -27, -29, -11,
    -- layer=1 filter=64 channel=122
    8, -2, 10, -2, -8, -2, 9, 10, 4,
    -- layer=1 filter=64 channel=123
    13, -12, 5, -15, -8, -20, -17, -19, -24,
    -- layer=1 filter=64 channel=124
    -5, -9, -13, -17, -13, -7, -3, -18, -12,
    -- layer=1 filter=64 channel=125
    -31, -29, -9, -28, -34, -39, -19, -25, -24,
    -- layer=1 filter=64 channel=126
    -63, -18, -36, -88, -57, -70, -92, -118, -53,
    -- layer=1 filter=64 channel=127
    -3, -10, 29, -12, 2, 3, -41, -18, -10,
    -- layer=1 filter=65 channel=0
    34, 8, -9, 26, -5, -5, 4, -7, -2,
    -- layer=1 filter=65 channel=1
    -7, 5, -12, -41, -40, -4, -10, 6, 16,
    -- layer=1 filter=65 channel=2
    -4, 16, 26, -21, -9, 12, -54, -54, -4,
    -- layer=1 filter=65 channel=3
    -2, 0, -1, 4, -10, 4, -6, 13, 10,
    -- layer=1 filter=65 channel=4
    7, 8, 6, 0, 9, -4, -3, -1, 13,
    -- layer=1 filter=65 channel=5
    -10, -1, 0, -78, -72, 11, -1, -8, 7,
    -- layer=1 filter=65 channel=6
    -35, -3, 18, -8, 25, 57, 34, 48, 63,
    -- layer=1 filter=65 channel=7
    24, -54, -64, 21, -49, -85, 1, -14, -74,
    -- layer=1 filter=65 channel=8
    2, 18, 14, -37, -11, -4, 0, 1, 4,
    -- layer=1 filter=65 channel=9
    -22, 18, 16, -35, -9, 16, -11, -13, 7,
    -- layer=1 filter=65 channel=10
    19, -80, -75, 0, -41, -105, 11, -10, -84,
    -- layer=1 filter=65 channel=11
    19, 12, -1, 12, 1, -23, 5, 2, 13,
    -- layer=1 filter=65 channel=12
    9, 10, 15, 18, -6, -25, -52, 5, -1,
    -- layer=1 filter=65 channel=13
    -22, 3, 18, -16, 23, 24, -1, 12, 19,
    -- layer=1 filter=65 channel=14
    10, -19, -39, 0, -57, -42, -51, 17, -63,
    -- layer=1 filter=65 channel=15
    -45, 18, -42, -13, -31, 19, -59, 28, 52,
    -- layer=1 filter=65 channel=16
    -3, -11, 3, -62, -58, -13, 3, -14, -14,
    -- layer=1 filter=65 channel=17
    47, 19, 2, 4, 22, 0, -6, -15, -25,
    -- layer=1 filter=65 channel=18
    35, 16, 1, 6, -7, -19, 8, -14, 11,
    -- layer=1 filter=65 channel=19
    -17, -6, 1, -45, -2, -24, 54, -20, -5,
    -- layer=1 filter=65 channel=20
    2, -1, 0, -11, 14, 10, -5, 9, 13,
    -- layer=1 filter=65 channel=21
    -41, -26, -7, -1, 0, -16, 3, 21, 9,
    -- layer=1 filter=65 channel=22
    -28, -6, -2, -33, 5, 16, -1, 13, 20,
    -- layer=1 filter=65 channel=23
    -20, -10, -47, 17, -20, -49, 16, -16, -44,
    -- layer=1 filter=65 channel=24
    -40, -14, 0, -35, 0, -24, -31, -10, -5,
    -- layer=1 filter=65 channel=25
    13, -64, -26, 6, -56, -69, 30, -38, -96,
    -- layer=1 filter=65 channel=26
    -21, 49, 24, 5, 27, 15, -18, 1, 20,
    -- layer=1 filter=65 channel=27
    38, 32, 20, 22, 18, 20, 7, 19, 47,
    -- layer=1 filter=65 channel=28
    6, -40, -60, 20, -20, -61, -4, 1, -59,
    -- layer=1 filter=65 channel=29
    8, 2, 0, 6, -5, 3, -10, -19, 2,
    -- layer=1 filter=65 channel=30
    48, 17, 5, -4, -3, -20, 31, -9, 6,
    -- layer=1 filter=65 channel=31
    -4, -52, -27, -32, -34, -24, -19, 2, 18,
    -- layer=1 filter=65 channel=32
    -1, 48, 18, 28, 26, 32, -2, 22, 33,
    -- layer=1 filter=65 channel=33
    9, 9, 16, 13, 36, 12, 31, 37, 11,
    -- layer=1 filter=65 channel=34
    -17, -13, 22, -5, 13, 30, 17, 28, 33,
    -- layer=1 filter=65 channel=35
    0, -7, -7, -13, -21, 3, -21, -3, -14,
    -- layer=1 filter=65 channel=36
    47, 17, 14, 24, 15, -7, 29, 15, 11,
    -- layer=1 filter=65 channel=37
    -2, -23, 2, -73, -55, 1, 13, -7, -10,
    -- layer=1 filter=65 channel=38
    -25, -5, 2, 4, 27, 14, 12, 30, 11,
    -- layer=1 filter=65 channel=39
    13, -2, -15, -5, 5, -16, -18, -3, -10,
    -- layer=1 filter=65 channel=40
    -6, -15, 14, 2, -6, 14, 0, 20, 26,
    -- layer=1 filter=65 channel=41
    53, 37, 9, 12, -15, 0, 22, -27, -5,
    -- layer=1 filter=65 channel=42
    12, -10, 19, 21, -6, -6, -101, -99, -27,
    -- layer=1 filter=65 channel=43
    0, 0, -19, -20, -55, -29, 7, -15, -22,
    -- layer=1 filter=65 channel=44
    -3, 67, 35, 39, 53, 18, 11, 28, 38,
    -- layer=1 filter=65 channel=45
    -29, -2, 0, -9, 9, 1, -19, 20, 33,
    -- layer=1 filter=65 channel=46
    -47, -81, -41, -42, -40, -16, 16, 2, 10,
    -- layer=1 filter=65 channel=47
    -45, -32, -41, -37, -38, 1, -31, -1, 35,
    -- layer=1 filter=65 channel=48
    0, -9, 8, 11, 7, 10, 3, 0, -1,
    -- layer=1 filter=65 channel=49
    -32, -29, -19, -22, -10, 28, 4, 16, 41,
    -- layer=1 filter=65 channel=50
    -5, 2, 28, 11, 3, 25, 21, 29, 3,
    -- layer=1 filter=65 channel=51
    3, -22, -20, 13, 15, 7, 9, 13, 12,
    -- layer=1 filter=65 channel=52
    10, 3, 1, -1, 0, 3, 0, 2, -1,
    -- layer=1 filter=65 channel=53
    -16, 1, -12, -12, -4, -10, -7, -5, 1,
    -- layer=1 filter=65 channel=54
    21, -67, 10, -28, -66, -68, 19, -71, -83,
    -- layer=1 filter=65 channel=55
    6, 0, -6, 11, -2, -6, 21, -10, -2,
    -- layer=1 filter=65 channel=56
    -9, 3, 6, 4, -10, 5, 11, 2, 1,
    -- layer=1 filter=65 channel=57
    7, -76, -46, -15, -16, -43, 10, 1, -31,
    -- layer=1 filter=65 channel=58
    -7, -112, -82, 12, -103, -105, 57, -44, -97,
    -- layer=1 filter=65 channel=59
    -5, 3, -13, -1, -7, -10, -1, -8, -8,
    -- layer=1 filter=65 channel=60
    17, 5, 12, 4, 3, 6, 20, 8, 23,
    -- layer=1 filter=65 channel=61
    -9, -12, -4, -1, 9, 0, 0, -9, -11,
    -- layer=1 filter=65 channel=62
    -2, 1, 14, -77, -29, -16, -15, -13, -27,
    -- layer=1 filter=65 channel=63
    32, 20, 2, 16, -9, -10, 18, 4, 7,
    -- layer=1 filter=65 channel=64
    -1, 3, 3, -10, -9, 6, 0, 0, -1,
    -- layer=1 filter=65 channel=65
    -5, -2, 5, -1, -4, -2, 15, 14, -6,
    -- layer=1 filter=65 channel=66
    22, 13, -5, 8, -10, -12, 9, -5, -7,
    -- layer=1 filter=65 channel=67
    -39, -31, -34, -37, -8, 0, -5, 11, 6,
    -- layer=1 filter=65 channel=68
    28, 69, 21, 48, 45, 30, 15, 19, 40,
    -- layer=1 filter=65 channel=69
    -30, 13, -25, -21, -11, -14, -52, 18, 10,
    -- layer=1 filter=65 channel=70
    -57, -60, -43, -44, -39, -8, -3, 11, 20,
    -- layer=1 filter=65 channel=71
    -31, -24, -39, -7, -33, -40, -5, -3, -26,
    -- layer=1 filter=65 channel=72
    18, 19, 11, -9, -3, -10, 36, -2, 15,
    -- layer=1 filter=65 channel=73
    1, 3, -2, -8, -13, -5, -10, -14, -3,
    -- layer=1 filter=65 channel=74
    32, 59, 29, 16, 6, -5, 33, 13, 0,
    -- layer=1 filter=65 channel=75
    29, -29, -4, -16, -49, -53, -21, -33, 4,
    -- layer=1 filter=65 channel=76
    21, 34, 5, 15, 25, 9, -2, -10, 0,
    -- layer=1 filter=65 channel=77
    -7, -25, -12, -8, -11, -16, 0, 1, 0,
    -- layer=1 filter=65 channel=78
    24, 0, -8, -13, -10, -18, -6, 15, -21,
    -- layer=1 filter=65 channel=79
    -8, -10, 11, -59, -32, -7, 5, 9, 2,
    -- layer=1 filter=65 channel=80
    2, 4, 7, 1, -13, -2, 1, 2, -3,
    -- layer=1 filter=65 channel=81
    -12, -16, -21, -11, -14, -8, -12, -10, -30,
    -- layer=1 filter=65 channel=82
    -35, -14, -9, -15, -3, 3, 0, 9, 11,
    -- layer=1 filter=65 channel=83
    -24, 19, -24, -5, 5, 16, -32, 5, 21,
    -- layer=1 filter=65 channel=84
    43, 64, 51, 24, 23, 27, 22, -8, 6,
    -- layer=1 filter=65 channel=85
    -9, -55, -34, 11, -61, -44, 37, -36, -63,
    -- layer=1 filter=65 channel=86
    29, 3, -16, 12, -24, -23, -7, -2, -12,
    -- layer=1 filter=65 channel=87
    13, -3, 19, -39, 21, -2, 33, -10, 15,
    -- layer=1 filter=65 channel=88
    -8, -12, -3, 2, 0, -2, -2, 19, 8,
    -- layer=1 filter=65 channel=89
    -29, -7, -3, 2, 8, 20, 12, 24, 11,
    -- layer=1 filter=65 channel=90
    2, 60, 14, 22, 32, 19, -6, 33, 34,
    -- layer=1 filter=65 channel=91
    -10, -13, 3, -7, -4, 6, 4, 4, 12,
    -- layer=1 filter=65 channel=92
    -20, 9, -41, 7, -40, 21, -52, 2, 15,
    -- layer=1 filter=65 channel=93
    -5, 1, -10, 2, -4, -15, 4, 1, -10,
    -- layer=1 filter=65 channel=94
    27, 6, -2, 30, 13, -4, -1, -7, -25,
    -- layer=1 filter=65 channel=95
    30, 51, 27, 34, 23, 27, 28, 5, 13,
    -- layer=1 filter=65 channel=96
    18, 1, 7, 0, -7, 12, 12, 0, 5,
    -- layer=1 filter=65 channel=97
    14, 14, -12, 9, 9, -7, -5, -4, -21,
    -- layer=1 filter=65 channel=98
    13, -4, 2, -34, -2, -6, 17, 8, -8,
    -- layer=1 filter=65 channel=99
    -9, -31, -74, -11, 8, -74, -14, 18, -46,
    -- layer=1 filter=65 channel=100
    29, 16, 4, 17, 10, -9, 11, 9, 29,
    -- layer=1 filter=65 channel=101
    -14, 10, -3, 3, 15, 16, 0, 24, 1,
    -- layer=1 filter=65 channel=102
    33, 16, 3, 32, 5, -2, 7, 1, -16,
    -- layer=1 filter=65 channel=103
    23, 13, 15, 0, 20, 0, 0, -2, 24,
    -- layer=1 filter=65 channel=104
    -14, -2, -27, 4, 8, -10, 28, 13, -14,
    -- layer=1 filter=65 channel=105
    26, 3, -1, 18, 9, -15, -10, -7, -21,
    -- layer=1 filter=65 channel=106
    -18, 28, 23, -1, 18, 26, -6, 24, 30,
    -- layer=1 filter=65 channel=107
    7, 17, 13, 3, 1, -5, 7, 15, 0,
    -- layer=1 filter=65 channel=108
    -4, 63, 20, 32, 46, 15, -16, 32, 26,
    -- layer=1 filter=65 channel=109
    -6, -5, 3, -1, -1, 6, 0, 1, 8,
    -- layer=1 filter=65 channel=110
    7, 11, -2, 4, -2, 1, 1, -2, -14,
    -- layer=1 filter=65 channel=111
    52, 24, 21, 5, 0, 0, 19, -3, -3,
    -- layer=1 filter=65 channel=112
    3, 27, 16, 21, -14, 7, -24, -16, -23,
    -- layer=1 filter=65 channel=113
    -41, -31, -1, -23, -21, 34, 2, -4, 31,
    -- layer=1 filter=65 channel=114
    0, 10, -18, -3, -28, 22, -25, -17, 0,
    -- layer=1 filter=65 channel=115
    23, -14, -34, 14, -26, -39, -4, -8, -45,
    -- layer=1 filter=65 channel=116
    -1, 3, -10, -6, 1, 0, 0, -4, 3,
    -- layer=1 filter=65 channel=117
    -1, -39, 4, -28, -35, -13, -72, -35, -22,
    -- layer=1 filter=65 channel=118
    39, 48, 20, -4, 27, 17, 16, 12, 29,
    -- layer=1 filter=65 channel=119
    3, 48, 29, 10, 43, 16, 9, 19, 36,
    -- layer=1 filter=65 channel=120
    -11, -47, 12, -10, -7, -3, 6, -2, -11,
    -- layer=1 filter=65 channel=121
    7, -31, -32, -30, -30, -39, -6, -4, 18,
    -- layer=1 filter=65 channel=122
    3, 4, -6, 7, 9, -1, 7, 4, 5,
    -- layer=1 filter=65 channel=123
    25, 7, -9, 3, -11, -14, 17, 8, 7,
    -- layer=1 filter=65 channel=124
    3, -17, -20, -2, -4, -10, -17, -15, -6,
    -- layer=1 filter=65 channel=125
    -62, -61, -29, -60, -52, 8, -9, 12, 39,
    -- layer=1 filter=65 channel=126
    10, -18, -28, -74, 0, -14, -49, -11, 4,
    -- layer=1 filter=65 channel=127
    27, 37, 31, 25, 15, -3, 4, 2, 25,
    -- layer=1 filter=66 channel=0
    -3, 3, -1, -11, 2, -5, 7, -10, -10,
    -- layer=1 filter=66 channel=1
    -13, -15, -3, -3, -21, -15, -6, -15, -5,
    -- layer=1 filter=66 channel=2
    0, 3, 1, -8, -2, -13, 11, 3, 5,
    -- layer=1 filter=66 channel=3
    2, -1, -3, 6, 7, 1, 4, -2, 6,
    -- layer=1 filter=66 channel=4
    -1, 0, 5, 0, 0, 6, -3, 4, -2,
    -- layer=1 filter=66 channel=5
    -4, -17, 5, -11, -5, -6, -1, 0, -13,
    -- layer=1 filter=66 channel=6
    -5, -8, -25, -7, -14, -5, -16, -23, -21,
    -- layer=1 filter=66 channel=7
    0, -6, 7, -14, 0, 18, -8, -2, -4,
    -- layer=1 filter=66 channel=8
    -5, 0, 0, -3, -8, -11, 2, -3, -18,
    -- layer=1 filter=66 channel=9
    -14, -6, -5, -1, -10, -13, -22, -8, 5,
    -- layer=1 filter=66 channel=10
    -8, -11, 16, -21, 4, 3, -7, -20, -7,
    -- layer=1 filter=66 channel=11
    -3, 4, -12, -12, 5, -5, 4, -5, 4,
    -- layer=1 filter=66 channel=12
    -5, -10, -23, -34, -3, 12, 3, -12, -1,
    -- layer=1 filter=66 channel=13
    -17, -4, -9, -6, -17, -8, -14, -19, -28,
    -- layer=1 filter=66 channel=14
    15, -6, 7, -7, -10, 19, -5, -1, 6,
    -- layer=1 filter=66 channel=15
    -12, -15, -19, -6, -10, 0, -24, -7, -8,
    -- layer=1 filter=66 channel=16
    0, -7, 0, -15, -5, -4, 0, -7, -15,
    -- layer=1 filter=66 channel=17
    -9, -5, -9, -1, -9, -6, 1, -5, -16,
    -- layer=1 filter=66 channel=18
    -16, 2, -11, -2, -23, -20, -17, -22, 4,
    -- layer=1 filter=66 channel=19
    -3, 0, -11, -17, -1, 0, 2, -16, 0,
    -- layer=1 filter=66 channel=20
    -1, -1, -8, -1, -8, -2, -20, -4, -19,
    -- layer=1 filter=66 channel=21
    -10, -23, -11, 1, -16, -4, -6, 2, 1,
    -- layer=1 filter=66 channel=22
    -1, -21, -17, -9, -13, 0, -1, -17, -15,
    -- layer=1 filter=66 channel=23
    3, 1, 0, 3, -6, 8, -5, -15, -7,
    -- layer=1 filter=66 channel=24
    -6, -5, -9, -2, -10, -10, -12, -13, -17,
    -- layer=1 filter=66 channel=25
    -6, -11, 12, -17, -11, 6, 7, -11, -13,
    -- layer=1 filter=66 channel=26
    -2, 5, 1, -10, -11, -11, -20, -11, -19,
    -- layer=1 filter=66 channel=27
    0, -9, 7, -2, 6, -3, -3, 3, 8,
    -- layer=1 filter=66 channel=28
    1, -11, 8, -6, -21, -7, -16, -15, -15,
    -- layer=1 filter=66 channel=29
    -10, 5, -11, -3, 0, -4, -4, -1, 1,
    -- layer=1 filter=66 channel=30
    -6, -9, -12, -7, -10, -12, 7, -8, -18,
    -- layer=1 filter=66 channel=31
    -13, -3, -6, -3, -17, -9, -14, -23, -12,
    -- layer=1 filter=66 channel=32
    -6, 2, -4, -2, -2, -6, -18, -11, -3,
    -- layer=1 filter=66 channel=33
    1, -5, -4, 2, 3, -6, -10, -4, 0,
    -- layer=1 filter=66 channel=34
    -7, -1, 1, 4, 5, 3, -1, -4, 0,
    -- layer=1 filter=66 channel=35
    -12, -10, 2, -3, -3, 1, 7, -3, -3,
    -- layer=1 filter=66 channel=36
    -1, -8, -7, -13, -13, -2, -14, 0, -8,
    -- layer=1 filter=66 channel=37
    3, -3, 3, -20, -7, -8, 6, 1, -27,
    -- layer=1 filter=66 channel=38
    -8, -8, -4, -1, -11, -25, -9, -16, -19,
    -- layer=1 filter=66 channel=39
    -2, -15, -11, -9, -13, -9, -15, -5, -2,
    -- layer=1 filter=66 channel=40
    -11, -13, -10, -18, -11, 1, -11, -15, -11,
    -- layer=1 filter=66 channel=41
    -4, 4, 3, 8, 0, 0, -7, 5, 15,
    -- layer=1 filter=66 channel=42
    -3, 0, 1, 10, -8, -6, 5, -4, 0,
    -- layer=1 filter=66 channel=43
    0, -7, -7, -14, -19, -7, -12, 2, -14,
    -- layer=1 filter=66 channel=44
    -10, -7, -3, -19, 1, 1, -22, 13, 3,
    -- layer=1 filter=66 channel=45
    -3, -14, -13, -10, -10, -21, -13, -7, -11,
    -- layer=1 filter=66 channel=46
    0, -12, 0, -17, -12, -10, 5, -17, -16,
    -- layer=1 filter=66 channel=47
    -12, 1, 4, 7, 0, -5, -11, -3, -4,
    -- layer=1 filter=66 channel=48
    -15, 0, -16, -7, -12, -2, -13, -17, -4,
    -- layer=1 filter=66 channel=49
    -4, -15, -4, 2, -8, -16, -11, -9, -16,
    -- layer=1 filter=66 channel=50
    -4, 0, 8, 0, -8, -8, -8, 6, -4,
    -- layer=1 filter=66 channel=51
    0, -4, 0, 0, -16, -7, -19, -9, -3,
    -- layer=1 filter=66 channel=52
    -5, 4, 4, -4, 7, 2, 1, -6, -8,
    -- layer=1 filter=66 channel=53
    -8, 1, 7, -11, -8, 1, -8, -6, 6,
    -- layer=1 filter=66 channel=54
    8, -17, 14, -23, -3, 8, 11, -25, -14,
    -- layer=1 filter=66 channel=55
    3, 1, 0, -1, 8, 3, -4, 1, 9,
    -- layer=1 filter=66 channel=56
    -3, -5, 2, -1, -1, -3, -11, 2, -11,
    -- layer=1 filter=66 channel=57
    -1, -12, 9, -13, -4, 7, -3, -10, -4,
    -- layer=1 filter=66 channel=58
    2, 0, -2, -10, -2, 12, -5, -20, 0,
    -- layer=1 filter=66 channel=59
    -5, -11, 5, 4, -2, -5, 6, -4, -2,
    -- layer=1 filter=66 channel=60
    -11, 1, -2, -9, 5, -7, 0, 2, 7,
    -- layer=1 filter=66 channel=61
    4, -3, 9, -10, -2, 7, 9, 4, -8,
    -- layer=1 filter=66 channel=62
    0, -16, -8, -22, 6, -12, 8, -7, -15,
    -- layer=1 filter=66 channel=63
    -14, 6, -9, 0, 0, -11, -6, -9, -4,
    -- layer=1 filter=66 channel=64
    6, -11, 0, 2, -2, -12, -11, -12, -5,
    -- layer=1 filter=66 channel=65
    2, -10, -8, -5, -10, -9, -11, -2, -1,
    -- layer=1 filter=66 channel=66
    0, -8, 4, 0, 1, 1, -13, 2, -6,
    -- layer=1 filter=66 channel=67
    12, 8, 3, 15, 15, 5, 15, 18, 4,
    -- layer=1 filter=66 channel=68
    -22, -3, -15, -10, 0, -1, -20, 3, -4,
    -- layer=1 filter=66 channel=69
    -16, -5, -18, -1, -15, -13, 0, -1, -25,
    -- layer=1 filter=66 channel=70
    -11, -17, 3, -5, 7, -16, -21, -13, -8,
    -- layer=1 filter=66 channel=71
    8, 4, -13, -6, -4, -12, 2, -4, 2,
    -- layer=1 filter=66 channel=72
    -4, 4, -3, -3, -12, 8, 6, -13, -7,
    -- layer=1 filter=66 channel=73
    8, -2, -11, 0, 2, -1, -1, -10, -11,
    -- layer=1 filter=66 channel=74
    -7, -2, -2, -15, -10, -2, -10, -6, -12,
    -- layer=1 filter=66 channel=75
    -8, 4, -7, -19, 0, 7, 2, -20, -1,
    -- layer=1 filter=66 channel=76
    -12, -4, 0, -5, -6, -11, -11, -9, 7,
    -- layer=1 filter=66 channel=77
    -11, -2, -6, -5, -8, -8, -12, 0, -15,
    -- layer=1 filter=66 channel=78
    -4, -12, -6, -7, 5, -9, -4, 8, 5,
    -- layer=1 filter=66 channel=79
    -14, -12, -6, -11, -13, -5, -4, -4, -17,
    -- layer=1 filter=66 channel=80
    -4, 3, 5, -3, -1, 10, -10, -2, 2,
    -- layer=1 filter=66 channel=81
    5, 4, -2, 2, 0, -6, -8, -13, -2,
    -- layer=1 filter=66 channel=82
    -12, -15, -4, -7, -4, -2, -11, -10, -3,
    -- layer=1 filter=66 channel=83
    -2, 5, -7, -8, 0, -8, -3, -7, -15,
    -- layer=1 filter=66 channel=84
    -14, 4, -9, 1, -10, -22, -14, -21, -19,
    -- layer=1 filter=66 channel=85
    -12, -9, -10, 2, -7, -2, -3, -15, 5,
    -- layer=1 filter=66 channel=86
    -12, -6, 9, -4, -1, -2, -4, -13, -11,
    -- layer=1 filter=66 channel=87
    -17, 5, 0, 0, -21, -15, -6, -24, 1,
    -- layer=1 filter=66 channel=88
    -6, -15, 2, -16, 0, -18, -4, -9, 4,
    -- layer=1 filter=66 channel=89
    -2, 1, -3, 1, -4, -1, -20, 1, 2,
    -- layer=1 filter=66 channel=90
    -21, -4, -1, -4, 1, -3, -29, 3, -4,
    -- layer=1 filter=66 channel=91
    -5, -17, -3, -16, -10, -19, -13, -11, -13,
    -- layer=1 filter=66 channel=92
    -1, -3, -2, 2, -3, 4, -8, -3, -10,
    -- layer=1 filter=66 channel=93
    -3, -20, -6, -17, -8, -8, -1, -10, -9,
    -- layer=1 filter=66 channel=94
    -1, -15, -2, 3, -12, -3, 2, -9, -11,
    -- layer=1 filter=66 channel=95
    -2, -6, -4, -3, -25, -15, -3, -23, -6,
    -- layer=1 filter=66 channel=96
    6, 7, -2, -5, 4, -7, 8, 0, 8,
    -- layer=1 filter=66 channel=97
    -8, -23, -12, -7, -13, -14, -8, -10, -5,
    -- layer=1 filter=66 channel=98
    -11, -20, -6, -16, -9, -7, 2, -16, -22,
    -- layer=1 filter=66 channel=99
    0, -1, 0, -4, -1, -13, 1, -12, -4,
    -- layer=1 filter=66 channel=100
    -13, 1, -8, -5, -2, -5, -8, 12, 2,
    -- layer=1 filter=66 channel=101
    -2, -7, -8, -2, -11, -17, -13, -16, 0,
    -- layer=1 filter=66 channel=102
    -4, 6, -12, 9, -1, 0, 13, 4, 7,
    -- layer=1 filter=66 channel=103
    1, 9, 3, 0, -11, 4, -7, -1, 11,
    -- layer=1 filter=66 channel=104
    7, -9, 0, -3, -10, -5, -10, 9, -2,
    -- layer=1 filter=66 channel=105
    -17, -9, 4, -8, -18, 0, -8, 0, -11,
    -- layer=1 filter=66 channel=106
    -16, 2, -22, 3, -9, -9, -24, -12, -12,
    -- layer=1 filter=66 channel=107
    1, -5, 0, 4, 6, 6, -2, 6, 3,
    -- layer=1 filter=66 channel=108
    -11, 4, -4, 0, 3, -5, -24, 10, -2,
    -- layer=1 filter=66 channel=109
    6, 5, 4, 7, -9, -2, 1, 3, -7,
    -- layer=1 filter=66 channel=110
    6, -5, 0, -2, -7, 0, -11, -2, 0,
    -- layer=1 filter=66 channel=111
    -12, -4, -16, 8, -18, 2, -3, -23, -7,
    -- layer=1 filter=66 channel=112
    6, -3, -9, -10, -3, -13, 2, -18, -5,
    -- layer=1 filter=66 channel=113
    -8, -11, 1, -4, -3, -2, 7, -6, 3,
    -- layer=1 filter=66 channel=114
    -2, -19, -7, 4, -2, -14, -7, -14, -22,
    -- layer=1 filter=66 channel=115
    -5, -6, -9, -16, -7, 6, 0, -9, -3,
    -- layer=1 filter=66 channel=116
    0, -4, -3, 0, 6, -6, 0, 9, 10,
    -- layer=1 filter=66 channel=117
    -18, -4, 0, 0, 2, -1, 0, -23, -28,
    -- layer=1 filter=66 channel=118
    -20, -1, -5, -8, -7, -8, -16, -12, -8,
    -- layer=1 filter=66 channel=119
    -16, -7, -8, -6, -3, -8, -24, -9, -9,
    -- layer=1 filter=66 channel=120
    -12, -16, -1, -17, -7, 2, 0, -7, -18,
    -- layer=1 filter=66 channel=121
    -21, -3, -13, -8, 2, -1, 8, -17, 4,
    -- layer=1 filter=66 channel=122
    2, 0, -2, 2, 3, -6, 3, 7, 1,
    -- layer=1 filter=66 channel=123
    -16, -8, -12, -7, 2, -2, 4, -2, 16,
    -- layer=1 filter=66 channel=124
    -9, 0, 4, -11, 5, -11, 5, -1, 6,
    -- layer=1 filter=66 channel=125
    -16, -11, -9, -9, 0, -12, -2, -6, -11,
    -- layer=1 filter=66 channel=126
    -5, -11, -6, -13, -20, -4, -3, -17, -3,
    -- layer=1 filter=66 channel=127
    -7, -8, -1, -1, -17, -9, -10, -20, -4,
    -- layer=1 filter=67 channel=0
    -6, 1, -7, -2, -6, -5, -2, 7, 6,
    -- layer=1 filter=67 channel=1
    0, 9, 5, -36, -22, -29, -30, -27, 2,
    -- layer=1 filter=67 channel=2
    -8, 30, 8, 2, 7, 10, 16, 28, 19,
    -- layer=1 filter=67 channel=3
    13, 4, 0, 16, 13, 0, 3, 12, -3,
    -- layer=1 filter=67 channel=4
    11, -7, 1, 2, 5, -1, 2, -7, 6,
    -- layer=1 filter=67 channel=5
    3, 12, 19, -43, -7, -26, -30, -41, -35,
    -- layer=1 filter=67 channel=6
    33, 48, 57, 29, 25, 78, 34, 7, -19,
    -- layer=1 filter=67 channel=7
    16, 74, 55, -10, 48, 12, 29, 28, 23,
    -- layer=1 filter=67 channel=8
    -24, -3, -9, -58, -36, -36, -38, -14, -11,
    -- layer=1 filter=67 channel=9
    -5, -11, -31, -17, -9, -7, -24, -5, -31,
    -- layer=1 filter=67 channel=10
    22, 59, 44, 0, 39, 11, 19, 13, 23,
    -- layer=1 filter=67 channel=11
    14, 8, -8, 21, 36, 21, 27, 28, 13,
    -- layer=1 filter=67 channel=12
    -32, 43, 16, -31, -19, 26, 73, 12, 43,
    -- layer=1 filter=67 channel=13
    -16, -13, 11, -4, -22, -8, -25, -23, -12,
    -- layer=1 filter=67 channel=14
    8, 22, 49, -30, 0, 17, -2, -9, 35,
    -- layer=1 filter=67 channel=15
    5, 20, 59, -30, 8, 8, -33, -29, -12,
    -- layer=1 filter=67 channel=16
    -18, -22, -29, -60, -36, -25, -38, -24, -55,
    -- layer=1 filter=67 channel=17
    -20, -19, -20, -6, -18, -18, -14, 0, -14,
    -- layer=1 filter=67 channel=18
    1, -25, -19, 0, 18, -7, -5, 11, -3,
    -- layer=1 filter=67 channel=19
    -14, -45, -44, -59, -84, -30, -46, -64, -95,
    -- layer=1 filter=67 channel=20
    -13, -20, -14, -39, -40, -19, -16, -32, -37,
    -- layer=1 filter=67 channel=21
    23, 17, 30, 6, 6, 12, 3, -6, 6,
    -- layer=1 filter=67 channel=22
    -28, -26, 19, -5, -58, -35, -11, -16, -3,
    -- layer=1 filter=67 channel=23
    -11, 34, 33, -10, 42, 6, -16, 45, 18,
    -- layer=1 filter=67 channel=24
    30, 56, 38, 2, 24, 48, 2, -5, 16,
    -- layer=1 filter=67 channel=25
    5, 28, -2, -44, -1, -19, 8, 16, -9,
    -- layer=1 filter=67 channel=26
    2, 28, 10, -6, 11, 6, -17, 8, 0,
    -- layer=1 filter=67 channel=27
    45, 47, 40, 61, 65, 52, 68, 56, 39,
    -- layer=1 filter=67 channel=28
    9, 33, 40, 10, 21, 9, 20, 24, 9,
    -- layer=1 filter=67 channel=29
    30, 25, 14, 33, 1, 4, 4, -5, -3,
    -- layer=1 filter=67 channel=30
    -33, -47, -48, -67, -48, -43, -65, -61, -64,
    -- layer=1 filter=67 channel=31
    0, -12, -12, -29, -14, -5, 7, -12, 25,
    -- layer=1 filter=67 channel=32
    15, 17, 24, 13, -3, 1, -44, 17, 17,
    -- layer=1 filter=67 channel=33
    11, 23, 6, 8, 15, 27, 16, 22, 19,
    -- layer=1 filter=67 channel=34
    28, 18, 14, 21, 19, 18, 13, 15, -8,
    -- layer=1 filter=67 channel=35
    20, 17, 8, 1, 13, 16, 12, 11, 8,
    -- layer=1 filter=67 channel=36
    24, 7, -4, 32, 22, 19, 32, 38, 32,
    -- layer=1 filter=67 channel=37
    6, 9, -4, -23, -5, -12, -11, -31, -65,
    -- layer=1 filter=67 channel=38
    -9, 0, 9, -26, -13, 13, -6, -26, -20,
    -- layer=1 filter=67 channel=39
    -1, 9, -3, 9, 5, 0, 15, 17, 6,
    -- layer=1 filter=67 channel=40
    -56, -27, -9, -60, -27, -24, -19, -37, -34,
    -- layer=1 filter=67 channel=41
    26, 31, 18, 34, -11, 0, -26, -8, -2,
    -- layer=1 filter=67 channel=42
    -4, -11, -6, -19, -21, -9, 0, 4, 0,
    -- layer=1 filter=67 channel=43
    -16, 3, 5, -46, 13, -40, 2, -6, -29,
    -- layer=1 filter=67 channel=44
    5, 39, 36, 7, 28, 18, -21, 25, 16,
    -- layer=1 filter=67 channel=45
    -22, 31, 27, -34, 5, 11, -35, -18, -9,
    -- layer=1 filter=67 channel=46
    -3, -21, 29, -62, -44, -5, -63, -49, -88,
    -- layer=1 filter=67 channel=47
    -9, 33, 40, -8, 10, -21, -20, 13, -4,
    -- layer=1 filter=67 channel=48
    13, 28, 22, -4, 24, 14, -6, -4, -8,
    -- layer=1 filter=67 channel=49
    16, 18, 32, -2, 10, 25, -15, -18, -16,
    -- layer=1 filter=67 channel=50
    23, 7, -2, 4, -8, 19, -3, 15, 7,
    -- layer=1 filter=67 channel=51
    13, 18, 20, -13, 0, -10, 1, -16, -8,
    -- layer=1 filter=67 channel=52
    -3, -2, -12, -8, -17, 20, -9, -17, -1,
    -- layer=1 filter=67 channel=53
    -8, -7, 6, -8, -6, -5, 2, 5, 5,
    -- layer=1 filter=67 channel=54
    5, 39, 3, -10, 4, 16, 14, 31, -10,
    -- layer=1 filter=67 channel=55
    30, 27, 7, 43, 46, 17, 23, 36, 29,
    -- layer=1 filter=67 channel=56
    -6, 6, 12, 2, -8, 5, 4, -7, 7,
    -- layer=1 filter=67 channel=57
    -18, 11, 29, -22, 18, -3, -8, -20, 5,
    -- layer=1 filter=67 channel=58
    -19, 59, 9, -24, 47, 9, 1, 40, 3,
    -- layer=1 filter=67 channel=59
    -1, -12, -1, 3, 4, 5, -18, -13, 0,
    -- layer=1 filter=67 channel=60
    -3, -4, 0, -2, -15, 18, -17, -12, 15,
    -- layer=1 filter=67 channel=61
    5, 7, 7, -3, 6, -7, -3, 11, -1,
    -- layer=1 filter=67 channel=62
    -44, -7, -30, -97, -45, -35, -31, -32, -34,
    -- layer=1 filter=67 channel=63
    32, -8, -5, 29, 31, 11, 30, 29, 26,
    -- layer=1 filter=67 channel=64
    -9, -7, 30, 11, -5, -7, 0, 0, 4,
    -- layer=1 filter=67 channel=65
    22, 25, 16, -1, 19, 2, 2, 0, -15,
    -- layer=1 filter=67 channel=66
    1, 1, -7, 11, 16, 10, 10, 16, 10,
    -- layer=1 filter=67 channel=67
    70, 71, 54, 28, 72, 83, 55, 41, 41,
    -- layer=1 filter=67 channel=68
    25, 46, 36, 7, 36, 36, -21, 37, 41,
    -- layer=1 filter=67 channel=69
    -33, 42, 13, -58, 7, 2, -23, -20, -8,
    -- layer=1 filter=67 channel=70
    48, 95, 59, 59, 67, 112, 45, 38, 74,
    -- layer=1 filter=67 channel=71
    39, 30, 42, 15, 34, 27, 12, 10, 6,
    -- layer=1 filter=67 channel=72
    -13, -10, -14, -4, -17, 8, -18, -19, -20,
    -- layer=1 filter=67 channel=73
    16, 7, 9, 9, 0, 18, 12, 16, 7,
    -- layer=1 filter=67 channel=74
    -33, -9, 21, -42, 13, 47, -24, -8, 0,
    -- layer=1 filter=67 channel=75
    -25, -14, 10, -40, -18, -26, -8, -12, -20,
    -- layer=1 filter=67 channel=76
    24, 3, -5, -4, 4, 2, -35, 11, -5,
    -- layer=1 filter=67 channel=77
    18, 39, 23, 2, 28, 12, -7, 2, -1,
    -- layer=1 filter=67 channel=78
    14, 1, 2, -9, -3, 13, 0, 13, 12,
    -- layer=1 filter=67 channel=79
    -30, -18, -38, -82, -35, -48, -38, -47, -62,
    -- layer=1 filter=67 channel=80
    -12, 0, -6, -3, -4, -17, 2, -1, 5,
    -- layer=1 filter=67 channel=81
    20, 23, 26, 14, 34, 16, 5, 18, -2,
    -- layer=1 filter=67 channel=82
    10, 27, 43, 28, 25, 16, 15, 7, 5,
    -- layer=1 filter=67 channel=83
    -1, 48, 8, -10, 13, -18, -3, -8, -4,
    -- layer=1 filter=67 channel=84
    -28, -52, -31, -17, -20, -15, -45, -2, -2,
    -- layer=1 filter=67 channel=85
    -24, 34, -3, 12, 21, 13, -35, 44, -7,
    -- layer=1 filter=67 channel=86
    10, -11, -16, 12, -5, -12, 3, 5, -6,
    -- layer=1 filter=67 channel=87
    -29, 2, -19, -41, -35, -38, -50, -35, -39,
    -- layer=1 filter=67 channel=88
    29, 40, 50, 4, 22, 46, -21, -7, -4,
    -- layer=1 filter=67 channel=89
    17, 27, 36, 7, 7, 14, -16, -7, 1,
    -- layer=1 filter=67 channel=90
    23, 64, 43, -5, 45, 25, -17, 30, 21,
    -- layer=1 filter=67 channel=91
    -21, -28, -18, -10, -42, -21, -4, -41, -41,
    -- layer=1 filter=67 channel=92
    41, 65, 7, 17, 37, -33, -9, 1, -11,
    -- layer=1 filter=67 channel=93
    7, 10, 3, -1, 4, -1, -8, -14, 2,
    -- layer=1 filter=67 channel=94
    -15, -25, -25, 0, -6, -13, -11, -12, -15,
    -- layer=1 filter=67 channel=95
    -34, -50, -32, -57, -17, -31, -61, -12, -21,
    -- layer=1 filter=67 channel=96
    13, 4, 8, 29, 18, -2, 20, 22, 6,
    -- layer=1 filter=67 channel=97
    6, -4, -7, 0, 0, -9, 8, 0, 1,
    -- layer=1 filter=67 channel=98
    -43, -36, -22, -52, -40, -55, -48, -40, -31,
    -- layer=1 filter=67 channel=99
    -27, 2, 50, -5, -11, 17, 8, -13, 54,
    -- layer=1 filter=67 channel=100
    25, 5, -2, 28, 24, 14, 24, 32, 7,
    -- layer=1 filter=67 channel=101
    -17, -21, -5, -19, -33, -3, -17, -33, -21,
    -- layer=1 filter=67 channel=102
    -7, -37, -36, -14, -34, -19, -22, -32, -30,
    -- layer=1 filter=67 channel=103
    26, 20, -8, 23, 39, 17, 24, 20, 12,
    -- layer=1 filter=67 channel=104
    -26, 25, 28, -12, 1, 0, -14, 17, 36,
    -- layer=1 filter=67 channel=105
    -11, -7, -13, -7, -1, 0, -5, 7, 6,
    -- layer=1 filter=67 channel=106
    -30, 6, 13, -19, -25, 6, -58, -21, -10,
    -- layer=1 filter=67 channel=107
    -9, 12, -8, 9, 1, -2, -1, -12, -3,
    -- layer=1 filter=67 channel=108
    25, 71, 65, 25, 39, 47, -22, 12, 53,
    -- layer=1 filter=67 channel=109
    -2, 6, -1, 2, 8, 0, 3, 6, 8,
    -- layer=1 filter=67 channel=110
    0, -1, -6, -17, -8, -9, -22, -9, -12,
    -- layer=1 filter=67 channel=111
    -27, -53, -44, -49, -36, -38, -55, -19, -33,
    -- layer=1 filter=67 channel=112
    -13, -20, -10, -33, -26, -13, -18, 26, 14,
    -- layer=1 filter=67 channel=113
    -6, -16, -12, -34, -31, -16, -30, -29, -14,
    -- layer=1 filter=67 channel=114
    14, 47, 34, 1, 29, 15, 22, 3, -11,
    -- layer=1 filter=67 channel=115
    -25, 0, -20, -14, 1, -19, 1, 11, -7,
    -- layer=1 filter=67 channel=116
    4, 9, -7, 8, -4, -5, -1, -1, -5,
    -- layer=1 filter=67 channel=117
    -37, 1, -9, -59, -43, -59, -27, -2, 17,
    -- layer=1 filter=67 channel=118
    -46, -53, -23, -65, -27, -14, -39, -16, -36,
    -- layer=1 filter=67 channel=119
    34, 51, 43, 10, 25, 38, -25, 24, 32,
    -- layer=1 filter=67 channel=120
    30, 44, 9, 0, 10, -7, 20, -6, -27,
    -- layer=1 filter=67 channel=121
    40, 33, 34, 27, 44, 44, 57, 40, 26,
    -- layer=1 filter=67 channel=122
    1, -5, -5, -9, -1, 9, 9, 4, -6,
    -- layer=1 filter=67 channel=123
    41, 40, 35, 46, 52, 41, 37, 48, 33,
    -- layer=1 filter=67 channel=124
    9, 0, 5, -6, -1, -2, -1, -1, -16,
    -- layer=1 filter=67 channel=125
    59, 67, 65, 43, 95, 80, 52, 28, 71,
    -- layer=1 filter=67 channel=126
    -6, 3, -8, -4, -33, -43, -43, -56, 7,
    -- layer=1 filter=67 channel=127
    -52, -81, -53, -76, -40, -50, -52, -37, -51,
    -- layer=1 filter=68 channel=0
    -18, -17, -5, 2, -7, 11, 5, -2, 14,
    -- layer=1 filter=68 channel=1
    -9, 5, -21, 6, 4, 9, 0, 1, 12,
    -- layer=1 filter=68 channel=2
    32, 36, 26, 32, 39, 26, 36, 42, -5,
    -- layer=1 filter=68 channel=3
    0, -10, -5, -4, -3, 1, -17, 0, -14,
    -- layer=1 filter=68 channel=4
    -2, -9, -2, 3, -8, 6, -1, -2, 6,
    -- layer=1 filter=68 channel=5
    1, -1, -34, -13, -3, 9, -3, -3, 11,
    -- layer=1 filter=68 channel=6
    -6, -12, -6, -15, -5, -4, -25, -20, -19,
    -- layer=1 filter=68 channel=7
    3, 41, 30, 30, 28, 25, 6, 34, 10,
    -- layer=1 filter=68 channel=8
    -3, 0, -23, 12, 2, 15, -7, 2, -3,
    -- layer=1 filter=68 channel=9
    9, -42, -2, -2, -13, -13, -7, -21, -16,
    -- layer=1 filter=68 channel=10
    14, 38, 29, 37, 24, 29, 8, 26, -7,
    -- layer=1 filter=68 channel=11
    -15, -28, -26, -8, -13, -12, -16, -3, -2,
    -- layer=1 filter=68 channel=12
    -45, -22, -2, -20, -33, -62, -21, -80, -8,
    -- layer=1 filter=68 channel=13
    11, 11, 6, 8, 23, 5, -5, -6, 1,
    -- layer=1 filter=68 channel=14
    -16, 18, -5, -12, -28, -14, 2, -21, -27,
    -- layer=1 filter=68 channel=15
    7, 8, -24, 3, 9, -25, -18, 2, -19,
    -- layer=1 filter=68 channel=16
    19, 28, -9, 15, 8, 17, 13, 3, 6,
    -- layer=1 filter=68 channel=17
    -9, 2, 7, 0, 17, 11, 15, 13, 6,
    -- layer=1 filter=68 channel=18
    -34, -38, -36, -24, 0, -4, -12, -20, 22,
    -- layer=1 filter=68 channel=19
    4, -60, -50, -22, -45, -25, 22, 14, 35,
    -- layer=1 filter=68 channel=20
    16, 21, 20, 8, 21, 19, 5, 19, -2,
    -- layer=1 filter=68 channel=21
    3, 11, 4, 4, -4, -8, 4, -15, 1,
    -- layer=1 filter=68 channel=22
    12, 13, 0, 18, 12, 19, 8, 6, -6,
    -- layer=1 filter=68 channel=23
    -22, -2, -1, -9, -1, -2, 1, -9, -8,
    -- layer=1 filter=68 channel=24
    15, -31, -19, -18, -19, -15, -17, -10, -18,
    -- layer=1 filter=68 channel=25
    15, 43, -4, 30, 17, 32, 0, 35, 9,
    -- layer=1 filter=68 channel=26
    4, -5, -9, 1, 0, -23, -6, 12, -2,
    -- layer=1 filter=68 channel=27
    -24, -20, -14, -32, -26, -37, -25, -40, -60,
    -- layer=1 filter=68 channel=28
    3, 27, 14, 30, 13, 18, 15, 26, -7,
    -- layer=1 filter=68 channel=29
    -24, -11, -4, -10, -14, 4, -2, 3, -5,
    -- layer=1 filter=68 channel=30
    -41, -58, -49, -40, -35, -44, -15, -21, 5,
    -- layer=1 filter=68 channel=31
    -27, -1, -20, -15, -21, -23, -30, -37, -10,
    -- layer=1 filter=68 channel=32
    -10, 7, -7, -11, 14, -45, -26, 17, -2,
    -- layer=1 filter=68 channel=33
    2, 0, -1, 11, 6, 0, 0, 8, 12,
    -- layer=1 filter=68 channel=34
    -22, -22, -3, -39, -9, -13, -37, -28, -17,
    -- layer=1 filter=68 channel=35
    20, 9, -1, 10, 20, 9, 9, 16, 0,
    -- layer=1 filter=68 channel=36
    -37, -39, -35, -33, -11, -20, -13, -9, -7,
    -- layer=1 filter=68 channel=37
    6, 14, -35, -5, 6, 13, -1, 10, 2,
    -- layer=1 filter=68 channel=38
    19, 9, 4, 19, 5, -3, 12, 3, 0,
    -- layer=1 filter=68 channel=39
    -2, -4, 0, -26, -18, -11, -12, -10, 0,
    -- layer=1 filter=68 channel=40
    6, -4, 0, -20, -13, -18, 1, -29, -7,
    -- layer=1 filter=68 channel=41
    -9, -38, 23, -33, 12, -44, -22, -20, -19,
    -- layer=1 filter=68 channel=42
    46, 47, 17, 39, 28, 33, 58, 37, -3,
    -- layer=1 filter=68 channel=43
    13, 21, -21, 22, -4, 26, -8, 6, -8,
    -- layer=1 filter=68 channel=44
    -7, -8, -12, -8, 16, -42, -13, 27, -8,
    -- layer=1 filter=68 channel=45
    11, 4, -5, -2, 10, -9, -8, 6, -22,
    -- layer=1 filter=68 channel=46
    0, -31, -29, -1, -2, -16, 18, 15, 21,
    -- layer=1 filter=68 channel=47
    -8, -4, -3, -1, 27, -17, -15, -12, -13,
    -- layer=1 filter=68 channel=48
    7, -3, 13, 16, -10, 2, 5, -9, -10,
    -- layer=1 filter=68 channel=49
    22, 11, 14, 7, -3, -5, 0, -22, -10,
    -- layer=1 filter=68 channel=50
    -2, -5, -2, -12, -10, -1, 2, -10, -6,
    -- layer=1 filter=68 channel=51
    3, 11, 17, 23, 7, 0, 1, -2, -11,
    -- layer=1 filter=68 channel=52
    -2, -3, 9, -16, -2, -2, 5, -7, 6,
    -- layer=1 filter=68 channel=53
    10, 7, 0, 18, 18, 17, -1, 13, 14,
    -- layer=1 filter=68 channel=54
    15, 35, -5, 12, 4, 29, -7, 11, -18,
    -- layer=1 filter=68 channel=55
    -16, -26, -32, -33, -24, -21, -21, -13, -44,
    -- layer=1 filter=68 channel=56
    7, 0, 1, -3, -1, 0, 5, 2, 5,
    -- layer=1 filter=68 channel=57
    11, 16, 22, 25, 14, 26, 3, 14, -7,
    -- layer=1 filter=68 channel=58
    5, 8, 6, -9, 1, 10, -13, 21, 2,
    -- layer=1 filter=68 channel=59
    1, 12, 16, -4, 5, 12, -4, 11, 5,
    -- layer=1 filter=68 channel=60
    11, 21, 6, 6, 0, -1, -1, -1, -6,
    -- layer=1 filter=68 channel=61
    6, -4, -8, -1, -3, -2, -5, -10, 0,
    -- layer=1 filter=68 channel=62
    9, 15, -21, 9, -3, 13, 8, 0, -6,
    -- layer=1 filter=68 channel=63
    -42, -37, -25, -23, -23, -29, -7, -6, 8,
    -- layer=1 filter=68 channel=64
    0, 10, 13, 10, 8, -4, -1, -5, 9,
    -- layer=1 filter=68 channel=65
    5, -7, -13, 3, -6, 0, -1, 6, 0,
    -- layer=1 filter=68 channel=66
    -32, -25, -21, -12, -19, 2, -7, -5, 3,
    -- layer=1 filter=68 channel=67
    9, -7, 9, -3, -36, -18, -21, -46, -32,
    -- layer=1 filter=68 channel=68
    0, -7, -15, -2, 11, -30, 0, 44, -5,
    -- layer=1 filter=68 channel=69
    11, 3, -18, -8, 12, -6, 5, 6, -19,
    -- layer=1 filter=68 channel=70
    -26, -36, -21, -34, -43, -32, -50, -35, -20,
    -- layer=1 filter=68 channel=71
    -16, -9, -11, -10, -27, -3, -6, -7, -2,
    -- layer=1 filter=68 channel=72
    -21, -71, -60, -44, -27, -37, -14, -37, 5,
    -- layer=1 filter=68 channel=73
    -2, -1, -4, -10, -3, -9, 8, 2, 4,
    -- layer=1 filter=68 channel=74
    -16, -35, -35, -14, 27, -17, -12, 6, 15,
    -- layer=1 filter=68 channel=75
    -44, -4, -45, 21, -42, -65, -1, -68, -35,
    -- layer=1 filter=68 channel=76
    -16, -3, -12, -4, 1, -17, 0, 4, 7,
    -- layer=1 filter=68 channel=77
    0, -1, 2, 6, 3, 2, 11, -1, -6,
    -- layer=1 filter=68 channel=78
    -5, -11, -5, 2, -5, 9, 4, -6, 14,
    -- layer=1 filter=68 channel=79
    5, 24, -3, 21, 15, 12, 4, 20, 4,
    -- layer=1 filter=68 channel=80
    5, 8, -6, -8, -6, 8, 1, -4, -8,
    -- layer=1 filter=68 channel=81
    -4, -18, 0, 0, -18, 0, -9, -6, -9,
    -- layer=1 filter=68 channel=82
    9, 10, 6, 11, -12, 4, 0, -17, 1,
    -- layer=1 filter=68 channel=83
    3, -13, 4, -10, 14, 5, -2, 18, -14,
    -- layer=1 filter=68 channel=84
    -60, -45, -83, -47, -29, -25, -26, -12, 13,
    -- layer=1 filter=68 channel=85
    23, -20, 31, -13, -11, 11, -19, -19, 6,
    -- layer=1 filter=68 channel=86
    -15, -6, 0, -6, -6, 4, -3, 12, 20,
    -- layer=1 filter=68 channel=87
    -2, -64, -63, -55, -35, -48, 0, -31, -11,
    -- layer=1 filter=68 channel=88
    2, 13, 6, -2, -14, -13, -4, -5, -12,
    -- layer=1 filter=68 channel=89
    -7, 0, -6, -11, -9, 0, 2, 7, 2,
    -- layer=1 filter=68 channel=90
    9, -13, -17, 3, 24, -40, -2, 29, -22,
    -- layer=1 filter=68 channel=91
    21, 23, 13, 17, 1, 12, 9, 13, 3,
    -- layer=1 filter=68 channel=92
    16, -50, -58, 18, 23, -110, 2, -11, -54,
    -- layer=1 filter=68 channel=93
    2, -7, 2, -7, -4, 2, -3, 0, 2,
    -- layer=1 filter=68 channel=94
    -10, 1, 5, -11, 6, 13, 8, 0, 17,
    -- layer=1 filter=68 channel=95
    -68, -63, -82, -50, -23, -40, -30, -27, 5,
    -- layer=1 filter=68 channel=96
    -4, -5, 4, -13, 1, -2, -14, -13, -4,
    -- layer=1 filter=68 channel=97
    -25, -16, -11, -2, 5, 6, 0, 15, 13,
    -- layer=1 filter=68 channel=98
    12, 25, 1, 33, 8, 21, 7, 20, 0,
    -- layer=1 filter=68 channel=99
    17, 4, -14, 14, 16, -16, 2, -3, -19,
    -- layer=1 filter=68 channel=100
    -17, -14, -21, -20, -19, -21, -3, 0, -11,
    -- layer=1 filter=68 channel=101
    10, 2, 18, 9, 3, 11, 12, -4, 8,
    -- layer=1 filter=68 channel=102
    -13, -10, -4, 15, 12, 9, 7, 22, 24,
    -- layer=1 filter=68 channel=103
    -13, -19, -7, -16, -12, -6, -8, 3, -2,
    -- layer=1 filter=68 channel=104
    -19, -18, -7, -9, -3, -15, -26, -5, -36,
    -- layer=1 filter=68 channel=105
    -28, -10, -1, -12, 4, -2, 10, -2, 11,
    -- layer=1 filter=68 channel=106
    0, 2, -6, 0, 4, -15, -8, 15, 4,
    -- layer=1 filter=68 channel=107
    -11, 6, -10, -10, -13, -15, -12, -12, -6,
    -- layer=1 filter=68 channel=108
    -4, -12, 13, -19, 31, -27, -21, 21, -13,
    -- layer=1 filter=68 channel=109
    7, -3, -6, -5, 1, -6, -8, 6, 2,
    -- layer=1 filter=68 channel=110
    -4, 7, 8, 4, 7, -1, 4, 8, 13,
    -- layer=1 filter=68 channel=111
    -43, -61, -41, -52, -10, -18, -10, -32, 9,
    -- layer=1 filter=68 channel=112
    -55, -31, -47, -19, -7, 0, -8, -9, 5,
    -- layer=1 filter=68 channel=113
    -8, 3, -3, 3, 8, 12, -23, 3, -16,
    -- layer=1 filter=68 channel=114
    -13, -50, -60, -63, -63, -49, -52, -45, -44,
    -- layer=1 filter=68 channel=115
    -13, -3, 10, 2, -7, 17, -2, 3, 2,
    -- layer=1 filter=68 channel=116
    0, 3, -9, 8, 1, 2, 4, -9, 4,
    -- layer=1 filter=68 channel=117
    -22, -67, -49, -30, -25, -13, 0, -12, -16,
    -- layer=1 filter=68 channel=118
    -41, -70, -49, -33, -14, -21, -14, -12, 7,
    -- layer=1 filter=68 channel=119
    -2, -3, -1, 1, 19, -21, -22, 31, -23,
    -- layer=1 filter=68 channel=120
    9, 14, 10, 7, 5, 3, 1, 2, -3,
    -- layer=1 filter=68 channel=121
    -2, -21, -24, -31, -40, -45, -6, -23, -26,
    -- layer=1 filter=68 channel=122
    8, -5, 5, 3, -3, -6, -1, -8, -9,
    -- layer=1 filter=68 channel=123
    -23, -13, -31, -28, -19, -38, -21, -19, -30,
    -- layer=1 filter=68 channel=124
    -4, 8, -6, -7, 1, 9, -11, -7, 4,
    -- layer=1 filter=68 channel=125
    -1, -1, 12, -17, -15, -18, -29, -14, -11,
    -- layer=1 filter=68 channel=126
    -14, -2, -9, 7, -13, 3, 5, -4, -18,
    -- layer=1 filter=68 channel=127
    -45, -57, -66, -37, -18, -11, -16, -33, 4,
    -- layer=1 filter=69 channel=0
    13, -4, 6, -3, 11, 8, -11, 4, 9,
    -- layer=1 filter=69 channel=1
    9, -7, 13, -11, -8, -15, 20, 8, -11,
    -- layer=1 filter=69 channel=2
    22, 34, 38, 7, -14, 5, 41, 37, 40,
    -- layer=1 filter=69 channel=3
    6, 1, 10, 7, -6, -3, -3, 9, 4,
    -- layer=1 filter=69 channel=4
    7, 6, -11, 0, -9, 5, -6, 0, -5,
    -- layer=1 filter=69 channel=5
    -13, -8, 7, -20, -52, -42, 52, 47, 35,
    -- layer=1 filter=69 channel=6
    -16, -5, -24, 5, 7, 34, 12, 36, 30,
    -- layer=1 filter=69 channel=7
    1, 2, -16, 27, 1, -37, 27, 24, 28,
    -- layer=1 filter=69 channel=8
    6, 26, 12, -17, -13, -13, 45, 13, -31,
    -- layer=1 filter=69 channel=9
    35, 5, 40, 30, 11, 0, -39, 17, -29,
    -- layer=1 filter=69 channel=10
    26, -1, -19, 48, 14, -31, 32, 52, 30,
    -- layer=1 filter=69 channel=11
    -5, -26, -8, -16, -8, -22, 5, -3, -31,
    -- layer=1 filter=69 channel=12
    -17, 60, 46, 72, 39, 25, -23, 14, 34,
    -- layer=1 filter=69 channel=13
    3, 11, 6, -19, 3, 40, -10, -12, -3,
    -- layer=1 filter=69 channel=14
    -20, -32, -14, 24, -1, -32, 22, 9, 3,
    -- layer=1 filter=69 channel=15
    -9, 26, 28, 19, -17, -27, 20, 56, 1,
    -- layer=1 filter=69 channel=16
    5, 21, 28, -24, -36, -36, 20, -4, -28,
    -- layer=1 filter=69 channel=17
    9, 9, 17, -15, 14, 31, -25, -26, -12,
    -- layer=1 filter=69 channel=18
    -15, -25, -1, 11, 11, -43, 39, 57, 67,
    -- layer=1 filter=69 channel=19
    16, 1, 15, 29, -34, -63, 1, 21, -3,
    -- layer=1 filter=69 channel=20
    3, 17, 16, -17, 33, 41, -23, 2, 0,
    -- layer=1 filter=69 channel=21
    11, 1, 14, -27, -7, 19, -14, -28, -6,
    -- layer=1 filter=69 channel=22
    0, 16, 14, -27, 20, 20, -16, -18, -37,
    -- layer=1 filter=69 channel=23
    -17, 14, -12, -6, -62, -24, 25, 20, 10,
    -- layer=1 filter=69 channel=24
    2, 5, 14, -16, -25, -30, -7, -57, -63,
    -- layer=1 filter=69 channel=25
    12, 9, 3, 4, -23, -34, 4, -28, -8,
    -- layer=1 filter=69 channel=26
    19, 18, 28, -11, -39, -27, 6, -48, -64,
    -- layer=1 filter=69 channel=27
    40, 44, 42, 49, 36, 39, 34, 33, 29,
    -- layer=1 filter=69 channel=28
    33, 5, 28, 22, 10, 1, -10, 7, 0,
    -- layer=1 filter=69 channel=29
    20, 18, 32, 27, 27, 26, 17, 22, 24,
    -- layer=1 filter=69 channel=30
    -27, -37, 1, 34, 8, -25, 21, 76, 62,
    -- layer=1 filter=69 channel=31
    -22, -9, -4, 17, -18, -18, 27, 58, 52,
    -- layer=1 filter=69 channel=32
    -12, -44, -15, 17, -55, -62, 14, -7, -28,
    -- layer=1 filter=69 channel=33
    -9, 16, 8, -16, 8, 9, -4, 11, -23,
    -- layer=1 filter=69 channel=34
    -25, 13, 10, -8, 5, 27, 0, 0, 9,
    -- layer=1 filter=69 channel=35
    6, 22, 5, 9, -22, 8, 1, -6, -10,
    -- layer=1 filter=69 channel=36
    -7, -17, -5, -21, -23, -20, -17, -24, -23,
    -- layer=1 filter=69 channel=37
    -13, 15, 5, -49, -73, -57, 35, 26, 23,
    -- layer=1 filter=69 channel=38
    2, 12, 7, 9, 25, 22, -30, 16, 15,
    -- layer=1 filter=69 channel=39
    -8, 5, 9, 7, -13, -18, -3, -24, -41,
    -- layer=1 filter=69 channel=40
    -29, -13, -17, 13, 15, 13, 17, 68, 63,
    -- layer=1 filter=69 channel=41
    -14, -70, -34, 31, -91, -75, 2, -39, -103,
    -- layer=1 filter=69 channel=42
    -8, 17, 39, 11, -4, 3, 23, 19, 25,
    -- layer=1 filter=69 channel=43
    5, 12, 36, -21, -43, -20, 15, -10, -39,
    -- layer=1 filter=69 channel=44
    7, -4, 17, 0, -56, -33, 43, -35, -48,
    -- layer=1 filter=69 channel=45
    0, 2, 26, -19, -5, -15, 6, -13, 0,
    -- layer=1 filter=69 channel=46
    12, 44, 62, 45, 12, -46, 54, 113, 64,
    -- layer=1 filter=69 channel=47
    -22, -11, -54, 9, -64, -34, 42, 19, 21,
    -- layer=1 filter=69 channel=48
    0, 5, -2, 3, 28, 26, -16, -12, 17,
    -- layer=1 filter=69 channel=49
    -2, 3, -24, 10, 0, 16, -2, 11, 2,
    -- layer=1 filter=69 channel=50
    -11, 4, 2, -18, 3, -4, -8, -6, -22,
    -- layer=1 filter=69 channel=51
    0, -11, -17, 23, 15, 23, -22, 14, 19,
    -- layer=1 filter=69 channel=52
    -4, -6, 9, -18, -17, -22, 5, -6, 0,
    -- layer=1 filter=69 channel=53
    -5, 7, 8, 5, 1, -1, 10, 9, 20,
    -- layer=1 filter=69 channel=54
    13, -14, 11, -25, -50, -71, 9, -36, 3,
    -- layer=1 filter=69 channel=55
    -1, -27, -24, 9, -4, -16, 15, -18, -47,
    -- layer=1 filter=69 channel=56
    2, 2, -3, -7, 0, 11, 3, -1, -2,
    -- layer=1 filter=69 channel=57
    10, 12, -16, 28, 27, -8, 9, 45, 33,
    -- layer=1 filter=69 channel=58
    -7, -42, -17, 13, -34, -79, 45, 12, 40,
    -- layer=1 filter=69 channel=59
    11, 13, -5, -2, -2, 0, -1, -20, -7,
    -- layer=1 filter=69 channel=60
    17, 10, 0, 4, 12, 9, 11, 3, 14,
    -- layer=1 filter=69 channel=61
    1, -11, -4, -3, 1, -6, -1, 5, -9,
    -- layer=1 filter=69 channel=62
    3, 8, 30, -40, -35, -38, 23, -21, -60,
    -- layer=1 filter=69 channel=63
    -17, -27, -15, -3, -29, -42, -9, -2, -23,
    -- layer=1 filter=69 channel=64
    17, 0, 4, -20, 0, 11, -4, -11, -13,
    -- layer=1 filter=69 channel=65
    9, 13, 26, -5, 11, 30, -24, -10, 1,
    -- layer=1 filter=69 channel=66
    -10, -4, -10, 11, -14, -14, 0, -8, -23,
    -- layer=1 filter=69 channel=67
    -9, -35, -24, 22, 18, 22, -5, -5, 31,
    -- layer=1 filter=69 channel=68
    14, 8, 19, -14, -57, -39, 24, -29, -35,
    -- layer=1 filter=69 channel=69
    23, 37, 50, -22, -45, -28, 53, 54, 3,
    -- layer=1 filter=69 channel=70
    27, 17, -6, 16, 19, 17, 18, 56, 71,
    -- layer=1 filter=69 channel=71
    13, -4, 19, -5, -15, -21, 13, -17, -27,
    -- layer=1 filter=69 channel=72
    -2, -9, 28, 17, -18, -9, -16, 47, 31,
    -- layer=1 filter=69 channel=73
    -7, -6, -2, -9, 4, -4, 4, 0, -5,
    -- layer=1 filter=69 channel=74
    -23, -2, -2, -4, -44, -22, 8, 19, 33,
    -- layer=1 filter=69 channel=75
    -60, 8, 30, 32, -1, -23, 24, 64, 49,
    -- layer=1 filter=69 channel=76
    14, -21, 15, 4, -3, -8, 17, -18, 24,
    -- layer=1 filter=69 channel=77
    8, -1, 6, -9, 6, 26, -17, -33, -10,
    -- layer=1 filter=69 channel=78
    -3, 0, -12, -13, 5, -9, -7, 2, 13,
    -- layer=1 filter=69 channel=79
    6, 37, 43, -32, -30, -17, 18, -16, -53,
    -- layer=1 filter=69 channel=80
    3, 4, 0, 5, 10, -2, -1, 0, 1,
    -- layer=1 filter=69 channel=81
    20, 26, 36, -11, -31, -3, -16, -67, -42,
    -- layer=1 filter=69 channel=82
    4, 7, 21, -12, 13, 16, -31, -28, 0,
    -- layer=1 filter=69 channel=83
    14, 28, 33, -14, -35, -12, 20, -3, -6,
    -- layer=1 filter=69 channel=84
    -14, -37, -19, 7, -12, -43, 19, 9, 37,
    -- layer=1 filter=69 channel=85
    -41, -1, -8, -16, -51, -34, 3, 8, -6,
    -- layer=1 filter=69 channel=86
    -10, -15, -12, -10, -13, -9, -16, -7, -26,
    -- layer=1 filter=69 channel=87
    43, -17, 22, 37, -8, -38, -21, 19, -4,
    -- layer=1 filter=69 channel=88
    0, 0, 1, -2, 4, 9, -1, -16, 2,
    -- layer=1 filter=69 channel=89
    13, 15, 12, -3, -5, 9, -8, -2, -11,
    -- layer=1 filter=69 channel=90
    9, 16, 33, -22, -43, -16, 36, -12, -51,
    -- layer=1 filter=69 channel=91
    -20, 1, 4, 10, 37, 32, -35, 19, 29,
    -- layer=1 filter=69 channel=92
    21, 35, 35, 16, 22, -9, 17, 45, 18,
    -- layer=1 filter=69 channel=93
    7, 14, 19, -8, 1, 18, -21, -32, -24,
    -- layer=1 filter=69 channel=94
    -11, 6, 1, 7, 15, 1, -6, 2, -2,
    -- layer=1 filter=69 channel=95
    -49, -30, -6, 18, -18, -29, 44, 41, 35,
    -- layer=1 filter=69 channel=96
    0, 15, 14, 13, 8, 12, 16, 19, 12,
    -- layer=1 filter=69 channel=97
    6, 11, 19, -22, -3, 18, -15, -29, -23,
    -- layer=1 filter=69 channel=98
    26, 30, 24, -14, 7, 25, -8, -48, -61,
    -- layer=1 filter=69 channel=99
    32, 0, 6, 25, 21, 3, 20, 64, 40,
    -- layer=1 filter=69 channel=100
    1, 9, 7, -5, -11, -38, -11, 2, -13,
    -- layer=1 filter=69 channel=101
    -4, 15, 6, -1, 16, 32, -10, 3, 27,
    -- layer=1 filter=69 channel=102
    4, -1, 6, 9, 33, 33, -23, 13, 29,
    -- layer=1 filter=69 channel=103
    13, -2, 13, 14, 16, -16, 20, 19, -18,
    -- layer=1 filter=69 channel=104
    15, -11, -18, 1, -35, -20, 16, 24, 25,
    -- layer=1 filter=69 channel=105
    5, 6, -5, 1, -4, 6, -12, -8, -10,
    -- layer=1 filter=69 channel=106
    -14, -4, -4, 0, 3, 22, 4, -10, 16,
    -- layer=1 filter=69 channel=107
    -10, 0, -13, -2, -5, 8, -4, -5, -11,
    -- layer=1 filter=69 channel=108
    24, 0, 12, 25, -50, -40, 33, -6, -41,
    -- layer=1 filter=69 channel=109
    4, -2, 0, 7, -9, 6, -7, 9, 6,
    -- layer=1 filter=69 channel=110
    10, 13, 4, 12, 2, 2, 0, 5, 0,
    -- layer=1 filter=69 channel=111
    0, -21, 3, 37, 10, -21, 46, 47, 69,
    -- layer=1 filter=69 channel=112
    -19, -27, -37, 12, -4, -40, 42, 22, 39,
    -- layer=1 filter=69 channel=113
    -4, 37, 14, -13, 25, 0, -12, 18, 13,
    -- layer=1 filter=69 channel=114
    4, 15, 24, 20, -19, -29, 34, 40, 0,
    -- layer=1 filter=69 channel=115
    0, 9, -23, 13, 10, -5, -5, 8, 0,
    -- layer=1 filter=69 channel=116
    -5, 0, 1, -3, 0, 0, 0, 4, -6,
    -- layer=1 filter=69 channel=117
    37, 9, -9, 60, 58, -2, 67, 64, 109,
    -- layer=1 filter=69 channel=118
    -32, -47, 0, 15, 3, -19, 26, 47, 52,
    -- layer=1 filter=69 channel=119
    16, -28, -6, 7, -62, -48, 10, -38, -52,
    -- layer=1 filter=69 channel=120
    15, 0, 1, -9, 10, 22, -18, -34, -8,
    -- layer=1 filter=69 channel=121
    11, 32, 53, 38, 28, -24, 20, 55, 36,
    -- layer=1 filter=69 channel=122
    0, -2, 8, -1, 0, -5, -2, 2, -7,
    -- layer=1 filter=69 channel=123
    3, 21, 22, 8, -17, -41, 22, 28, 1,
    -- layer=1 filter=69 channel=124
    26, 21, 15, 20, 8, 28, 7, 18, 12,
    -- layer=1 filter=69 channel=125
    -1, -3, -35, -18, 27, -11, -12, 32, 43,
    -- layer=1 filter=69 channel=126
    46, 32, 19, -30, 21, 34, -19, -32, -20,
    -- layer=1 filter=69 channel=127
    -45, -13, 3, 30, -15, -44, 40, 57, 59,
    -- layer=1 filter=70 channel=0
    -1, -9, 13, 4, 4, -13, -24, -29, -18,
    -- layer=1 filter=70 channel=1
    1, -4, 0, -11, -26, -11, -20, -4, -2,
    -- layer=1 filter=70 channel=2
    -18, -9, 11, -18, -7, -9, 31, 14, 18,
    -- layer=1 filter=70 channel=3
    -1, 0, 10, -3, 16, -2, 20, 5, 15,
    -- layer=1 filter=70 channel=4
    -1, -6, 2, -8, 3, -9, -7, 5, 10,
    -- layer=1 filter=70 channel=5
    -2, -5, -4, -26, -10, -25, 3, -10, -14,
    -- layer=1 filter=70 channel=6
    -28, -27, -37, 22, 33, 23, 33, 38, 36,
    -- layer=1 filter=70 channel=7
    -22, -6, 30, -3, -41, 35, -6, -48, -15,
    -- layer=1 filter=70 channel=8
    -3, -13, 9, 11, -2, -2, 7, -5, -9,
    -- layer=1 filter=70 channel=9
    -11, -22, -37, 8, -28, -8, -2, -12, 10,
    -- layer=1 filter=70 channel=10
    -15, -11, 27, -3, -63, 8, -6, -47, -11,
    -- layer=1 filter=70 channel=11
    31, 30, 16, 14, 12, 1, -15, -12, -7,
    -- layer=1 filter=70 channel=12
    -61, -21, -42, 12, -22, -43, -63, -26, 23,
    -- layer=1 filter=70 channel=13
    -9, -18, -13, 0, 12, 24, 7, 16, 9,
    -- layer=1 filter=70 channel=14
    2, -1, 9, 0, -18, 19, 29, -8, -11,
    -- layer=1 filter=70 channel=15
    -50, -44, -21, -13, -34, -60, -3, 11, -22,
    -- layer=1 filter=70 channel=16
    9, 5, 2, 19, 7, -10, 3, 3, 14,
    -- layer=1 filter=70 channel=17
    1, 8, 21, 5, 14, 8, -36, -25, -34,
    -- layer=1 filter=70 channel=18
    25, 20, 17, 29, 25, 33, -4, 20, 6,
    -- layer=1 filter=70 channel=19
    23, 16, 0, 4, 11, 30, 35, 22, 20,
    -- layer=1 filter=70 channel=20
    -11, -26, 0, -5, 16, 16, 9, 21, 7,
    -- layer=1 filter=70 channel=21
    -63, -60, -44, -18, -27, 0, 45, 31, 25,
    -- layer=1 filter=70 channel=22
    -23, -18, 4, 32, 41, 46, 9, 30, 34,
    -- layer=1 filter=70 channel=23
    -17, 1, 11, -5, -15, -18, 7, -5, -20,
    -- layer=1 filter=70 channel=24
    -14, -41, -23, -25, -18, -7, 28, 13, 20,
    -- layer=1 filter=70 channel=25
    -18, -6, 14, -11, -50, -3, -14, -44, -2,
    -- layer=1 filter=70 channel=26
    3, 10, 4, 17, 24, 33, 1, 7, -7,
    -- layer=1 filter=70 channel=27
    20, 19, 15, 1, 7, 4, -5, -10, 4,
    -- layer=1 filter=70 channel=28
    -28, -15, 5, 1, -49, 12, -4, -56, -19,
    -- layer=1 filter=70 channel=29
    -7, -3, 7, -1, 9, 10, 23, 8, 8,
    -- layer=1 filter=70 channel=30
    35, 1, 13, 40, 11, 21, 0, 25, 10,
    -- layer=1 filter=70 channel=31
    -20, -26, -7, 8, 16, 20, 12, 18, 34,
    -- layer=1 filter=70 channel=32
    -4, 8, -14, -9, 2, 14, 1, -1, -15,
    -- layer=1 filter=70 channel=33
    0, 9, 7, 22, 30, 24, 13, 3, 12,
    -- layer=1 filter=70 channel=34
    4, -5, 0, 15, 32, 23, 24, 32, 12,
    -- layer=1 filter=70 channel=35
    -14, -18, -18, -2, -7, -10, 0, -10, -7,
    -- layer=1 filter=70 channel=36
    21, 26, 28, 12, -3, 19, -10, -26, -10,
    -- layer=1 filter=70 channel=37
    6, -2, 2, -1, -11, -4, 0, -5, 13,
    -- layer=1 filter=70 channel=38
    -20, -40, -14, -10, 9, 10, 33, 23, 41,
    -- layer=1 filter=70 channel=39
    18, 14, 10, 9, 0, -2, -1, -15, -5,
    -- layer=1 filter=70 channel=40
    1, 1, -7, 62, 52, 48, 39, 58, 47,
    -- layer=1 filter=70 channel=41
    -8, 12, -32, 3, -11, -3, -31, -6, -35,
    -- layer=1 filter=70 channel=42
    3, 8, 16, -14, 2, 8, 16, -1, -14,
    -- layer=1 filter=70 channel=43
    -3, -5, -16, 5, 5, 4, -6, 0, -2,
    -- layer=1 filter=70 channel=44
    -12, -5, 12, 4, 10, 28, 0, 2, -25,
    -- layer=1 filter=70 channel=45
    -16, -21, -22, -6, 0, -23, 6, 13, 12,
    -- layer=1 filter=70 channel=46
    3, -4, -10, 3, 27, 11, 66, 69, 47,
    -- layer=1 filter=70 channel=47
    -41, -40, -43, -17, -25, 1, 23, 24, 15,
    -- layer=1 filter=70 channel=48
    -15, -39, -8, -8, -17, -14, 8, 13, 6,
    -- layer=1 filter=70 channel=49
    -23, -30, -25, -7, -26, -5, 14, 34, 13,
    -- layer=1 filter=70 channel=50
    -2, -2, 0, 23, 13, 14, 1, 3, 20,
    -- layer=1 filter=70 channel=51
    -38, -43, -4, 7, -30, 10, 33, 26, 30,
    -- layer=1 filter=70 channel=52
    -1, 0, -8, 11, -5, 14, 4, 19, 1,
    -- layer=1 filter=70 channel=53
    -4, 5, -2, -4, -13, -10, -5, -5, 1,
    -- layer=1 filter=70 channel=54
    -14, -6, -4, -13, -42, -24, -4, -28, -17,
    -- layer=1 filter=70 channel=55
    25, 18, 24, 0, 6, 6, -31, -35, -11,
    -- layer=1 filter=70 channel=56
    -6, 3, -10, 0, -4, -8, -1, -5, -9,
    -- layer=1 filter=70 channel=57
    -6, -20, 26, 21, -20, 24, 16, -2, 12,
    -- layer=1 filter=70 channel=58
    -45, -74, 11, -22, -64, -15, 0, -41, -32,
    -- layer=1 filter=70 channel=59
    -6, 0, 4, -1, -6, -8, -4, 2, 5,
    -- layer=1 filter=70 channel=60
    1, -5, -4, -1, 4, -11, 2, 1, 12,
    -- layer=1 filter=70 channel=61
    -2, 17, 4, 0, 15, 0, 15, 5, 14,
    -- layer=1 filter=70 channel=62
    9, -8, 8, 13, 8, -5, 0, 6, 7,
    -- layer=1 filter=70 channel=63
    24, 29, 11, 10, 0, 10, -22, -13, -10,
    -- layer=1 filter=70 channel=64
    -3, -3, 2, -12, -14, 3, 6, 0, -3,
    -- layer=1 filter=70 channel=65
    -30, -20, -30, 7, -7, -3, 28, 12, 19,
    -- layer=1 filter=70 channel=66
    21, 16, 11, 4, -11, -12, -19, -17, -21,
    -- layer=1 filter=70 channel=67
    -12, -61, -67, 3, -53, -36, 5, -3, 9,
    -- layer=1 filter=70 channel=68
    -12, -13, 12, 15, -6, 35, -15, -17, -15,
    -- layer=1 filter=70 channel=69
    -2, -18, 0, -6, -11, -35, 18, 3, -12,
    -- layer=1 filter=70 channel=70
    -9, -31, -47, 39, 2, 16, 46, 59, 41,
    -- layer=1 filter=70 channel=71
    -19, -23, -12, -14, -23, -13, 16, 21, 9,
    -- layer=1 filter=70 channel=72
    -11, -3, -26, 26, 18, 25, 15, 24, 5,
    -- layer=1 filter=70 channel=73
    1, -12, -5, -9, -11, -2, -14, -6, -12,
    -- layer=1 filter=70 channel=74
    3, -10, -31, 27, 15, 16, -1, -14, 30,
    -- layer=1 filter=70 channel=75
    4, -12, -14, -1, 0, 18, 22, 16, 32,
    -- layer=1 filter=70 channel=76
    -12, 1, -15, 2, 3, 3, -29, -33, -33,
    -- layer=1 filter=70 channel=77
    -13, -24, -18, -7, -16, -21, 33, 18, 11,
    -- layer=1 filter=70 channel=78
    5, 11, 9, 6, -7, 0, -17, -18, -7,
    -- layer=1 filter=70 channel=79
    4, -2, 3, 16, 2, -16, -2, 7, 4,
    -- layer=1 filter=70 channel=80
    0, 6, -2, 0, -10, 9, 1, -2, 1,
    -- layer=1 filter=70 channel=81
    -17, -25, -22, 5, 0, -16, 32, 15, 10,
    -- layer=1 filter=70 channel=82
    -56, -51, -51, -15, -29, -31, 27, 18, 26,
    -- layer=1 filter=70 channel=83
    -4, -13, 17, -10, -26, -25, -26, -18, -35,
    -- layer=1 filter=70 channel=84
    5, 9, 11, 57, 50, 36, -6, 26, 19,
    -- layer=1 filter=70 channel=85
    -17, -36, 21, -17, -46, -6, -15, -23, -13,
    -- layer=1 filter=70 channel=86
    22, 32, 24, -4, 3, -10, -28, -39, -35,
    -- layer=1 filter=70 channel=87
    -4, -36, -37, -14, -18, -12, 20, 43, 13,
    -- layer=1 filter=70 channel=88
    -30, -42, -42, -28, -37, -32, -2, 1, -11,
    -- layer=1 filter=70 channel=89
    -39, -38, -45, -14, -3, -11, 30, 21, 16,
    -- layer=1 filter=70 channel=90
    -9, -12, 6, -3, -22, 6, -7, -22, -27,
    -- layer=1 filter=70 channel=91
    -21, -30, -16, -4, -7, 8, 11, 16, 9,
    -- layer=1 filter=70 channel=92
    -53, -31, -19, -13, -31, -17, -13, -28, -46,
    -- layer=1 filter=70 channel=93
    -22, -30, -5, -13, -22, -22, 4, -5, 5,
    -- layer=1 filter=70 channel=94
    14, 16, 20, -5, -6, 3, -22, -13, -29,
    -- layer=1 filter=70 channel=95
    27, 10, 17, 30, 28, 51, 12, 17, 37,
    -- layer=1 filter=70 channel=96
    4, 5, 10, 3, -6, 11, 5, -12, -1,
    -- layer=1 filter=70 channel=97
    0, 9, 10, 0, -2, -3, -12, -19, -24,
    -- layer=1 filter=70 channel=98
    -13, -31, 2, 21, 16, -9, 21, 9, 26,
    -- layer=1 filter=70 channel=99
    -31, -34, 21, -5, -38, -18, -17, -39, -14,
    -- layer=1 filter=70 channel=100
    14, 12, 4, 13, 9, 22, -15, -6, -7,
    -- layer=1 filter=70 channel=101
    -33, -29, -7, -6, -9, -6, 11, 31, 10,
    -- layer=1 filter=70 channel=102
    2, -8, -3, -8, -17, -11, -17, -20, -23,
    -- layer=1 filter=70 channel=103
    21, 29, 14, 29, 23, 13, -7, -9, -6,
    -- layer=1 filter=70 channel=104
    -19, 0, -3, -8, -5, -31, 8, -5, -27,
    -- layer=1 filter=70 channel=105
    12, 12, 14, 0, -12, 1, -18, -33, -25,
    -- layer=1 filter=70 channel=106
    -36, -13, -25, -1, 8, 5, 10, 30, 25,
    -- layer=1 filter=70 channel=107
    6, 3, -2, 15, 3, 12, 6, -3, 6,
    -- layer=1 filter=70 channel=108
    -20, -16, -23, -7, -15, -4, 0, -20, -33,
    -- layer=1 filter=70 channel=109
    -8, 4, -1, 10, -8, -10, 8, -1, -7,
    -- layer=1 filter=70 channel=110
    -3, -6, 4, 6, 0, 0, -2, 3, -6,
    -- layer=1 filter=70 channel=111
    14, 10, 10, 37, 7, 28, -24, 9, 8,
    -- layer=1 filter=70 channel=112
    -7, -10, 5, 27, 8, 10, -28, -9, 9,
    -- layer=1 filter=70 channel=113
    -21, -23, -5, 5, 10, 25, 24, 46, 20,
    -- layer=1 filter=70 channel=114
    20, 6, -11, -7, 5, -29, 5, -14, -23,
    -- layer=1 filter=70 channel=115
    2, 25, 37, 2, 8, -1, -20, -38, -31,
    -- layer=1 filter=70 channel=116
    4, 9, -7, 0, 9, -9, -13, 2, 6,
    -- layer=1 filter=70 channel=117
    10, 3, 35, 67, 30, 38, -30, -3, 5,
    -- layer=1 filter=70 channel=118
    30, 5, -17, 18, 24, 30, -3, 14, 26,
    -- layer=1 filter=70 channel=119
    -6, 1, -9, -13, -14, 11, -13, -14, -30,
    -- layer=1 filter=70 channel=120
    -20, -35, -26, 10, -17, -19, 28, 20, 31,
    -- layer=1 filter=70 channel=121
    15, 19, -1, -1, -18, 7, 28, 31, 15,
    -- layer=1 filter=70 channel=122
    9, 8, -9, -9, -6, 4, -8, -4, -7,
    -- layer=1 filter=70 channel=123
    8, 19, 10, 14, 6, 24, 5, 8, -5,
    -- layer=1 filter=70 channel=124
    -6, -15, -12, -17, -13, -15, -2, -18, -6,
    -- layer=1 filter=70 channel=125
    -18, -26, -40, 14, -5, -3, 48, 51, 23,
    -- layer=1 filter=70 channel=126
    10, -20, 11, 24, 10, 13, 17, 29, 39,
    -- layer=1 filter=70 channel=127
    31, 13, 20, 45, 36, 38, 8, 16, 26,
    -- layer=1 filter=71 channel=0
    7, 6, 3, 6, 8, -4, -11, 2, 3,
    -- layer=1 filter=71 channel=1
    -4, -4, 8, -5, -2, 1, -9, -12, 4,
    -- layer=1 filter=71 channel=2
    9, -10, -1, 3, -3, 1, 4, -2, -5,
    -- layer=1 filter=71 channel=3
    8, -3, 5, 10, -6, 4, 0, -10, 9,
    -- layer=1 filter=71 channel=4
    -2, -11, -5, 8, 7, 4, -11, 7, 4,
    -- layer=1 filter=71 channel=5
    -3, -3, 0, -8, -6, 4, 0, 1, -11,
    -- layer=1 filter=71 channel=6
    6, 2, 6, 2, -3, -11, -11, 0, 1,
    -- layer=1 filter=71 channel=7
    -13, -4, 0, -2, 2, -5, -7, -17, -5,
    -- layer=1 filter=71 channel=8
    0, -9, 3, -5, -9, -7, 0, 3, -12,
    -- layer=1 filter=71 channel=9
    0, 1, 0, 0, -7, 8, -11, -6, 3,
    -- layer=1 filter=71 channel=10
    -1, 8, -9, -7, -6, -8, -10, -4, -10,
    -- layer=1 filter=71 channel=11
    1, -6, 8, -11, -2, 6, -10, 9, 9,
    -- layer=1 filter=71 channel=12
    11, -6, 9, -5, 5, -1, -6, 7, 2,
    -- layer=1 filter=71 channel=13
    7, 6, -1, 6, -10, -11, -9, 4, -1,
    -- layer=1 filter=71 channel=14
    -10, 4, 3, -8, -11, 9, 8, 2, 0,
    -- layer=1 filter=71 channel=15
    1, 0, 6, -12, -3, -4, 7, 3, -12,
    -- layer=1 filter=71 channel=16
    3, -11, -8, -11, -9, -7, -5, -5, -3,
    -- layer=1 filter=71 channel=17
    4, 3, 6, -10, -5, -4, -1, -8, -5,
    -- layer=1 filter=71 channel=18
    -9, -5, -7, -6, 0, 5, -5, -9, 2,
    -- layer=1 filter=71 channel=19
    -5, -7, -7, -1, 5, 0, -2, 8, -4,
    -- layer=1 filter=71 channel=20
    -10, 6, -2, 3, -1, -3, -1, -5, 2,
    -- layer=1 filter=71 channel=21
    0, 4, 4, 6, -5, -2, -1, 5, 2,
    -- layer=1 filter=71 channel=22
    3, 7, 5, 0, 1, 8, 8, 0, 8,
    -- layer=1 filter=71 channel=23
    1, -5, 4, 2, 2, -13, -8, -2, -5,
    -- layer=1 filter=71 channel=24
    6, -5, 4, -13, 3, 5, -1, 3, -11,
    -- layer=1 filter=71 channel=25
    -8, -8, 3, -2, 0, 9, -7, 4, 0,
    -- layer=1 filter=71 channel=26
    -6, 4, 4, -12, -11, 0, 8, 4, 6,
    -- layer=1 filter=71 channel=27
    -9, -10, -4, 1, -7, 0, -3, 10, 5,
    -- layer=1 filter=71 channel=28
    4, 2, 3, 6, -8, -5, -11, -10, 3,
    -- layer=1 filter=71 channel=29
    3, 5, 1, -7, -14, 0, 3, -8, 8,
    -- layer=1 filter=71 channel=30
    -9, 7, -10, 0, -8, -10, -3, -7, -11,
    -- layer=1 filter=71 channel=31
    2, -7, -7, 4, 0, 3, -8, -3, 6,
    -- layer=1 filter=71 channel=32
    -5, 4, 3, 4, -4, 1, -6, -9, -1,
    -- layer=1 filter=71 channel=33
    2, 7, 8, 4, 9, 3, 5, -1, -1,
    -- layer=1 filter=71 channel=34
    -12, -3, 3, 5, 6, -7, 3, -10, -8,
    -- layer=1 filter=71 channel=35
    -9, 4, -1, 6, 7, -9, -1, -4, -6,
    -- layer=1 filter=71 channel=36
    -8, 7, -3, 0, 2, 7, 2, 0, -5,
    -- layer=1 filter=71 channel=37
    0, -6, 7, -3, 7, -2, 7, -2, -1,
    -- layer=1 filter=71 channel=38
    -6, -10, -11, -10, 1, -12, -4, 0, 1,
    -- layer=1 filter=71 channel=39
    -11, -3, 8, 6, 1, -4, -6, -10, -4,
    -- layer=1 filter=71 channel=40
    -5, 7, -2, -10, -9, -2, -6, 7, -6,
    -- layer=1 filter=71 channel=41
    -6, -9, 3, 6, -11, 5, 4, -10, 0,
    -- layer=1 filter=71 channel=42
    8, 6, 10, 6, -7, 11, -4, 0, -6,
    -- layer=1 filter=71 channel=43
    -2, -8, 7, 1, 10, 7, -9, -11, -8,
    -- layer=1 filter=71 channel=44
    2, -9, -6, -4, -9, -10, -4, -2, -9,
    -- layer=1 filter=71 channel=45
    5, 6, 7, 2, -10, 1, -7, 0, -4,
    -- layer=1 filter=71 channel=46
    -11, -9, -3, -4, -5, 4, -9, 7, -2,
    -- layer=1 filter=71 channel=47
    6, -4, -5, 6, -1, 1, 1, -9, -6,
    -- layer=1 filter=71 channel=48
    0, 1, 4, 4, -10, 0, -12, -11, -11,
    -- layer=1 filter=71 channel=49
    -11, 1, 5, -10, -2, 6, -7, 8, -4,
    -- layer=1 filter=71 channel=50
    2, 5, -1, 7, 6, -11, -8, -10, 9,
    -- layer=1 filter=71 channel=51
    -7, -5, -2, -4, -3, -1, 0, -4, 0,
    -- layer=1 filter=71 channel=52
    2, -7, 0, -8, -3, 6, 9, 4, 0,
    -- layer=1 filter=71 channel=53
    -2, 1, -7, 0, -7, -8, -10, -4, -7,
    -- layer=1 filter=71 channel=54
    -4, -7, -3, -9, 0, 0, 7, -11, -11,
    -- layer=1 filter=71 channel=55
    -5, -5, -6, 4, 1, -5, -1, 4, -9,
    -- layer=1 filter=71 channel=56
    1, -1, -9, -6, -5, -9, -9, -2, -7,
    -- layer=1 filter=71 channel=57
    -5, -3, 5, -3, -6, 1, -10, -2, 0,
    -- layer=1 filter=71 channel=58
    7, -2, -3, 8, 5, -4, -3, 3, 8,
    -- layer=1 filter=71 channel=59
    3, 0, -6, -5, -10, 7, 0, -9, -4,
    -- layer=1 filter=71 channel=60
    -1, 7, -11, -4, 0, -1, 4, -7, 0,
    -- layer=1 filter=71 channel=61
    5, -3, 10, -6, 9, -2, 6, -3, -5,
    -- layer=1 filter=71 channel=62
    -10, -10, -1, -1, 4, -11, -3, 2, -6,
    -- layer=1 filter=71 channel=63
    0, -12, 0, -11, 3, -7, 2, -7, -7,
    -- layer=1 filter=71 channel=64
    1, 2, 6, 8, 3, -9, 2, 5, -4,
    -- layer=1 filter=71 channel=65
    -9, 0, -12, -11, 8, 5, -7, 0, -12,
    -- layer=1 filter=71 channel=66
    0, 7, 1, 4, -10, -1, -6, 3, -10,
    -- layer=1 filter=71 channel=67
    9, -5, -4, -6, 2, 6, 1, -7, 0,
    -- layer=1 filter=71 channel=68
    -8, -2, -12, 7, -1, 2, -2, -11, 4,
    -- layer=1 filter=71 channel=69
    -4, -5, 4, -8, -13, -11, -7, 7, -8,
    -- layer=1 filter=71 channel=70
    0, 0, 2, -4, 9, -6, 8, 2, -4,
    -- layer=1 filter=71 channel=71
    -12, 0, 6, -3, -1, -11, 0, 5, 0,
    -- layer=1 filter=71 channel=72
    -6, 0, -4, 0, -10, 4, -4, -9, -5,
    -- layer=1 filter=71 channel=73
    6, 7, -7, 0, 6, -10, 8, -11, 2,
    -- layer=1 filter=71 channel=74
    -11, -3, -6, -10, 1, -9, 7, -2, -7,
    -- layer=1 filter=71 channel=75
    -8, -2, -8, 6, 5, -3, -10, 1, -1,
    -- layer=1 filter=71 channel=76
    -5, -8, -10, -12, 0, -10, -10, -8, 7,
    -- layer=1 filter=71 channel=77
    -1, 8, -4, -5, -2, 7, 1, -4, 3,
    -- layer=1 filter=71 channel=78
    0, 0, 5, 4, 0, 8, -10, 1, 6,
    -- layer=1 filter=71 channel=79
    -4, -2, -6, -7, 5, 0, 7, 2, -8,
    -- layer=1 filter=71 channel=80
    -10, 5, 3, -8, -6, -7, -8, 7, 8,
    -- layer=1 filter=71 channel=81
    8, 7, -11, 2, -2, -9, -1, 1, 5,
    -- layer=1 filter=71 channel=82
    8, 5, -2, 8, -2, -4, -9, -5, 1,
    -- layer=1 filter=71 channel=83
    2, 8, -7, 2, 2, -4, 6, 4, 5,
    -- layer=1 filter=71 channel=84
    -6, 3, 2, -1, 3, 1, 6, -4, -12,
    -- layer=1 filter=71 channel=85
    7, -13, -13, -11, -10, 7, 5, 4, 0,
    -- layer=1 filter=71 channel=86
    7, 3, -6, 6, 0, 0, 2, -3, -9,
    -- layer=1 filter=71 channel=87
    8, -10, 2, 4, 5, -2, -3, -9, 3,
    -- layer=1 filter=71 channel=88
    -1, -8, -9, -7, -5, 1, -7, -4, 9,
    -- layer=1 filter=71 channel=89
    -3, -8, -7, -10, 3, -8, -11, 4, 6,
    -- layer=1 filter=71 channel=90
    -9, 4, -8, -7, -8, 6, 1, -5, -8,
    -- layer=1 filter=71 channel=91
    6, -6, -11, 8, -7, 1, -11, -8, 5,
    -- layer=1 filter=71 channel=92
    -6, 0, 8, 0, -10, 1, 4, 8, -1,
    -- layer=1 filter=71 channel=93
    -1, -2, 3, -2, -4, -7, 0, 0, -13,
    -- layer=1 filter=71 channel=94
    -5, -9, -6, -1, -2, 0, 2, 0, 4,
    -- layer=1 filter=71 channel=95
    0, 1, 2, -7, 5, 5, -8, -9, 6,
    -- layer=1 filter=71 channel=96
    -5, -5, 3, -8, -1, 0, -6, 7, 6,
    -- layer=1 filter=71 channel=97
    6, -1, -2, 6, 0, -5, -3, -10, -10,
    -- layer=1 filter=71 channel=98
    -6, 4, 8, -2, -9, 1, -10, 4, -6,
    -- layer=1 filter=71 channel=99
    -2, -3, 1, -11, 4, 7, 2, 0, 2,
    -- layer=1 filter=71 channel=100
    2, -3, 1, 3, 3, 1, -8, -1, 8,
    -- layer=1 filter=71 channel=101
    0, -6, 4, -2, -5, 2, 9, 7, -2,
    -- layer=1 filter=71 channel=102
    2, 1, 6, 1, -5, -3, 3, -3, -1,
    -- layer=1 filter=71 channel=103
    -4, -5, 3, 7, 7, -2, 0, -9, -4,
    -- layer=1 filter=71 channel=104
    3, -4, -4, 7, -1, 4, -10, 7, -6,
    -- layer=1 filter=71 channel=105
    -1, 5, -8, -1, -7, 4, -12, 4, 4,
    -- layer=1 filter=71 channel=106
    -1, 0, 1, 1, 4, 6, 8, -10, -6,
    -- layer=1 filter=71 channel=107
    -1, -4, -7, -3, -9, -6, -2, 1, 9,
    -- layer=1 filter=71 channel=108
    -6, -8, 3, -6, 6, 0, 3, 8, -4,
    -- layer=1 filter=71 channel=109
    -4, 9, -6, -7, -3, 8, 5, 0, 2,
    -- layer=1 filter=71 channel=110
    5, -9, -4, -10, 1, 6, -1, -5, 5,
    -- layer=1 filter=71 channel=111
    -4, -9, -13, 3, -3, -8, -2, 4, 0,
    -- layer=1 filter=71 channel=112
    0, 4, -3, 5, -6, -8, -1, -4, -2,
    -- layer=1 filter=71 channel=113
    4, -4, 4, 4, 6, 2, 2, -1, 2,
    -- layer=1 filter=71 channel=114
    -4, 10, 7, 8, -3, 3, 9, 1, 3,
    -- layer=1 filter=71 channel=115
    -7, 5, 2, 7, -8, -11, -6, 1, -7,
    -- layer=1 filter=71 channel=116
    1, -1, -2, -10, 0, 7, -6, -4, 6,
    -- layer=1 filter=71 channel=117
    -12, -10, -4, 7, -11, 2, 3, -2, -2,
    -- layer=1 filter=71 channel=118
    -7, -3, -9, -1, -1, -4, -7, -1, -7,
    -- layer=1 filter=71 channel=119
    0, 7, -13, 1, -9, -4, 4, -5, -8,
    -- layer=1 filter=71 channel=120
    8, -3, -4, -7, 5, 5, -1, -1, -1,
    -- layer=1 filter=71 channel=121
    -10, -9, -11, 0, -7, -9, -1, 0, 5,
    -- layer=1 filter=71 channel=122
    4, -1, 7, -10, 6, -4, -3, -5, -8,
    -- layer=1 filter=71 channel=123
    -11, 5, 2, -8, -12, -1, -8, -8, 5,
    -- layer=1 filter=71 channel=124
    4, -8, -7, -11, 1, -5, 2, 2, 0,
    -- layer=1 filter=71 channel=125
    -4, 5, 4, 0, 5, -10, 9, -7, -8,
    -- layer=1 filter=71 channel=126
    2, -13, -5, -10, -6, -5, 7, -1, 3,
    -- layer=1 filter=71 channel=127
    -5, -10, 3, -1, 7, -5, -10, 0, 0,
    -- layer=1 filter=72 channel=0
    -12, -15, 9, -15, -6, -6, 7, 3, -8,
    -- layer=1 filter=72 channel=1
    -1, -9, -27, 13, -8, 16, -4, -11, -11,
    -- layer=1 filter=72 channel=2
    8, 5, 7, -1, 1, 17, -9, -8, -7,
    -- layer=1 filter=72 channel=3
    0, -16, 1, 1, 4, 4, 5, -8, -2,
    -- layer=1 filter=72 channel=4
    -6, 0, -2, -11, -3, -14, -7, -8, 4,
    -- layer=1 filter=72 channel=5
    3, 9, -8, 2, -4, 17, 18, 11, 0,
    -- layer=1 filter=72 channel=6
    -23, -13, 3, -40, -24, -44, -52, -42, -17,
    -- layer=1 filter=72 channel=7
    -48, -74, -67, -85, -120, -75, -81, -75, -59,
    -- layer=1 filter=72 channel=8
    10, -8, -22, 11, 14, 31, 8, 3, 24,
    -- layer=1 filter=72 channel=9
    -25, -22, -65, -42, -28, -20, -23, -46, -1,
    -- layer=1 filter=72 channel=10
    -41, -45, -39, -30, -80, -38, -38, -56, -58,
    -- layer=1 filter=72 channel=11
    -19, 4, 2, 5, -3, 4, -10, -15, -4,
    -- layer=1 filter=72 channel=12
    -70, -57, -38, -10, -36, -18, 11, -12, 10,
    -- layer=1 filter=72 channel=13
    1, 4, 5, 1, 0, -5, 9, 7, 12,
    -- layer=1 filter=72 channel=14
    4, -26, -12, -7, -50, 0, -2, -6, -56,
    -- layer=1 filter=72 channel=15
    13, -8, 20, -10, -21, -12, -27, -37, -41,
    -- layer=1 filter=72 channel=16
    16, 4, 1, 22, 23, 10, 25, 23, 15,
    -- layer=1 filter=72 channel=17
    -23, -19, -22, -13, -4, -15, -12, 0, -11,
    -- layer=1 filter=72 channel=18
    12, 9, 25, 12, 17, 22, -10, -24, -13,
    -- layer=1 filter=72 channel=19
    13, 7, 39, 7, 3, -14, -4, -27, 5,
    -- layer=1 filter=72 channel=20
    -9, 2, -4, -6, 2, 5, 9, 18, 0,
    -- layer=1 filter=72 channel=21
    -9, 5, -19, 9, 15, 4, -2, 15, -1,
    -- layer=1 filter=72 channel=22
    -1, -5, 5, 7, -3, 4, 4, -5, -5,
    -- layer=1 filter=72 channel=23
    -23, -44, -48, -49, -33, -55, -40, -48, -24,
    -- layer=1 filter=72 channel=24
    -3, 3, -7, 14, 8, 19, 13, 13, 30,
    -- layer=1 filter=72 channel=25
    -25, -35, -33, -12, -29, -41, -17, -15, 0,
    -- layer=1 filter=72 channel=26
    8, -8, 0, 10, -36, -3, -1, 9, -9,
    -- layer=1 filter=72 channel=27
    -31, -29, -33, -13, -6, -5, 9, 10, 8,
    -- layer=1 filter=72 channel=28
    -31, -33, -35, -19, -40, -25, -4, -28, -5,
    -- layer=1 filter=72 channel=29
    -41, -31, -46, -23, -28, -21, -19, -26, -12,
    -- layer=1 filter=72 channel=30
    37, 15, 15, 5, 10, 8, 31, -10, 7,
    -- layer=1 filter=72 channel=31
    0, -18, 3, 16, 21, 8, 15, 15, 23,
    -- layer=1 filter=72 channel=32
    10, -33, -29, -28, -79, -19, -20, -48, -41,
    -- layer=1 filter=72 channel=33
    -22, -12, 0, -8, -2, -7, 4, -8, -23,
    -- layer=1 filter=72 channel=34
    -36, -31, -33, -30, -18, -31, -10, -22, -18,
    -- layer=1 filter=72 channel=35
    3, 4, -7, -12, -8, -11, 1, -4, 1,
    -- layer=1 filter=72 channel=36
    0, 2, 6, 2, -2, 4, -10, -1, -8,
    -- layer=1 filter=72 channel=37
    17, 8, 10, -11, 4, 13, 13, -1, 4,
    -- layer=1 filter=72 channel=38
    5, 9, 9, 5, 0, 8, 8, 4, 10,
    -- layer=1 filter=72 channel=39
    -22, -12, -11, -7, -3, -5, 4, 6, 19,
    -- layer=1 filter=72 channel=40
    13, -3, 15, -40, -7, -15, 17, -15, -6,
    -- layer=1 filter=72 channel=41
    1, -27, -31, -19, -32, -23, -32, -59, 14,
    -- layer=1 filter=72 channel=42
    4, -1, 10, 15, 1, 20, -23, -11, -16,
    -- layer=1 filter=72 channel=43
    -16, -5, -34, 25, 2, 19, 5, -6, 5,
    -- layer=1 filter=72 channel=44
    -24, -72, -64, -19, -97, -8, -24, -41, -42,
    -- layer=1 filter=72 channel=45
    -7, -5, 2, 12, 1, 16, -5, -17, -14,
    -- layer=1 filter=72 channel=46
    35, 29, 32, 18, -5, -22, 11, -7, -11,
    -- layer=1 filter=72 channel=47
    24, -39, -13, -34, -15, -30, -14, -29, -18,
    -- layer=1 filter=72 channel=48
    4, 1, -2, 8, 9, -8, 4, 7, 5,
    -- layer=1 filter=72 channel=49
    28, 10, 18, 16, 2, 16, 7, 9, 15,
    -- layer=1 filter=72 channel=50
    -4, -11, -15, -7, -3, -28, 10, 13, -2,
    -- layer=1 filter=72 channel=51
    -4, 2, 3, 1, 6, -1, 5, 2, -4,
    -- layer=1 filter=72 channel=52
    0, 17, 23, 26, 22, 29, 2, 8, 2,
    -- layer=1 filter=72 channel=53
    -3, -5, 0, -6, -10, 7, -2, -4, -3,
    -- layer=1 filter=72 channel=54
    -20, -26, -34, -4, -20, -29, -1, -11, 3,
    -- layer=1 filter=72 channel=55
    -3, 12, 4, 2, 11, 7, 5, 8, 24,
    -- layer=1 filter=72 channel=56
    9, -8, 7, -8, -7, -9, 2, -8, -7,
    -- layer=1 filter=72 channel=57
    -1, -26, -3, -12, -39, -17, 12, -21, -13,
    -- layer=1 filter=72 channel=58
    -54, -98, -63, -86, -62, -67, -66, -71, -51,
    -- layer=1 filter=72 channel=59
    -7, -11, 1, 8, 0, -10, 5, 5, 1,
    -- layer=1 filter=72 channel=60
    -11, -3, -10, -13, -6, -21, -7, -7, -6,
    -- layer=1 filter=72 channel=61
    3, -1, 3, 3, -2, -1, 5, -4, 1,
    -- layer=1 filter=72 channel=62
    9, -13, -21, 10, 7, 17, 17, -1, 4,
    -- layer=1 filter=72 channel=63
    -11, 8, -1, 4, 13, -4, 7, 7, 2,
    -- layer=1 filter=72 channel=64
    -3, -1, 0, -12, -17, -7, 0, 0, -1,
    -- layer=1 filter=72 channel=65
    -1, -12, -4, -15, 5, 0, -5, -5, -7,
    -- layer=1 filter=72 channel=66
    -5, 2, 0, -4, -5, 13, 2, 3, 2,
    -- layer=1 filter=72 channel=67
    -3, -6, -14, -27, -26, -38, -41, -41, -44,
    -- layer=1 filter=72 channel=68
    -47, -77, -69, -70, -106, -60, -60, -51, -47,
    -- layer=1 filter=72 channel=69
    18, 7, 11, 13, -5, 24, 28, 8, -2,
    -- layer=1 filter=72 channel=70
    8, -14, 25, -20, -34, -5, -35, -33, -32,
    -- layer=1 filter=72 channel=71
    -5, -11, -15, 20, 6, 14, 11, 0, -1,
    -- layer=1 filter=72 channel=72
    18, 6, 20, 24, 32, 5, -7, -38, 17,
    -- layer=1 filter=72 channel=73
    6, -5, 2, -9, 3, 0, 12, -5, 0,
    -- layer=1 filter=72 channel=74
    -14, -4, -13, -14, -5, -3, -21, -12, -9,
    -- layer=1 filter=72 channel=75
    6, -17, -5, 21, 2, 34, 22, 12, 5,
    -- layer=1 filter=72 channel=76
    -8, -11, -18, -5, -14, -19, -12, -19, -8,
    -- layer=1 filter=72 channel=77
    -5, -14, -9, -4, 0, 16, -7, -6, 4,
    -- layer=1 filter=72 channel=78
    -8, -19, 1, 0, -6, -17, -7, -3, 0,
    -- layer=1 filter=72 channel=79
    11, -13, 5, 16, 10, 7, 13, 14, 2,
    -- layer=1 filter=72 channel=80
    -6, -8, -3, -11, 1, -19, -26, -13, -9,
    -- layer=1 filter=72 channel=81
    -5, -26, -30, 0, 1, 1, 9, -4, 8,
    -- layer=1 filter=72 channel=82
    5, -7, 0, 16, 1, 16, 1, 14, 0,
    -- layer=1 filter=72 channel=83
    -1, -24, -4, 15, -12, 4, -15, -19, -16,
    -- layer=1 filter=72 channel=84
    3, 16, 8, 5, 9, 8, -22, 0, -2,
    -- layer=1 filter=72 channel=85
    -2, -23, -32, -48, -33, -27, -28, -34, -3,
    -- layer=1 filter=72 channel=86
    7, 4, 0, 3, -7, -7, 0, -1, 0,
    -- layer=1 filter=72 channel=87
    22, 7, 12, -11, 16, -28, 7, -20, 8,
    -- layer=1 filter=72 channel=88
    -9, 7, -9, -11, 12, 0, -7, -3, 7,
    -- layer=1 filter=72 channel=89
    5, 8, -8, 2, 11, 4, -4, 0, -1,
    -- layer=1 filter=72 channel=90
    -48, -101, -72, -16, -93, -21, -42, -41, -62,
    -- layer=1 filter=72 channel=91
    21, 8, 17, 14, 4, 2, 18, 11, 16,
    -- layer=1 filter=72 channel=92
    -67, -44, -7, -85, -65, -15, -44, -59, -20,
    -- layer=1 filter=72 channel=93
    3, 6, 6, 16, 10, 18, 20, 23, 26,
    -- layer=1 filter=72 channel=94
    -1, -7, 2, -8, -13, -7, -12, -20, -10,
    -- layer=1 filter=72 channel=95
    20, 9, 23, -3, 0, 27, -5, -3, -11,
    -- layer=1 filter=72 channel=96
    -14, -3, -8, -3, -3, 0, -17, -2, 7,
    -- layer=1 filter=72 channel=97
    0, -6, -4, -2, 8, 8, 8, 0, 5,
    -- layer=1 filter=72 channel=98
    19, 2, 1, 25, 24, 13, 0, 1, 0,
    -- layer=1 filter=72 channel=99
    -49, -5, -10, -31, -21, -37, 16, -42, -43,
    -- layer=1 filter=72 channel=100
    -2, -14, -2, -5, 6, 3, 8, 6, -8,
    -- layer=1 filter=72 channel=101
    13, 15, 0, 4, 15, 11, 18, 3, 12,
    -- layer=1 filter=72 channel=102
    -6, -11, -1, -22, -28, -26, -8, -14, -29,
    -- layer=1 filter=72 channel=103
    -21, -14, -10, -8, -5, 8, -18, -14, -10,
    -- layer=1 filter=72 channel=104
    29, 7, 4, -18, 10, 2, -9, -30, -11,
    -- layer=1 filter=72 channel=105
    -9, 6, 9, 8, 2, 11, 0, 6, -2,
    -- layer=1 filter=72 channel=106
    29, 7, 10, 0, 4, 8, 8, 6, 11,
    -- layer=1 filter=72 channel=107
    0, 0, 0, 18, 2, 15, 0, -5, 8,
    -- layer=1 filter=72 channel=108
    -6, -89, -44, -16, -73, -33, -15, -59, -29,
    -- layer=1 filter=72 channel=109
    -6, -3, -10, 2, 2, -3, 1, -9, -4,
    -- layer=1 filter=72 channel=110
    2, 0, -6, 3, -14, -4, -10, -9, 0,
    -- layer=1 filter=72 channel=111
    5, 10, 4, 2, 8, 16, 19, 0, -14,
    -- layer=1 filter=72 channel=112
    -6, 13, 15, 15, 0, 12, -29, -12, -20,
    -- layer=1 filter=72 channel=113
    -8, -11, 16, 7, 12, 2, 1, 10, 15,
    -- layer=1 filter=72 channel=114
    0, -2, -10, 2, -17, -12, 9, -14, -9,
    -- layer=1 filter=72 channel=115
    -7, -9, 3, -10, 0, -5, -4, -8, 2,
    -- layer=1 filter=72 channel=116
    -10, -1, -3, -2, -6, 6, 7, -7, 4,
    -- layer=1 filter=72 channel=117
    6, 20, 42, 44, 28, 10, 27, -15, -36,
    -- layer=1 filter=72 channel=118
    33, 29, 23, 17, 1, 4, 24, -8, 21,
    -- layer=1 filter=72 channel=119
    -2, -74, -63, -45, -88, -59, -37, -80, -34,
    -- layer=1 filter=72 channel=120
    2, 1, -12, 9, 15, 10, -1, 16, 14,
    -- layer=1 filter=72 channel=121
    20, 18, 0, 17, 8, 5, 34, 4, 3,
    -- layer=1 filter=72 channel=122
    7, 1, -7, 4, -7, 1, 7, 4, -7,
    -- layer=1 filter=72 channel=123
    10, -3, -7, -7, 8, 18, 23, 7, 5,
    -- layer=1 filter=72 channel=124
    -11, -17, -16, -15, -25, -13, -10, -8, -13,
    -- layer=1 filter=72 channel=125
    15, 4, 13, -26, -20, -33, -7, -45, -33,
    -- layer=1 filter=72 channel=126
    0, -12, -21, 37, 0, 14, -4, -7, 3,
    -- layer=1 filter=72 channel=127
    45, 33, 34, 19, 47, 28, 18, 13, 4,
    -- layer=1 filter=73 channel=0
    -7, -7, 4, -1, -10, 3, 0, 6, 0,
    -- layer=1 filter=73 channel=1
    6, 2, 2, 2, 6, -9, -11, -5, 5,
    -- layer=1 filter=73 channel=2
    -4, 0, -5, -13, -10, -8, 0, -15, -15,
    -- layer=1 filter=73 channel=3
    -8, -3, 0, -7, -6, 5, -3, 4, 0,
    -- layer=1 filter=73 channel=4
    2, -9, 8, -6, 2, -3, -10, -6, 8,
    -- layer=1 filter=73 channel=5
    7, -8, 1, -3, -10, 12, -5, 8, 1,
    -- layer=1 filter=73 channel=6
    6, 2, -15, 5, -6, 0, -7, 3, -3,
    -- layer=1 filter=73 channel=7
    -8, -9, -9, 1, -9, 0, 0, 1, -12,
    -- layer=1 filter=73 channel=8
    -3, 5, 6, -6, -9, -4, -7, 6, -12,
    -- layer=1 filter=73 channel=9
    -8, 4, 0, -7, -8, -3, -11, -8, -4,
    -- layer=1 filter=73 channel=10
    3, -7, 1, -5, -17, -14, -13, 2, -11,
    -- layer=1 filter=73 channel=11
    -3, 6, 7, 8, 6, 6, 3, -9, -4,
    -- layer=1 filter=73 channel=12
    2, 7, -9, 0, -6, -10, 5, 10, -1,
    -- layer=1 filter=73 channel=13
    -12, 0, -2, -6, -10, 4, 2, -6, -3,
    -- layer=1 filter=73 channel=14
    0, 7, -10, -5, -13, -8, -2, 1, -2,
    -- layer=1 filter=73 channel=15
    -5, 3, -1, -1, 6, -9, 6, -4, 2,
    -- layer=1 filter=73 channel=16
    -3, 2, -6, -8, -10, -4, -1, 6, 7,
    -- layer=1 filter=73 channel=17
    -6, 2, 2, 4, -3, 1, 5, -3, -2,
    -- layer=1 filter=73 channel=18
    -4, -8, -10, -3, 4, 0, -3, 4, -3,
    -- layer=1 filter=73 channel=19
    5, 2, 1, -2, 0, -3, 4, 7, -3,
    -- layer=1 filter=73 channel=20
    8, 6, 2, -7, 3, -10, -3, -5, 4,
    -- layer=1 filter=73 channel=21
    0, 0, -4, -2, 4, -11, -6, 2, -11,
    -- layer=1 filter=73 channel=22
    -10, 0, -3, 5, 3, 1, -3, -7, 0,
    -- layer=1 filter=73 channel=23
    -3, 5, -3, -6, 6, 2, -10, 6, 0,
    -- layer=1 filter=73 channel=24
    -5, 7, -11, 0, -10, -11, 7, -6, -7,
    -- layer=1 filter=73 channel=25
    -11, -1, -3, -10, -9, -2, -1, 2, -12,
    -- layer=1 filter=73 channel=26
    1, -8, -4, 0, 1, -11, 0, -5, 4,
    -- layer=1 filter=73 channel=27
    -4, 1, 5, -1, 8, -1, 8, -6, 1,
    -- layer=1 filter=73 channel=28
    6, -7, -9, -9, -5, -1, 5, -9, 3,
    -- layer=1 filter=73 channel=29
    8, -6, -6, -9, -10, 5, -2, -6, -4,
    -- layer=1 filter=73 channel=30
    -12, 1, -1, -10, -7, -6, 2, 0, -11,
    -- layer=1 filter=73 channel=31
    -2, 2, -3, -11, 1, -1, -7, 4, -5,
    -- layer=1 filter=73 channel=32
    5, 4, 0, 8, 7, -9, -10, -11, -8,
    -- layer=1 filter=73 channel=33
    -6, -4, -3, 9, 8, 5, 9, -3, 11,
    -- layer=1 filter=73 channel=34
    7, 9, 0, -3, -2, 6, 3, -8, -2,
    -- layer=1 filter=73 channel=35
    -6, -11, 3, -7, -4, 0, 4, -6, 4,
    -- layer=1 filter=73 channel=36
    -8, -9, -1, -2, -10, 0, 0, -5, -5,
    -- layer=1 filter=73 channel=37
    -9, 2, 1, -7, -7, 0, 0, 8, 0,
    -- layer=1 filter=73 channel=38
    5, 5, -14, -5, -2, -5, -1, 0, -4,
    -- layer=1 filter=73 channel=39
    -11, -11, 3, 2, 6, 5, -3, 2, -7,
    -- layer=1 filter=73 channel=40
    6, -5, -7, 7, 0, 0, 1, -9, -11,
    -- layer=1 filter=73 channel=41
    -1, -5, -7, 1, 8, -4, -7, -9, -2,
    -- layer=1 filter=73 channel=42
    0, -5, -4, -10, -9, -1, -9, -17, -8,
    -- layer=1 filter=73 channel=43
    0, 8, -10, 0, 0, -7, 0, -7, -10,
    -- layer=1 filter=73 channel=44
    -1, 5, 3, -8, -1, -2, -7, 0, -5,
    -- layer=1 filter=73 channel=45
    -1, -3, -7, 0, -5, -10, 1, -6, -3,
    -- layer=1 filter=73 channel=46
    -2, 3, -1, -8, -7, 1, -1, -8, 0,
    -- layer=1 filter=73 channel=47
    -9, 8, -2, -8, -7, -5, -4, -8, -11,
    -- layer=1 filter=73 channel=48
    -5, -11, -6, -2, -3, -5, 4, -8, 4,
    -- layer=1 filter=73 channel=49
    3, -8, 4, 0, -1, -9, -8, -11, -2,
    -- layer=1 filter=73 channel=50
    7, -6, 2, -2, -8, -5, -11, 1, 2,
    -- layer=1 filter=73 channel=51
    -6, -3, -10, 6, -7, 4, 4, 2, 5,
    -- layer=1 filter=73 channel=52
    0, 5, -5, 5, -3, -7, 9, -7, -10,
    -- layer=1 filter=73 channel=53
    0, 0, -11, 0, -1, -10, -6, -8, -10,
    -- layer=1 filter=73 channel=54
    -7, -7, -3, 6, 2, -3, -6, -3, -1,
    -- layer=1 filter=73 channel=55
    -5, 0, -5, -16, -8, 0, -16, -2, -10,
    -- layer=1 filter=73 channel=56
    -2, 3, -5, -8, 1, -11, 0, 0, 1,
    -- layer=1 filter=73 channel=57
    -10, -2, 0, -7, 0, 2, 2, -1, 4,
    -- layer=1 filter=73 channel=58
    -3, 5, -12, -1, -9, -1, -7, -3, -8,
    -- layer=1 filter=73 channel=59
    -1, 8, 3, -8, -5, 3, 7, -5, -6,
    -- layer=1 filter=73 channel=60
    -1, 1, -7, 6, -1, -3, -4, 8, 8,
    -- layer=1 filter=73 channel=61
    2, -2, 9, 1, 10, 4, 1, -8, -5,
    -- layer=1 filter=73 channel=62
    5, -8, -5, 2, -8, 9, -5, -7, -8,
    -- layer=1 filter=73 channel=63
    0, -1, 1, 1, 5, 9, 2, 0, -10,
    -- layer=1 filter=73 channel=64
    -1, -3, -1, 0, -2, -7, -11, -8, 7,
    -- layer=1 filter=73 channel=65
    3, -11, -1, -4, 0, -11, 6, -7, -5,
    -- layer=1 filter=73 channel=66
    -11, -4, -8, -3, 8, -4, 0, -7, -9,
    -- layer=1 filter=73 channel=67
    -10, 3, 4, 9, 0, 3, 2, 0, -3,
    -- layer=1 filter=73 channel=68
    -7, 4, 4, -1, 7, 0, -4, -5, -1,
    -- layer=1 filter=73 channel=69
    -3, 0, 5, -13, 5, -6, -8, -3, -7,
    -- layer=1 filter=73 channel=70
    -3, 1, -9, -6, 2, -3, -4, -12, 3,
    -- layer=1 filter=73 channel=71
    3, -9, -5, -5, 3, -6, -7, -11, 3,
    -- layer=1 filter=73 channel=72
    -9, 1, -3, 3, 4, -9, 5, -4, 0,
    -- layer=1 filter=73 channel=73
    -10, 1, 8, -2, 8, -6, 0, -2, 0,
    -- layer=1 filter=73 channel=74
    4, -6, 7, -3, 6, 0, 0, 0, 1,
    -- layer=1 filter=73 channel=75
    0, 1, 0, 2, -14, 2, -6, -3, 4,
    -- layer=1 filter=73 channel=76
    -2, -6, -4, -2, -10, -10, 8, 7, 8,
    -- layer=1 filter=73 channel=77
    -10, 5, 3, 3, -1, -4, -9, -6, -5,
    -- layer=1 filter=73 channel=78
    -3, -7, 4, 9, -2, -11, 4, -4, 5,
    -- layer=1 filter=73 channel=79
    -1, 2, -5, -10, -5, -11, -2, 7, 4,
    -- layer=1 filter=73 channel=80
    -8, 0, -2, -7, -6, -1, 0, -9, -2,
    -- layer=1 filter=73 channel=81
    -1, 0, -1, 8, 1, -8, 0, -1, 7,
    -- layer=1 filter=73 channel=82
    -12, -9, -7, 0, -4, -5, -9, 7, -3,
    -- layer=1 filter=73 channel=83
    8, -1, -5, 3, -4, 5, -9, 8, -7,
    -- layer=1 filter=73 channel=84
    -1, 2, 3, 0, -15, -12, -1, -9, 2,
    -- layer=1 filter=73 channel=85
    7, -8, 0, -2, -2, 5, -4, -1, -1,
    -- layer=1 filter=73 channel=86
    -9, 5, -8, 2, -11, -6, -6, 7, 3,
    -- layer=1 filter=73 channel=87
    -4, 7, 5, 2, 5, -4, 1, 6, -1,
    -- layer=1 filter=73 channel=88
    -6, -7, 0, -8, -11, -5, 0, 6, -1,
    -- layer=1 filter=73 channel=89
    1, 4, -6, 6, 4, -1, -7, -10, -2,
    -- layer=1 filter=73 channel=90
    -3, -10, 4, -7, -7, -3, 6, 7, -5,
    -- layer=1 filter=73 channel=91
    -5, -1, -2, -4, -11, 2, -6, -10, -11,
    -- layer=1 filter=73 channel=92
    -9, -8, -3, -2, 0, -1, 7, 0, -6,
    -- layer=1 filter=73 channel=93
    0, 6, 3, 1, 3, -11, -9, -8, -9,
    -- layer=1 filter=73 channel=94
    7, 0, -5, -1, 7, -9, -7, -7, -9,
    -- layer=1 filter=73 channel=95
    -1, 4, -8, -11, 3, -6, 6, 3, -1,
    -- layer=1 filter=73 channel=96
    5, 0, 6, -2, 7, -2, 5, -8, -1,
    -- layer=1 filter=73 channel=97
    7, -2, -2, 0, 0, 4, 0, 7, -1,
    -- layer=1 filter=73 channel=98
    -6, 5, 5, 9, 0, 8, 0, -7, -9,
    -- layer=1 filter=73 channel=99
    -2, -1, 6, -1, -4, 5, -11, 5, 4,
    -- layer=1 filter=73 channel=100
    0, -7, -9, 0, 5, 0, 2, 2, 3,
    -- layer=1 filter=73 channel=101
    -9, -5, 4, 6, 8, -9, -2, -9, 2,
    -- layer=1 filter=73 channel=102
    6, -6, -1, -2, 0, -2, 0, 5, 4,
    -- layer=1 filter=73 channel=103
    -10, -5, -7, 5, 1, 8, -11, -12, -9,
    -- layer=1 filter=73 channel=104
    -9, -5, -5, -8, 5, -8, -2, -10, 7,
    -- layer=1 filter=73 channel=105
    8, 5, 1, 4, 1, 5, -10, 3, -9,
    -- layer=1 filter=73 channel=106
    1, 0, -12, -7, -12, 0, 2, 0, -3,
    -- layer=1 filter=73 channel=107
    6, -3, 7, -4, -4, 8, -10, -7, 2,
    -- layer=1 filter=73 channel=108
    -9, 12, 3, 1, 0, -8, -4, -5, -11,
    -- layer=1 filter=73 channel=109
    -5, 6, 1, -8, -2, 0, -6, 1, -2,
    -- layer=1 filter=73 channel=110
    5, -9, 8, -7, -7, -3, 3, -4, -8,
    -- layer=1 filter=73 channel=111
    1, -14, 2, -2, -16, -6, 5, 8, 4,
    -- layer=1 filter=73 channel=112
    -11, 8, -9, -9, 4, -4, -9, 1, -8,
    -- layer=1 filter=73 channel=113
    0, -6, -1, -1, -12, -10, 0, 3, -10,
    -- layer=1 filter=73 channel=114
    2, 2, 2, 0, 4, -9, -4, -6, -9,
    -- layer=1 filter=73 channel=115
    -11, -11, 5, -4, -11, 5, 1, -2, -11,
    -- layer=1 filter=73 channel=116
    8, 9, 9, 0, -7, -6, -6, -5, 0,
    -- layer=1 filter=73 channel=117
    -10, -1, 7, 3, -9, 6, 7, -8, 4,
    -- layer=1 filter=73 channel=118
    -5, -2, -4, -6, -5, -13, -3, 3, -2,
    -- layer=1 filter=73 channel=119
    -3, -1, 1, -4, 5, 0, -9, 1, -1,
    -- layer=1 filter=73 channel=120
    7, -5, -5, 6, 7, -5, -4, -3, 5,
    -- layer=1 filter=73 channel=121
    7, 4, -3, -9, -7, -14, -4, 0, -3,
    -- layer=1 filter=73 channel=122
    -9, 1, 1, 10, -5, 8, 2, 1, 0,
    -- layer=1 filter=73 channel=123
    -5, 8, -10, 5, -12, 1, -7, -4, -3,
    -- layer=1 filter=73 channel=124
    -4, -5, 0, -9, 4, -5, -7, -7, 6,
    -- layer=1 filter=73 channel=125
    2, 6, -2, 12, 3, -2, 5, 5, -7,
    -- layer=1 filter=73 channel=126
    6, 7, 9, -6, -5, 4, -9, -1, 0,
    -- layer=1 filter=73 channel=127
    1, 7, -10, 2, -7, -10, 0, 7, -7,
    -- layer=1 filter=74 channel=0
    2, -8, 6, -5, -8, 5, 3, 4, -11,
    -- layer=1 filter=74 channel=1
    -12, 7, 5, 7, 8, 2, -10, -2, -7,
    -- layer=1 filter=74 channel=2
    -4, -10, -2, 1, 0, 1, -13, 2, -9,
    -- layer=1 filter=74 channel=3
    -5, -9, -1, 3, 4, 1, 10, -3, -7,
    -- layer=1 filter=74 channel=4
    -5, 8, -7, -7, -2, -4, 6, 1, 5,
    -- layer=1 filter=74 channel=5
    -7, -9, 4, -6, 4, 3, -7, -1, -7,
    -- layer=1 filter=74 channel=6
    -2, 5, -9, -7, -5, 4, -7, -5, 10,
    -- layer=1 filter=74 channel=7
    -12, 0, 7, -14, -9, -7, 2, 0, -8,
    -- layer=1 filter=74 channel=8
    -6, -1, -7, -10, -6, -1, -6, -8, -3,
    -- layer=1 filter=74 channel=9
    1, -8, -15, 2, -4, -5, -14, -9, 1,
    -- layer=1 filter=74 channel=10
    0, -2, -7, -13, -5, -1, -10, -11, 0,
    -- layer=1 filter=74 channel=11
    0, 4, -7, 2, -1, -5, 1, -1, 0,
    -- layer=1 filter=74 channel=12
    3, -14, -2, -13, -7, 0, 0, 2, 5,
    -- layer=1 filter=74 channel=13
    -12, 1, 4, 5, -8, 2, -4, -10, 3,
    -- layer=1 filter=74 channel=14
    3, 0, -7, -10, -5, -10, -12, 0, -6,
    -- layer=1 filter=74 channel=15
    -3, -5, -2, -11, -6, 2, 4, -2, -4,
    -- layer=1 filter=74 channel=16
    -6, 1, -7, 8, -3, -5, 1, -7, 4,
    -- layer=1 filter=74 channel=17
    -3, -11, -2, -6, -12, -8, -11, 2, -3,
    -- layer=1 filter=74 channel=18
    -5, 1, -7, -12, -10, 0, 9, -7, -7,
    -- layer=1 filter=74 channel=19
    -4, -10, 5, 6, -1, -10, 7, 7, 4,
    -- layer=1 filter=74 channel=20
    -10, 7, -1, 0, -9, -3, 4, 2, 4,
    -- layer=1 filter=74 channel=21
    2, -11, -8, -1, -12, -14, -7, 3, -13,
    -- layer=1 filter=74 channel=22
    2, 3, 5, 0, -3, -5, -1, -10, -8,
    -- layer=1 filter=74 channel=23
    6, 1, -6, -6, -9, 3, 2, 2, 2,
    -- layer=1 filter=74 channel=24
    -3, 0, -8, -12, -5, 1, -14, 2, 1,
    -- layer=1 filter=74 channel=25
    -14, -2, 5, -12, -12, 6, 10, 2, -7,
    -- layer=1 filter=74 channel=26
    -4, -13, 0, -7, -12, -12, -3, 4, -12,
    -- layer=1 filter=74 channel=27
    -2, -8, -4, -5, -13, 1, -5, -8, -11,
    -- layer=1 filter=74 channel=28
    -12, 5, -7, -1, -6, 0, -2, -11, 3,
    -- layer=1 filter=74 channel=29
    5, 1, 1, 7, -5, -11, -10, 0, -2,
    -- layer=1 filter=74 channel=30
    6, -4, 0, 1, 10, 0, -5, 2, 7,
    -- layer=1 filter=74 channel=31
    -5, 0, -14, -8, -13, 1, 0, -3, 1,
    -- layer=1 filter=74 channel=32
    2, 1, -9, 8, 5, -8, 7, -1, 0,
    -- layer=1 filter=74 channel=33
    -5, -5, -7, 4, 10, 2, -1, -4, 5,
    -- layer=1 filter=74 channel=34
    0, -5, -12, 5, -10, 0, -9, -8, -6,
    -- layer=1 filter=74 channel=35
    -4, 5, -4, 0, 8, -9, 6, -5, -1,
    -- layer=1 filter=74 channel=36
    7, -3, 7, -9, -11, 6, -7, -8, -4,
    -- layer=1 filter=74 channel=37
    -2, -5, -8, 0, -3, -8, 5, 2, -11,
    -- layer=1 filter=74 channel=38
    -7, -7, 1, -9, -8, -10, -8, 2, 7,
    -- layer=1 filter=74 channel=39
    -6, -8, 7, 4, -3, -4, -10, 0, 0,
    -- layer=1 filter=74 channel=40
    -12, 0, -1, -5, -9, 0, -2, -15, -1,
    -- layer=1 filter=74 channel=41
    -3, 0, 1, -9, -2, 4, 2, 1, -9,
    -- layer=1 filter=74 channel=42
    -1, -6, 0, -11, -14, -8, -12, -6, 0,
    -- layer=1 filter=74 channel=43
    2, -5, 7, 0, -11, -2, -6, -5, 5,
    -- layer=1 filter=74 channel=44
    -6, 6, -5, -7, -5, -1, -2, -11, 7,
    -- layer=1 filter=74 channel=45
    5, 0, -9, 1, 4, -5, -10, -9, -15,
    -- layer=1 filter=74 channel=46
    6, 1, -14, 0, 2, -6, -5, -2, -1,
    -- layer=1 filter=74 channel=47
    1, -5, -15, -1, -4, -9, 4, -8, -6,
    -- layer=1 filter=74 channel=48
    -5, 4, 5, -8, -8, -11, 2, 5, 0,
    -- layer=1 filter=74 channel=49
    -5, -3, 0, 1, 1, -3, -15, 0, -14,
    -- layer=1 filter=74 channel=50
    2, 0, -8, -9, -8, 4, 5, -6, 7,
    -- layer=1 filter=74 channel=51
    -5, -8, 0, -5, 0, 2, 3, 2, -13,
    -- layer=1 filter=74 channel=52
    -9, 10, -3, -5, -9, 0, 6, 0, -9,
    -- layer=1 filter=74 channel=53
    -4, 0, 6, 0, -9, -2, -2, -12, 2,
    -- layer=1 filter=74 channel=54
    -13, -9, 1, 1, 2, -7, 1, 0, 0,
    -- layer=1 filter=74 channel=55
    -8, 2, -12, -6, -12, -17, -5, 0, -5,
    -- layer=1 filter=74 channel=56
    -6, 4, 3, -8, -7, 7, -8, -2, -4,
    -- layer=1 filter=74 channel=57
    -9, -2, -3, -2, -13, 1, -7, 0, 5,
    -- layer=1 filter=74 channel=58
    -4, -9, -1, -11, -3, 1, -8, 1, 0,
    -- layer=1 filter=74 channel=59
    -10, 5, 2, -1, 0, 7, 0, 6, 0,
    -- layer=1 filter=74 channel=60
    3, -6, -2, -2, -4, 1, 7, 7, 5,
    -- layer=1 filter=74 channel=61
    -5, -3, 2, 7, 7, 4, 6, -6, 7,
    -- layer=1 filter=74 channel=62
    -9, 3, -2, 0, -9, -4, 9, 3, 4,
    -- layer=1 filter=74 channel=63
    -7, -4, 1, -4, 8, 4, 0, -5, -2,
    -- layer=1 filter=74 channel=64
    -3, -1, 0, 4, -6, -2, -10, -3, -6,
    -- layer=1 filter=74 channel=65
    -7, -10, -5, 0, 0, 5, -6, -2, -1,
    -- layer=1 filter=74 channel=66
    -12, -10, 0, -8, -10, -6, -12, 2, 4,
    -- layer=1 filter=74 channel=67
    -10, -2, -5, 1, -9, -7, 3, 10, 8,
    -- layer=1 filter=74 channel=68
    0, -3, -4, 7, -5, -10, -9, 3, 7,
    -- layer=1 filter=74 channel=69
    -7, -3, 0, -11, -13, -10, -1, -4, -6,
    -- layer=1 filter=74 channel=70
    4, 7, -1, -10, -6, 2, 6, -6, 6,
    -- layer=1 filter=74 channel=71
    3, -3, -1, 0, 5, -1, -7, 1, 2,
    -- layer=1 filter=74 channel=72
    1, 8, 4, 3, -12, -8, -9, 8, -12,
    -- layer=1 filter=74 channel=73
    5, -5, 4, -3, -11, -4, -5, -5, -5,
    -- layer=1 filter=74 channel=74
    3, -6, -1, 0, -12, -8, -6, -4, -2,
    -- layer=1 filter=74 channel=75
    -7, 0, -2, 3, -11, -11, 0, 2, -9,
    -- layer=1 filter=74 channel=76
    -6, 0, 7, 0, -11, -12, -2, 0, 4,
    -- layer=1 filter=74 channel=77
    2, 1, -6, 3, 5, -5, 7, 5, -4,
    -- layer=1 filter=74 channel=78
    -3, 1, -4, 7, 7, 1, 5, -11, 4,
    -- layer=1 filter=74 channel=79
    0, -3, 1, -9, 2, 0, -5, 6, -11,
    -- layer=1 filter=74 channel=80
    -10, 0, 3, 3, 0, 4, 7, 4, -2,
    -- layer=1 filter=74 channel=81
    3, 3, -5, -7, -2, -1, -2, -6, -1,
    -- layer=1 filter=74 channel=82
    5, -12, 2, 5, 2, -5, 1, -12, -6,
    -- layer=1 filter=74 channel=83
    -10, 0, -3, -4, -8, 6, -7, 1, -1,
    -- layer=1 filter=74 channel=84
    0, 0, 8, -10, 5, -5, 6, 0, -9,
    -- layer=1 filter=74 channel=85
    -3, -6, -8, 4, 2, 5, -12, -9, 4,
    -- layer=1 filter=74 channel=86
    -6, -6, 9, 4, -10, -10, -8, -11, 2,
    -- layer=1 filter=74 channel=87
    3, -11, 0, -2, -11, -11, 4, -5, -6,
    -- layer=1 filter=74 channel=88
    -15, -12, -5, 0, 2, -4, -6, -7, -11,
    -- layer=1 filter=74 channel=89
    2, -3, 1, 4, -11, 3, 2, 0, -6,
    -- layer=1 filter=74 channel=90
    -12, -12, 3, -7, 8, -1, -12, -2, -3,
    -- layer=1 filter=74 channel=91
    0, -10, -3, -2, -11, -8, 4, -10, -7,
    -- layer=1 filter=74 channel=92
    -10, -1, -9, -4, 2, 0, -14, -12, 0,
    -- layer=1 filter=74 channel=93
    -12, -10, -4, -3, -3, 0, -10, -11, -3,
    -- layer=1 filter=74 channel=94
    6, -9, -7, -9, 6, 5, -7, 2, -1,
    -- layer=1 filter=74 channel=95
    5, 2, -10, -10, 0, 0, -7, 3, 8,
    -- layer=1 filter=74 channel=96
    -3, -5, -12, -1, -10, 6, 0, -11, 7,
    -- layer=1 filter=74 channel=97
    0, 1, 1, -5, 5, 5, -2, -4, -11,
    -- layer=1 filter=74 channel=98
    3, -5, 0, 2, -4, -5, 9, -3, -13,
    -- layer=1 filter=74 channel=99
    2, -10, -4, -7, 5, -3, 3, 6, -1,
    -- layer=1 filter=74 channel=100
    -12, -10, -8, -9, 6, 0, 5, 6, -2,
    -- layer=1 filter=74 channel=101
    -8, -2, -4, -2, 0, 3, 1, -12, -5,
    -- layer=1 filter=74 channel=102
    -1, -7, -8, -10, 5, -3, -1, 3, 8,
    -- layer=1 filter=74 channel=103
    -7, -7, -3, -5, 4, -4, 0, 5, -9,
    -- layer=1 filter=74 channel=104
    -9, -10, -8, -12, -11, -1, -4, -11, -1,
    -- layer=1 filter=74 channel=105
    -12, 2, -3, 3, -7, 4, -1, -5, 1,
    -- layer=1 filter=74 channel=106
    -10, -2, 4, -12, 5, -9, -4, -12, -2,
    -- layer=1 filter=74 channel=107
    7, 8, 2, 1, -7, 1, 10, -6, -7,
    -- layer=1 filter=74 channel=108
    5, -1, -9, 3, -1, -3, -10, 6, 0,
    -- layer=1 filter=74 channel=109
    1, 11, 9, 8, 3, -7, 0, -5, 0,
    -- layer=1 filter=74 channel=110
    6, 2, 7, -9, -4, -9, -2, 3, 5,
    -- layer=1 filter=74 channel=111
    -10, 4, 6, -5, 0, -10, 5, -10, 0,
    -- layer=1 filter=74 channel=112
    0, 0, -3, -11, -1, -3, -9, -12, 1,
    -- layer=1 filter=74 channel=113
    -14, -9, -11, -2, -9, -4, -14, -9, -11,
    -- layer=1 filter=74 channel=114
    0, -9, 2, 6, -9, -9, 1, -8, 4,
    -- layer=1 filter=74 channel=115
    -2, 0, 4, 3, 7, 2, -9, -6, 4,
    -- layer=1 filter=74 channel=116
    0, -1, -7, 8, -8, -6, -7, -1, 5,
    -- layer=1 filter=74 channel=117
    0, -8, -8, 2, -5, 6, -7, 0, -5,
    -- layer=1 filter=74 channel=118
    3, 2, 0, 2, -1, 5, -7, 3, 4,
    -- layer=1 filter=74 channel=119
    -12, 1, -8, 1, 0, -1, -6, -6, -10,
    -- layer=1 filter=74 channel=120
    -16, 2, 0, -5, 4, 4, -5, -18, -7,
    -- layer=1 filter=74 channel=121
    -14, -14, -6, -3, -13, -4, -16, -4, 0,
    -- layer=1 filter=74 channel=122
    0, 4, -7, -9, 0, -1, -2, -2, 8,
    -- layer=1 filter=74 channel=123
    -14, 3, 4, 3, -15, -15, -11, 2, -10,
    -- layer=1 filter=74 channel=124
    -6, -10, 1, -3, 0, -9, -8, -7, -5,
    -- layer=1 filter=74 channel=125
    1, -7, 8, -13, 2, 2, -12, 0, 0,
    -- layer=1 filter=74 channel=126
    3, 6, 8, -3, 3, -2, 4, 1, -6,
    -- layer=1 filter=74 channel=127
    -8, -6, 9, -1, 3, -2, -4, -7, 5,
    -- layer=1 filter=75 channel=0
    -18, -19, -7, 0, 4, 21, -5, 12, 9,
    -- layer=1 filter=75 channel=1
    -16, 26, 19, 12, 2, 25, 18, 18, -28,
    -- layer=1 filter=75 channel=2
    20, 24, 36, 15, -11, 33, 19, 30, 39,
    -- layer=1 filter=75 channel=3
    8, -1, -3, -8, -6, 5, 1, 10, 11,
    -- layer=1 filter=75 channel=4
    2, 10, 1, -7, -6, 6, -1, 1, -8,
    -- layer=1 filter=75 channel=5
    0, 54, 46, 27, 31, 30, 35, 29, -35,
    -- layer=1 filter=75 channel=6
    48, 73, 53, 50, -32, -47, 5, -58, 0,
    -- layer=1 filter=75 channel=7
    -21, -3, 14, 14, 23, -36, 9, 46, -18,
    -- layer=1 filter=75 channel=8
    1, 32, 34, 5, 19, 34, 30, 9, -24,
    -- layer=1 filter=75 channel=9
    17, 38, 12, 29, 15, 14, 1, 22, 7,
    -- layer=1 filter=75 channel=10
    12, 15, 25, 2, 29, -23, 8, 36, -11,
    -- layer=1 filter=75 channel=11
    -23, -24, -27, 4, 23, 28, 9, 14, 20,
    -- layer=1 filter=75 channel=12
    13, 0, 3, 6, 7, -50, 26, 1, 18,
    -- layer=1 filter=75 channel=13
    36, 7, 9, 4, -18, -25, -5, -38, -52,
    -- layer=1 filter=75 channel=14
    -42, -28, 26, 3, 5, -51, -18, 13, -14,
    -- layer=1 filter=75 channel=15
    7, -7, 1, -6, -13, 15, 27, -1, -33,
    -- layer=1 filter=75 channel=16
    -28, 18, 22, 3, 34, 19, 34, 27, -39,
    -- layer=1 filter=75 channel=17
    19, 10, 16, -10, 5, 24, -17, -18, 11,
    -- layer=1 filter=75 channel=18
    -28, -12, -26, 26, 16, 2, 30, 23, 30,
    -- layer=1 filter=75 channel=19
    27, 21, 47, 20, 49, 2, 7, 19, -23,
    -- layer=1 filter=75 channel=20
    18, 20, -4, -1, -27, -19, -6, -36, -14,
    -- layer=1 filter=75 channel=21
    -16, 6, -19, -7, -44, -9, -34, -45, -68,
    -- layer=1 filter=75 channel=22
    6, 8, -11, 0, -25, -2, -12, -29, -24,
    -- layer=1 filter=75 channel=23
    -18, -14, -18, -27, 24, -35, -1, 22, -6,
    -- layer=1 filter=75 channel=24
    11, -17, -22, -35, -11, -18, -15, -77, -61,
    -- layer=1 filter=75 channel=25
    -2, 21, 8, 24, 35, -7, 24, 39, -45,
    -- layer=1 filter=75 channel=26
    8, -24, -23, -19, -42, -27, -12, -33, -42,
    -- layer=1 filter=75 channel=27
    -31, -4, 0, 9, 10, 2, 28, 29, 11,
    -- layer=1 filter=75 channel=28
    -29, 11, 14, -8, 10, -32, 5, 34, -49,
    -- layer=1 filter=75 channel=29
    -22, -18, -7, -20, -23, -3, -12, -22, -11,
    -- layer=1 filter=75 channel=30
    -11, -28, -9, 20, 7, -13, -10, 0, 22,
    -- layer=1 filter=75 channel=31
    6, 27, 29, 20, -7, -49, 0, -18, -10,
    -- layer=1 filter=75 channel=32
    23, -24, -11, 5, -58, -53, 6, -7, -34,
    -- layer=1 filter=75 channel=33
    3, 10, 0, 7, 7, 1, 11, 2, -2,
    -- layer=1 filter=75 channel=34
    33, 3, -2, 34, 6, 1, 14, 19, 6,
    -- layer=1 filter=75 channel=35
    -8, 2, -5, -15, -11, -10, 2, 0, -7,
    -- layer=1 filter=75 channel=36
    -9, -15, 0, 17, 15, 30, 29, 38, 46,
    -- layer=1 filter=75 channel=37
    10, 51, 32, 19, 55, 36, 53, 33, -41,
    -- layer=1 filter=75 channel=38
    47, 28, -2, 14, -25, -30, -16, -50, -43,
    -- layer=1 filter=75 channel=39
    -30, 7, 0, -12, 24, 19, 22, 17, 6,
    -- layer=1 filter=75 channel=40
    -12, 3, 3, 6, -17, -84, -30, -32, -25,
    -- layer=1 filter=75 channel=41
    39, 21, -30, 30, -18, -36, 19, 1, -24,
    -- layer=1 filter=75 channel=42
    14, 34, 48, 8, 29, 26, 23, 34, 41,
    -- layer=1 filter=75 channel=43
    -34, 37, 27, 0, 8, 18, 37, 34, -28,
    -- layer=1 filter=75 channel=44
    20, -36, -8, -28, -61, -25, -8, -18, -40,
    -- layer=1 filter=75 channel=45
    5, 1, 8, -31, -6, 0, 9, -21, -52,
    -- layer=1 filter=75 channel=46
    38, 23, 69, 9, 48, 58, 50, 13, -11,
    -- layer=1 filter=75 channel=47
    35, 19, 16, 12, 19, -25, 23, 9, 19,
    -- layer=1 filter=75 channel=48
    2, -13, -21, -21, -9, -30, -35, -28, -30,
    -- layer=1 filter=75 channel=49
    20, 21, 36, 13, 0, 3, 10, -3, 10,
    -- layer=1 filter=75 channel=50
    4, -23, 3, 8, 4, -21, 0, 15, 9,
    -- layer=1 filter=75 channel=51
    -8, -13, -1, -38, -19, -65, -38, -30, -41,
    -- layer=1 filter=75 channel=52
    5, -17, -31, 2, -7, 20, 10, 10, -2,
    -- layer=1 filter=75 channel=53
    0, -1, 17, 4, 1, 14, 1, -4, 9,
    -- layer=1 filter=75 channel=54
    0, 39, 41, 20, 55, 2, 38, 59, -46,
    -- layer=1 filter=75 channel=55
    -20, -22, -6, 7, 7, 13, 15, 9, 21,
    -- layer=1 filter=75 channel=56
    -9, -9, -7, -6, -6, -9, 7, 7, -3,
    -- layer=1 filter=75 channel=57
    8, 6, 27, 11, 20, -55, -1, 19, -23,
    -- layer=1 filter=75 channel=58
    2, 0, -4, -11, 29, -40, -8, 36, -20,
    -- layer=1 filter=75 channel=59
    -5, 0, 12, 5, 1, -5, -11, -4, 1,
    -- layer=1 filter=75 channel=60
    1, 14, 6, 2, 15, 7, 15, 13, 5,
    -- layer=1 filter=75 channel=61
    4, -10, -2, -3, 7, -9, 3, 9, 0,
    -- layer=1 filter=75 channel=62
    -4, 46, 20, 15, 37, 32, 44, 10, -35,
    -- layer=1 filter=75 channel=63
    -29, -46, -33, 21, 3, 6, 28, 40, 31,
    -- layer=1 filter=75 channel=64
    9, 24, 12, 7, 10, 9, 15, 4, -10,
    -- layer=1 filter=75 channel=65
    -4, 6, -25, -15, -25, -21, -31, -37, -22,
    -- layer=1 filter=75 channel=66
    -5, -5, -3, 7, 12, 24, 10, 24, 21,
    -- layer=1 filter=75 channel=67
    4, 18, 31, 28, 18, 0, 45, 27, -2,
    -- layer=1 filter=75 channel=68
    4, -27, -24, -22, -61, -19, -13, 0, -31,
    -- layer=1 filter=75 channel=69
    -14, 8, 19, -15, 0, 21, 43, 0, -46,
    -- layer=1 filter=75 channel=70
    34, 45, 26, 7, -40, -47, 38, -46, -2,
    -- layer=1 filter=75 channel=71
    -33, -22, -17, -20, -28, -13, -13, -9, -42,
    -- layer=1 filter=75 channel=72
    28, -7, 37, 31, 1, -1, 2, 3, 23,
    -- layer=1 filter=75 channel=73
    -9, 0, 0, -1, -6, 5, 4, -6, -5,
    -- layer=1 filter=75 channel=74
    -16, 33, -19, 15, -29, -19, -12, 9, -12,
    -- layer=1 filter=75 channel=75
    -22, -9, 16, 31, 3, -35, 19, 39, 26,
    -- layer=1 filter=75 channel=76
    1, -23, -44, 0, -2, 1, -21, 15, 12,
    -- layer=1 filter=75 channel=77
    -2, -15, -42, -13, -16, -37, -30, -44, -33,
    -- layer=1 filter=75 channel=78
    -6, 0, -1, 0, -15, -19, 15, 7, -10,
    -- layer=1 filter=75 channel=79
    -3, 31, 9, -3, 23, 7, 45, 11, -29,
    -- layer=1 filter=75 channel=80
    5, -11, 6, 2, 3, 7, 4, -11, -14,
    -- layer=1 filter=75 channel=81
    -32, -17, -35, -24, -21, -21, 4, -28, -30,
    -- layer=1 filter=75 channel=82
    7, 10, -24, -25, -37, -30, -42, -56, -60,
    -- layer=1 filter=75 channel=83
    4, -13, 18, -27, -12, 1, 8, -18, -29,
    -- layer=1 filter=75 channel=84
    -40, -10, -43, 32, 1, -30, 0, 22, 11,
    -- layer=1 filter=75 channel=85
    30, 39, 4, 14, 41, 2, 12, 40, -18,
    -- layer=1 filter=75 channel=86
    -24, 2, 7, -5, 23, 26, 16, 28, 15,
    -- layer=1 filter=75 channel=87
    46, 49, 74, 18, 54, 4, 22, -1, 14,
    -- layer=1 filter=75 channel=88
    29, 11, 22, -2, -4, 1, -7, -7, 2,
    -- layer=1 filter=75 channel=89
    3, -4, -28, -13, -24, -43, -46, -29, -48,
    -- layer=1 filter=75 channel=90
    29, -29, -1, -27, -31, -1, -10, -55, -64,
    -- layer=1 filter=75 channel=91
    19, 13, -6, 12, -9, -41, -20, -45, -47,
    -- layer=1 filter=75 channel=92
    21, -1, -18, 26, -41, -33, -14, 21, -19,
    -- layer=1 filter=75 channel=93
    -20, -9, -28, -28, -15, -22, -18, -25, -32,
    -- layer=1 filter=75 channel=94
    -10, -10, 2, 14, 30, 34, 3, 34, 41,
    -- layer=1 filter=75 channel=95
    -41, -7, -31, 21, -11, -21, -10, 31, 19,
    -- layer=1 filter=75 channel=96
    -4, -10, -5, 8, 2, 15, 11, 2, 12,
    -- layer=1 filter=75 channel=97
    -12, -20, 0, -7, 0, 1, 8, 7, -2,
    -- layer=1 filter=75 channel=98
    4, 25, 9, 2, 25, 21, 2, -6, -35,
    -- layer=1 filter=75 channel=99
    -29, -43, -6, -42, -22, -7, -31, 2, -31,
    -- layer=1 filter=75 channel=100
    -23, -12, -7, 27, 12, 9, 34, 27, 28,
    -- layer=1 filter=75 channel=101
    23, 6, 7, -6, -35, -35, -29, -42, -41,
    -- layer=1 filter=75 channel=102
    -4, -5, 12, 3, 19, 34, -14, -6, 34,
    -- layer=1 filter=75 channel=103
    -14, 0, -6, 24, 11, -6, 7, 27, 19,
    -- layer=1 filter=75 channel=104
    34, 19, 10, -3, 31, 3, 20, 40, 14,
    -- layer=1 filter=75 channel=105
    -25, -25, -3, 6, 4, 9, -7, 15, 11,
    -- layer=1 filter=75 channel=106
    34, 16, 8, 0, -51, -55, -24, -32, -41,
    -- layer=1 filter=75 channel=107
    5, 16, 13, 15, -1, 6, -7, -20, -15,
    -- layer=1 filter=75 channel=108
    11, -35, -26, -28, -59, -37, -17, -45, -46,
    -- layer=1 filter=75 channel=109
    8, 3, 3, 4, -5, -9, 5, -4, 10,
    -- layer=1 filter=75 channel=110
    -9, -7, -11, -1, -2, 0, 3, -12, -10,
    -- layer=1 filter=75 channel=111
    -29, -21, -29, 27, 26, -17, 0, 9, 21,
    -- layer=1 filter=75 channel=112
    -20, -16, -22, 35, 30, -3, 22, 23, 23,
    -- layer=1 filter=75 channel=113
    38, 17, 28, 15, 9, -13, 9, -17, -11,
    -- layer=1 filter=75 channel=114
    -32, 14, 28, 2, 22, 32, 51, 26, -24,
    -- layer=1 filter=75 channel=115
    -22, -12, 14, -9, 20, 20, -2, 36, 29,
    -- layer=1 filter=75 channel=116
    4, -5, -5, 7, -7, -3, 0, -2, -9,
    -- layer=1 filter=75 channel=117
    -45, -61, -29, 19, 46, -24, 13, 7, 40,
    -- layer=1 filter=75 channel=118
    -14, 2, -16, 1, -11, -7, -1, 6, -9,
    -- layer=1 filter=75 channel=119
    18, -32, -21, -13, -59, -28, 0, -43, -44,
    -- layer=1 filter=75 channel=120
    13, 18, -8, -7, -1, -39, -20, -23, -34,
    -- layer=1 filter=75 channel=121
    -15, -9, -13, -5, -3, 0, 1, 17, 17,
    -- layer=1 filter=75 channel=122
    11, -3, -10, 3, 5, 9, -4, 2, 8,
    -- layer=1 filter=75 channel=123
    -30, -37, -38, 18, 12, -5, 21, 32, 16,
    -- layer=1 filter=75 channel=124
    7, 6, 5, 1, -11, 2, -3, -6, 0,
    -- layer=1 filter=75 channel=125
    35, 40, 26, 1, -18, -43, 0, -7, -25,
    -- layer=1 filter=75 channel=126
    19, 35, 0, 30, 45, 38, 17, -30, -25,
    -- layer=1 filter=75 channel=127
    -35, -3, -17, 19, 15, -17, 0, 18, 10,
    -- layer=1 filter=76 channel=0
    -4, 2, -16, -8, 2, -9, 6, 6, -13,
    -- layer=1 filter=76 channel=1
    -26, 13, -20, 13, 3, -14, 32, -31, 16,
    -- layer=1 filter=76 channel=2
    18, 14, 21, -35, -13, 7, -5, -5, 3,
    -- layer=1 filter=76 channel=3
    -13, 0, 0, -13, 7, 3, -12, 7, 1,
    -- layer=1 filter=76 channel=4
    -4, -12, -22, -13, 0, -11, 0, -19, -6,
    -- layer=1 filter=76 channel=5
    -16, 20, -9, 2, -3, 7, 34, -35, 10,
    -- layer=1 filter=76 channel=6
    -3, -16, 12, 11, 6, 0, 27, 25, 8,
    -- layer=1 filter=76 channel=7
    40, -4, -23, 57, -12, 18, 40, -24, 39,
    -- layer=1 filter=76 channel=8
    -15, 4, -12, 0, 1, -10, -2, -29, 23,
    -- layer=1 filter=76 channel=9
    -38, -10, 11, -39, 13, -22, -66, -23, -18,
    -- layer=1 filter=76 channel=10
    22, -20, -34, 56, -28, 1, 37, -24, 0,
    -- layer=1 filter=76 channel=11
    -11, 7, 6, -14, 4, 13, -12, 27, 5,
    -- layer=1 filter=76 channel=12
    -1, -36, -7, -19, -36, 14, -25, -25, 25,
    -- layer=1 filter=76 channel=13
    -21, 5, 22, -31, 12, 2, -15, 24, 14,
    -- layer=1 filter=76 channel=14
    13, -5, 5, 5, -33, -29, 10, -13, 9,
    -- layer=1 filter=76 channel=15
    -11, 12, -1, -21, 8, 45, 7, -17, 2,
    -- layer=1 filter=76 channel=16
    -2, 15, -16, 20, -21, -3, 7, -37, -1,
    -- layer=1 filter=76 channel=17
    -7, -13, -8, -15, -1, -19, -24, 0, -8,
    -- layer=1 filter=76 channel=18
    12, -7, 1, -15, -24, 0, -21, -9, -1,
    -- layer=1 filter=76 channel=19
    15, -23, -32, -12, -39, 0, -2, -7, -15,
    -- layer=1 filter=76 channel=20
    5, -1, -15, 5, -6, -5, 14, 9, 0,
    -- layer=1 filter=76 channel=21
    5, -4, -24, 26, -5, -28, 20, -5, -20,
    -- layer=1 filter=76 channel=22
    13, 10, -20, 9, 13, -21, 27, 2, -12,
    -- layer=1 filter=76 channel=23
    14, 13, -7, 45, 14, 59, 26, 18, 27,
    -- layer=1 filter=76 channel=24
    -12, 7, 20, -44, 19, 29, -30, 38, 23,
    -- layer=1 filter=76 channel=25
    30, -21, -37, 55, -42, -11, 56, -35, 4,
    -- layer=1 filter=76 channel=26
    -62, -4, 34, -91, 22, 30, -69, 25, 26,
    -- layer=1 filter=76 channel=27
    6, 11, 3, 10, 0, -1, -7, -1, -3,
    -- layer=1 filter=76 channel=28
    12, -8, -52, 42, -6, -43, 43, -14, -13,
    -- layer=1 filter=76 channel=29
    23, 28, 27, 14, 2, 8, 14, 10, 6,
    -- layer=1 filter=76 channel=30
    15, -34, 9, -22, -31, 14, -35, -20, -15,
    -- layer=1 filter=76 channel=31
    7, 2, 24, 2, -1, -14, 2, 8, 0,
    -- layer=1 filter=76 channel=32
    -38, 16, 44, -72, 34, 48, -44, 55, 48,
    -- layer=1 filter=76 channel=33
    -4, 4, 2, 7, -2, -8, 0, 0, 10,
    -- layer=1 filter=76 channel=34
    -21, -27, -2, -21, -1, -31, -25, -13, 2,
    -- layer=1 filter=76 channel=35
    0, 13, -3, -13, 11, 13, 9, -7, 2,
    -- layer=1 filter=76 channel=36
    -2, 2, -3, -18, 21, 10, -17, 17, 1,
    -- layer=1 filter=76 channel=37
    7, 7, -18, 3, -15, 8, 18, -4, 15,
    -- layer=1 filter=76 channel=38
    1, 2, -9, 4, 12, -25, 14, 2, -15,
    -- layer=1 filter=76 channel=39
    -8, 10, -6, 8, 5, -13, 5, 6, 8,
    -- layer=1 filter=76 channel=40
    27, -2, 0, 9, -10, -37, 7, -9, -29,
    -- layer=1 filter=76 channel=41
    39, -5, 41, -30, 0, 19, -21, 18, 21,
    -- layer=1 filter=76 channel=42
    13, 0, 17, -2, -44, 12, -11, -38, 5,
    -- layer=1 filter=76 channel=43
    8, -13, -33, 23, -7, -2, 50, -48, 25,
    -- layer=1 filter=76 channel=44
    -73, 4, 36, -102, 42, 36, -43, 31, 30,
    -- layer=1 filter=76 channel=45
    -16, 2, -16, -32, 22, 1, -4, 17, 16,
    -- layer=1 filter=76 channel=46
    21, -8, -28, 7, -15, 44, 34, -9, 5,
    -- layer=1 filter=76 channel=47
    16, 27, 23, 21, 33, 43, -17, 22, 29,
    -- layer=1 filter=76 channel=48
    21, -16, -6, 21, 2, -25, 13, 1, -6,
    -- layer=1 filter=76 channel=49
    7, 6, 9, -4, -3, 7, 4, 4, -2,
    -- layer=1 filter=76 channel=50
    0, 10, 3, -4, -14, 1, -13, 0, -13,
    -- layer=1 filter=76 channel=51
    18, -18, -36, 38, -19, -46, 36, -13, -27,
    -- layer=1 filter=76 channel=52
    4, 18, -6, -12, 6, 1, 6, 2, -4,
    -- layer=1 filter=76 channel=53
    -3, 3, -15, 2, 13, 3, -3, 0, -16,
    -- layer=1 filter=76 channel=54
    18, -9, -34, 45, -30, 19, 39, -15, 21,
    -- layer=1 filter=76 channel=55
    -5, 4, 16, -12, 7, 24, -13, 23, 17,
    -- layer=1 filter=76 channel=56
    15, 16, -7, -2, 5, 2, 7, 1, 0,
    -- layer=1 filter=76 channel=57
    45, -18, -51, 54, -33, -12, 41, -6, 1,
    -- layer=1 filter=76 channel=58
    48, 1, 48, 101, -20, 97, 43, 8, 56,
    -- layer=1 filter=76 channel=59
    2, 1, -36, -4, 1, -29, 1, 2, -1,
    -- layer=1 filter=76 channel=60
    -1, 10, 8, 12, 11, -10, 11, 10, 3,
    -- layer=1 filter=76 channel=61
    -12, -1, 1, -16, -11, 4, -10, -9, -6,
    -- layer=1 filter=76 channel=62
    -9, -16, -37, -3, -19, 4, 7, -32, 10,
    -- layer=1 filter=76 channel=63
    7, -1, 10, 0, 28, 18, -10, 12, 7,
    -- layer=1 filter=76 channel=64
    13, 3, -14, 1, 8, -20, 15, -5, 1,
    -- layer=1 filter=76 channel=65
    -1, -2, -21, 22, 6, -17, 21, 3, -12,
    -- layer=1 filter=76 channel=66
    0, 3, 2, 0, 19, -16, 2, 12, -3,
    -- layer=1 filter=76 channel=67
    -34, -17, 1, 10, -19, 3, 1, 6, 24,
    -- layer=1 filter=76 channel=68
    -50, 38, 41, -82, 57, 37, -21, 59, 43,
    -- layer=1 filter=76 channel=69
    -24, 26, -4, -43, 19, 21, -10, 15, 17,
    -- layer=1 filter=76 channel=70
    5, -15, 13, 9, -23, -12, 19, 7, 1,
    -- layer=1 filter=76 channel=71
    4, 9, -13, 6, -22, -18, 11, -16, -5,
    -- layer=1 filter=76 channel=72
    44, -24, 0, -13, -36, -5, 0, -15, -15,
    -- layer=1 filter=76 channel=73
    0, -4, -2, 0, 12, -9, -4, 12, 3,
    -- layer=1 filter=76 channel=74
    -27, 12, -1, -44, 29, -10, -10, 36, -8,
    -- layer=1 filter=76 channel=75
    -3, -26, 11, -31, -37, 1, -10, -29, 12,
    -- layer=1 filter=76 channel=76
    -13, -3, 28, -43, 16, 10, -39, 14, -5,
    -- layer=1 filter=76 channel=77
    0, -2, -22, 19, 18, -36, 14, 17, -18,
    -- layer=1 filter=76 channel=78
    -6, 12, -24, 0, 12, -38, -2, -2, -10,
    -- layer=1 filter=76 channel=79
    4, -7, -14, 10, -18, 4, -3, -26, 12,
    -- layer=1 filter=76 channel=80
    -4, 5, 7, 15, -12, -11, 2, 5, -1,
    -- layer=1 filter=76 channel=81
    15, -7, -28, 5, -6, -8, 12, 8, 0,
    -- layer=1 filter=76 channel=82
    1, 1, -1, 6, -1, -17, 32, 1, -16,
    -- layer=1 filter=76 channel=83
    -34, 3, -26, -19, 18, 8, 12, -2, -10,
    -- layer=1 filter=76 channel=84
    -5, 3, 33, -41, 0, 21, -34, 15, 10,
    -- layer=1 filter=76 channel=85
    43, -9, 15, 66, -8, 42, 18, 5, 29,
    -- layer=1 filter=76 channel=86
    -15, 6, -2, -4, -1, 2, 0, 6, 4,
    -- layer=1 filter=76 channel=87
    25, -4, 39, 23, -2, 15, 6, 15, 8,
    -- layer=1 filter=76 channel=88
    3, -14, 0, 7, -9, -9, 3, 0, -12,
    -- layer=1 filter=76 channel=89
    -11, 7, -6, 3, 0, -8, 14, 9, -7,
    -- layer=1 filter=76 channel=90
    -36, 34, 31, -99, 61, 45, -23, 44, 47,
    -- layer=1 filter=76 channel=91
    26, -12, -17, 26, -10, -24, 12, -6, -30,
    -- layer=1 filter=76 channel=92
    -18, -22, -25, -60, 17, -7, -5, 15, 6,
    -- layer=1 filter=76 channel=93
    5, -8, -6, 9, -7, -11, 0, -3, -14,
    -- layer=1 filter=76 channel=94
    2, 5, -16, 1, -4, -18, 6, -6, -20,
    -- layer=1 filter=76 channel=95
    -25, 8, 24, -36, 2, 22, -37, 7, -11,
    -- layer=1 filter=76 channel=96
    -14, 15, 9, 1, 1, 16, -3, 12, 0,
    -- layer=1 filter=76 channel=97
    8, 5, -3, 7, 4, -10, 0, -7, -16,
    -- layer=1 filter=76 channel=98
    1, -29, -52, 25, 0, -29, 20, -43, 4,
    -- layer=1 filter=76 channel=99
    0, 29, -24, 32, 43, -30, -4, 39, -7,
    -- layer=1 filter=76 channel=100
    -24, -1, 2, -36, 17, 13, -3, 28, 6,
    -- layer=1 filter=76 channel=101
    -7, 7, -8, 9, 3, -4, 22, -7, -24,
    -- layer=1 filter=76 channel=102
    8, 16, -1, 4, -6, -35, 9, -6, -30,
    -- layer=1 filter=76 channel=103
    -23, -3, -10, -16, -4, -5, -9, 12, -4,
    -- layer=1 filter=76 channel=104
    -3, 3, 35, 5, 1, 40, -3, 12, 19,
    -- layer=1 filter=76 channel=105
    0, 4, -25, 4, -5, -29, 0, -2, -25,
    -- layer=1 filter=76 channel=106
    -36, 9, 25, -32, 19, 19, -19, 30, 17,
    -- layer=1 filter=76 channel=107
    5, 14, 3, 0, 1, 5, 5, 5, 28,
    -- layer=1 filter=76 channel=108
    -28, 13, 47, -92, 39, 59, -55, 33, 43,
    -- layer=1 filter=76 channel=109
    6, -2, -3, 8, -8, -2, -9, -10, -8,
    -- layer=1 filter=76 channel=110
    2, 5, -23, 2, -8, -21, 14, -5, -24,
    -- layer=1 filter=76 channel=111
    -3, 4, 17, -23, -17, -6, -44, -11, -33,
    -- layer=1 filter=76 channel=112
    -11, 15, 19, -24, 19, 16, -18, 7, -11,
    -- layer=1 filter=76 channel=113
    30, -1, 4, 18, -7, -8, 32, -9, -4,
    -- layer=1 filter=76 channel=114
    -26, 29, 5, -29, 19, 7, 14, -4, -8,
    -- layer=1 filter=76 channel=115
    18, 0, -43, 29, -25, -39, 17, -13, -23,
    -- layer=1 filter=76 channel=116
    4, -1, 0, -9, 2, -7, -7, 6, 0,
    -- layer=1 filter=76 channel=117
    -23, -20, -9, -11, -24, -48, -76, -40, -46,
    -- layer=1 filter=76 channel=118
    -16, 0, 38, -41, 10, 11, -29, 14, 7,
    -- layer=1 filter=76 channel=119
    -32, 14, 49, -72, 56, 65, -53, 61, 46,
    -- layer=1 filter=76 channel=120
    20, -15, -38, 49, -28, -29, 35, -11, -16,
    -- layer=1 filter=76 channel=121
    13, -13, 0, -6, -23, -2, -21, 18, 29,
    -- layer=1 filter=76 channel=122
    5, -4, -5, -7, -9, 7, 2, 2, 0,
    -- layer=1 filter=76 channel=123
    14, 0, 4, 0, -3, 17, 10, 13, 35,
    -- layer=1 filter=76 channel=124
    0, 10, 7, -9, 4, -1, 5, -11, -6,
    -- layer=1 filter=76 channel=125
    8, -18, 3, 36, -28, -2, 14, 15, 3,
    -- layer=1 filter=76 channel=126
    0, -22, -40, -4, 18, -23, -7, -42, -4,
    -- layer=1 filter=76 channel=127
    -7, 6, 26, -30, -4, 9, -21, 5, 4,
    -- layer=1 filter=77 channel=0
    -1, 2, 5, 0, 0, 7, -5, 5, 4,
    -- layer=1 filter=77 channel=1
    -11, -3, -4, 5, 3, -10, 0, -4, 5,
    -- layer=1 filter=77 channel=2
    -4, -10, 0, -6, 0, 0, 3, -8, 3,
    -- layer=1 filter=77 channel=3
    8, 7, 3, 0, 6, -8, 0, -3, -3,
    -- layer=1 filter=77 channel=4
    1, -11, -6, 1, 7, -7, 0, -8, 1,
    -- layer=1 filter=77 channel=5
    0, -5, -8, -2, -8, 11, 3, 2, -6,
    -- layer=1 filter=77 channel=6
    -2, -2, -6, 0, 3, 5, 1, 0, -4,
    -- layer=1 filter=77 channel=7
    -4, 8, 5, 8, -10, -7, 0, 3, 2,
    -- layer=1 filter=77 channel=8
    -10, 7, -9, -8, 8, 3, 7, -10, 8,
    -- layer=1 filter=77 channel=9
    -1, 9, 0, 6, 0, 2, 0, -1, -11,
    -- layer=1 filter=77 channel=10
    -2, 5, -7, 2, -2, 5, 0, 3, -6,
    -- layer=1 filter=77 channel=11
    1, -4, -9, -3, -8, -3, 9, 0, -8,
    -- layer=1 filter=77 channel=12
    -6, -10, 6, -2, 4, -7, -5, -9, 9,
    -- layer=1 filter=77 channel=13
    6, -10, -9, -10, 6, 9, -1, 7, 1,
    -- layer=1 filter=77 channel=14
    4, -10, -8, -5, -9, 0, -9, -3, 3,
    -- layer=1 filter=77 channel=15
    6, -3, 5, -7, 5, -1, -2, 1, 2,
    -- layer=1 filter=77 channel=16
    -5, 5, 0, -7, 10, 7, 1, 8, -7,
    -- layer=1 filter=77 channel=17
    -4, 1, 1, 1, -3, -4, -9, 7, -3,
    -- layer=1 filter=77 channel=18
    -6, -3, -2, -5, 1, 2, -8, 0, 1,
    -- layer=1 filter=77 channel=19
    0, 1, -1, 0, 3, 1, 2, -10, 6,
    -- layer=1 filter=77 channel=20
    2, 6, 6, 0, 2, 0, 2, -8, 0,
    -- layer=1 filter=77 channel=21
    5, -9, 0, -6, 0, 5, -11, -3, -2,
    -- layer=1 filter=77 channel=22
    6, -3, 8, 5, -3, 5, 1, -8, -1,
    -- layer=1 filter=77 channel=23
    -10, -8, -8, 2, 0, -6, 8, -7, -2,
    -- layer=1 filter=77 channel=24
    -3, -7, 6, -1, 7, -10, -10, -10, -2,
    -- layer=1 filter=77 channel=25
    6, 1, -7, 0, -5, 1, 1, -10, -10,
    -- layer=1 filter=77 channel=26
    -2, -6, -10, 0, -2, -7, -1, 6, -5,
    -- layer=1 filter=77 channel=27
    10, -2, -2, 2, -3, 0, 0, 4, -7,
    -- layer=1 filter=77 channel=28
    -2, -8, 6, 8, -2, -4, -10, -7, -8,
    -- layer=1 filter=77 channel=29
    -7, 5, 5, 3, 8, 3, 0, -6, 0,
    -- layer=1 filter=77 channel=30
    -6, -6, 6, 0, -7, 3, -12, -8, 5,
    -- layer=1 filter=77 channel=31
    -2, -6, -7, 5, 2, -3, -4, -7, -10,
    -- layer=1 filter=77 channel=32
    -7, -9, -9, -5, -5, -7, 1, 6, 9,
    -- layer=1 filter=77 channel=33
    2, 2, 0, 10, -9, 0, -8, 8, 2,
    -- layer=1 filter=77 channel=34
    -2, -8, 1, -7, -3, 5, 3, 2, -6,
    -- layer=1 filter=77 channel=35
    -5, -3, 4, -8, -2, -7, 5, -6, -5,
    -- layer=1 filter=77 channel=36
    8, 4, 2, -11, -4, -2, -1, -10, 3,
    -- layer=1 filter=77 channel=37
    -6, 4, -6, 0, -3, 6, -3, -9, -9,
    -- layer=1 filter=77 channel=38
    -4, -5, 3, 2, -9, 3, 8, 4, 2,
    -- layer=1 filter=77 channel=39
    -8, -3, 5, 0, 7, -4, 3, -5, -4,
    -- layer=1 filter=77 channel=40
    -6, -5, 9, -1, 5, 1, 3, 4, -1,
    -- layer=1 filter=77 channel=41
    9, -9, -1, -3, 1, 0, 4, 6, 0,
    -- layer=1 filter=77 channel=42
    3, -6, -7, 0, 0, -13, -6, 6, 0,
    -- layer=1 filter=77 channel=43
    -12, 0, 3, -10, -7, -9, -9, -1, -3,
    -- layer=1 filter=77 channel=44
    -9, -2, -3, 2, -3, -5, -2, -11, -7,
    -- layer=1 filter=77 channel=45
    -4, 5, -1, 4, 6, -1, 0, 4, -6,
    -- layer=1 filter=77 channel=46
    -5, -4, 0, -1, 3, 0, -14, 5, 8,
    -- layer=1 filter=77 channel=47
    1, 5, -8, -5, -10, 4, -2, -10, -12,
    -- layer=1 filter=77 channel=48
    -5, -5, -11, 2, -12, 6, 0, 6, 2,
    -- layer=1 filter=77 channel=49
    -10, -13, 0, -12, -10, 6, -10, -6, 7,
    -- layer=1 filter=77 channel=50
    2, -3, -10, 0, 1, -4, 5, 8, 8,
    -- layer=1 filter=77 channel=51
    -8, 0, -4, -2, -5, 3, 0, 3, -2,
    -- layer=1 filter=77 channel=52
    7, -3, 1, 0, 5, -9, -2, 6, -8,
    -- layer=1 filter=77 channel=53
    -12, 0, -8, -6, 2, -6, 7, -10, -1,
    -- layer=1 filter=77 channel=54
    7, 0, 3, 0, 5, 3, 8, 1, 5,
    -- layer=1 filter=77 channel=55
    -7, -2, 1, -5, 9, 10, 12, 8, -2,
    -- layer=1 filter=77 channel=56
    6, -1, -6, 8, -10, 7, -6, 7, -1,
    -- layer=1 filter=77 channel=57
    -11, -4, -8, -4, 8, -10, -9, 6, -9,
    -- layer=1 filter=77 channel=58
    6, -7, 2, 6, -5, -4, 9, -2, 5,
    -- layer=1 filter=77 channel=59
    -2, -13, 2, 7, -3, 3, 6, 0, 8,
    -- layer=1 filter=77 channel=60
    -5, -3, 2, 6, -7, 7, -8, 0, -11,
    -- layer=1 filter=77 channel=61
    -8, 10, -8, 3, -4, -9, 6, -2, -3,
    -- layer=1 filter=77 channel=62
    8, 0, 0, 3, -4, 5, -7, 2, -1,
    -- layer=1 filter=77 channel=63
    7, -13, 7, 0, -3, -12, -10, 4, -9,
    -- layer=1 filter=77 channel=64
    -9, -8, 2, 0, -6, 3, 4, -3, 1,
    -- layer=1 filter=77 channel=65
    1, 5, 0, -8, -1, 4, -5, -3, -8,
    -- layer=1 filter=77 channel=66
    -7, 7, 2, 2, -5, 4, 3, -12, -8,
    -- layer=1 filter=77 channel=67
    -1, 3, 11, -5, -8, 1, 2, 0, -2,
    -- layer=1 filter=77 channel=68
    -11, -4, 5, -7, 1, 5, -11, 1, -11,
    -- layer=1 filter=77 channel=69
    6, -9, 12, -3, 5, 1, 3, 5, 4,
    -- layer=1 filter=77 channel=70
    8, -2, 8, -2, -3, -4, 0, 4, 8,
    -- layer=1 filter=77 channel=71
    -8, 0, -12, -9, -1, -6, -12, 5, 4,
    -- layer=1 filter=77 channel=72
    -1, -3, -11, 5, 0, -8, -7, 0, 0,
    -- layer=1 filter=77 channel=73
    -5, -11, -7, 2, 5, -12, 0, -11, 4,
    -- layer=1 filter=77 channel=74
    1, 6, -5, -3, -3, 3, -1, -5, 4,
    -- layer=1 filter=77 channel=75
    4, 0, 1, -3, -3, 10, -6, -7, -11,
    -- layer=1 filter=77 channel=76
    -5, 2, -7, 3, -8, -2, 2, -1, -9,
    -- layer=1 filter=77 channel=77
    -9, -8, -3, -7, -8, -3, 7, 2, -5,
    -- layer=1 filter=77 channel=78
    4, -1, -8, 0, -4, 5, 4, -10, 0,
    -- layer=1 filter=77 channel=79
    -4, 4, -10, 5, 0, -6, 9, -10, -11,
    -- layer=1 filter=77 channel=80
    -8, 4, 0, -8, 8, -3, -1, 8, 3,
    -- layer=1 filter=77 channel=81
    2, 3, -8, 0, 3, 4, 7, 1, -11,
    -- layer=1 filter=77 channel=82
    1, 7, 1, -1, -1, 0, -10, -8, 6,
    -- layer=1 filter=77 channel=83
    -11, -1, 5, 8, -2, -10, 8, 2, -2,
    -- layer=1 filter=77 channel=84
    4, 6, -5, 3, -8, -1, 3, -9, -5,
    -- layer=1 filter=77 channel=85
    4, -2, -13, 6, 8, 7, -9, -4, -1,
    -- layer=1 filter=77 channel=86
    -6, -11, -4, 6, 2, -9, 0, -4, -8,
    -- layer=1 filter=77 channel=87
    -7, -1, -5, 3, -10, 8, 5, -6, 2,
    -- layer=1 filter=77 channel=88
    -4, -10, 1, 2, 3, 6, -7, 3, 8,
    -- layer=1 filter=77 channel=89
    -2, 0, 6, -7, -8, -2, -6, -9, -2,
    -- layer=1 filter=77 channel=90
    -6, 1, -10, -8, -11, -7, 1, -7, -12,
    -- layer=1 filter=77 channel=91
    -2, 3, -10, 0, 5, -9, -4, -4, 0,
    -- layer=1 filter=77 channel=92
    -11, 6, 0, -2, -2, 1, -1, 7, -3,
    -- layer=1 filter=77 channel=93
    -8, -13, -12, -3, -7, 1, 1, 7, 7,
    -- layer=1 filter=77 channel=94
    -9, -4, -6, 7, 1, -3, 6, -3, 4,
    -- layer=1 filter=77 channel=95
    6, -3, -13, 1, -9, 1, -10, 5, 1,
    -- layer=1 filter=77 channel=96
    -8, 6, -6, 0, 3, 5, 0, -10, -11,
    -- layer=1 filter=77 channel=97
    6, 6, 4, -1, 4, -12, -9, 4, 6,
    -- layer=1 filter=77 channel=98
    3, 1, -13, 5, -3, -1, 4, -6, 7,
    -- layer=1 filter=77 channel=99
    -13, 1, 1, 5, 7, 3, -7, -6, -8,
    -- layer=1 filter=77 channel=100
    -10, 0, 5, 1, 5, -11, 0, -6, -4,
    -- layer=1 filter=77 channel=101
    0, 3, -4, -13, -4, -3, -12, -2, 6,
    -- layer=1 filter=77 channel=102
    -6, 0, -10, -7, -10, 0, -12, 0, -6,
    -- layer=1 filter=77 channel=103
    4, 8, -1, -3, 3, -1, -8, 2, 8,
    -- layer=1 filter=77 channel=104
    -8, -1, 3, 4, 3, 6, 3, -5, -9,
    -- layer=1 filter=77 channel=105
    3, 4, 0, 0, -7, -4, -11, 8, 5,
    -- layer=1 filter=77 channel=106
    -4, 7, 1, 2, -6, -4, -2, -6, 5,
    -- layer=1 filter=77 channel=107
    -9, 5, -7, 5, -5, 3, -2, 10, 7,
    -- layer=1 filter=77 channel=108
    -2, -1, 10, -6, 7, -6, 3, 1, -1,
    -- layer=1 filter=77 channel=109
    9, 10, -3, -11, 3, 9, -6, 6, 4,
    -- layer=1 filter=77 channel=110
    -10, 2, 4, 7, -4, 1, -1, -12, -3,
    -- layer=1 filter=77 channel=111
    -8, -9, 0, 3, -8, -2, 5, -12, 6,
    -- layer=1 filter=77 channel=112
    -6, -8, 2, 5, 7, -5, 5, 2, -5,
    -- layer=1 filter=77 channel=113
    -2, -2, 7, -9, -8, -1, -3, -2, -11,
    -- layer=1 filter=77 channel=114
    0, 10, 4, 12, 2, 1, -7, -11, 6,
    -- layer=1 filter=77 channel=115
    -5, -4, -12, -12, 8, -2, 6, 0, -5,
    -- layer=1 filter=77 channel=116
    5, -7, 3, 9, 1, -2, 6, -4, 4,
    -- layer=1 filter=77 channel=117
    -5, 8, -10, -12, -7, -3, -2, -4, -2,
    -- layer=1 filter=77 channel=118
    0, 5, 3, -12, -2, 1, -3, 6, 1,
    -- layer=1 filter=77 channel=119
    -9, -11, 3, 8, 0, -7, 8, 6, 4,
    -- layer=1 filter=77 channel=120
    1, -11, -3, -6, -6, 5, -11, -9, 0,
    -- layer=1 filter=77 channel=121
    -9, 6, -8, 7, 8, -9, -3, 9, 1,
    -- layer=1 filter=77 channel=122
    1, -9, 8, 4, -9, -5, 7, -1, -2,
    -- layer=1 filter=77 channel=123
    4, -8, 0, 3, -1, -9, -3, -7, 4,
    -- layer=1 filter=77 channel=124
    0, -4, 4, 0, -7, -6, -6, -8, -5,
    -- layer=1 filter=77 channel=125
    2, 7, 0, -10, -5, 1, -2, -8, 6,
    -- layer=1 filter=77 channel=126
    5, -10, 0, -2, -6, -9, 0, -5, -5,
    -- layer=1 filter=77 channel=127
    2, 2, 5, 8, 5, -1, 1, -11, 9,
    -- layer=1 filter=78 channel=0
    -3, -9, 0, -10, 10, 14, -11, -13, 12,
    -- layer=1 filter=78 channel=1
    -35, -6, -28, -6, -41, -5, -4, -26, -43,
    -- layer=1 filter=78 channel=2
    29, 16, -9, 37, -10, -5, 36, 4, 7,
    -- layer=1 filter=78 channel=3
    0, -1, -19, -7, 2, -11, -8, 7, -1,
    -- layer=1 filter=78 channel=4
    -5, -2, 5, 2, 3, 0, 0, 7, -2,
    -- layer=1 filter=78 channel=5
    -28, 0, -27, 8, -59, -38, -23, -57, -75,
    -- layer=1 filter=78 channel=6
    10, -13, 2, -1, 1, 8, 1, -15, 9,
    -- layer=1 filter=78 channel=7
    66, 48, 37, 49, 59, 20, 28, 99, 21,
    -- layer=1 filter=78 channel=8
    -22, -32, -43, -24, -66, -23, -7, -64, -69,
    -- layer=1 filter=78 channel=9
    -22, -52, 36, -6, 15, -53, 24, 14, -37,
    -- layer=1 filter=78 channel=10
    60, 27, 33, 14, 75, -2, 21, 76, 36,
    -- layer=1 filter=78 channel=11
    10, 13, -9, 0, 9, 0, 0, 2, 1,
    -- layer=1 filter=78 channel=12
    5, -40, -62, 6, -68, 6, -42, -6, 13,
    -- layer=1 filter=78 channel=13
    -6, -4, -5, -11, 0, 1, 5, -10, 20,
    -- layer=1 filter=78 channel=14
    18, -13, 45, -4, -7, -23, -50, 34, -31,
    -- layer=1 filter=78 channel=15
    33, -25, 18, 15, -46, 0, 23, -41, 9,
    -- layer=1 filter=78 channel=16
    -8, -17, -24, -7, -46, -28, -10, -47, -42,
    -- layer=1 filter=78 channel=17
    3, 12, -13, -17, -16, -3, -13, -21, -12,
    -- layer=1 filter=78 channel=18
    23, -15, -18, -13, -14, -45, -51, -44, -41,
    -- layer=1 filter=78 channel=19
    -41, -58, -19, -9, -64, -91, 5, -61, 43,
    -- layer=1 filter=78 channel=20
    -12, -3, -12, -12, -24, 5, -5, -10, 9,
    -- layer=1 filter=78 channel=21
    -15, 17, 11, -1, 1, 39, -13, 12, 14,
    -- layer=1 filter=78 channel=22
    3, 15, -20, -2, -32, -8, 18, -18, -4,
    -- layer=1 filter=78 channel=23
    73, 51, 52, 125, 59, 79, 46, 95, 64,
    -- layer=1 filter=78 channel=24
    -18, -7, 7, -31, 1, 7, -8, -43, 6,
    -- layer=1 filter=78 channel=25
    21, 26, 2, 23, 20, -4, 6, 63, 14,
    -- layer=1 filter=78 channel=26
    -14, -6, 0, -20, -43, -6, 11, -21, 3,
    -- layer=1 filter=78 channel=27
    -5, -22, 11, 2, -10, 23, -23, -6, 17,
    -- layer=1 filter=78 channel=28
    17, 27, 17, 12, 36, 13, -7, 68, 27,
    -- layer=1 filter=78 channel=29
    -11, -18, -11, -32, -21, -13, -35, -14, -17,
    -- layer=1 filter=78 channel=30
    -6, -34, -10, -33, -5, -110, -51, -53, -48,
    -- layer=1 filter=78 channel=31
    19, -33, -40, 20, -41, -40, -27, -18, -42,
    -- layer=1 filter=78 channel=32
    -14, 19, 19, -14, -18, 15, -5, -8, 11,
    -- layer=1 filter=78 channel=33
    0, -35, -33, 11, -10, -4, 20, 16, 17,
    -- layer=1 filter=78 channel=34
    42, 5, -4, -5, 15, 0, 9, 16, 23,
    -- layer=1 filter=78 channel=35
    0, -10, -8, -12, 0, -10, -11, 1, -3,
    -- layer=1 filter=78 channel=36
    11, 5, 0, 11, 11, 3, 2, -4, 22,
    -- layer=1 filter=78 channel=37
    -7, -12, -46, -4, -57, -60, -16, -76, -20,
    -- layer=1 filter=78 channel=38
    10, 0, 19, 6, 17, -3, 0, 10, 7,
    -- layer=1 filter=78 channel=39
    3, 9, 2, 3, -6, 15, -6, -2, 3,
    -- layer=1 filter=78 channel=40
    45, -4, -22, -6, -1, -68, -16, -10, -34,
    -- layer=1 filter=78 channel=41
    -4, -27, 27, -28, -2, 5, -14, 14, -5,
    -- layer=1 filter=78 channel=42
    30, 18, -10, 46, 4, 2, 24, 2, -3,
    -- layer=1 filter=78 channel=43
    -8, 10, -24, 31, -19, 2, 6, -26, -31,
    -- layer=1 filter=78 channel=44
    -9, 6, -3, -3, -29, 5, 24, -9, 3,
    -- layer=1 filter=78 channel=45
    -22, 15, -1, -21, -10, 26, 21, -23, 31,
    -- layer=1 filter=78 channel=46
    -28, -38, -53, 16, -80, -79, -24, -26, -7,
    -- layer=1 filter=78 channel=47
    95, 24, 61, 65, 20, 30, 37, 40, 38,
    -- layer=1 filter=78 channel=48
    -13, -23, 20, -14, 1, 19, -26, 7, 9,
    -- layer=1 filter=78 channel=49
    28, -15, -1, 0, 4, 6, 24, -7, 6,
    -- layer=1 filter=78 channel=50
    -9, -4, -5, 0, 5, -16, 10, 5, 12,
    -- layer=1 filter=78 channel=51
    4, 8, 22, -10, 14, -9, -7, 14, 12,
    -- layer=1 filter=78 channel=52
    13, -2, -1, 1, -5, -6, -7, 17, 10,
    -- layer=1 filter=78 channel=53
    -1, -20, -9, 10, -16, 1, -7, 3, -7,
    -- layer=1 filter=78 channel=54
    18, 1, -8, 25, -2, -43, -3, 10, 20,
    -- layer=1 filter=78 channel=55
    25, 0, 5, 9, 6, 19, 15, 7, 10,
    -- layer=1 filter=78 channel=56
    18, 8, 13, 0, 4, 13, 0, 1, -6,
    -- layer=1 filter=78 channel=57
    72, 22, 4, 21, 47, -5, 24, 48, 10,
    -- layer=1 filter=78 channel=58
    119, 40, 61, 98, 76, 54, 51, 80, 60,
    -- layer=1 filter=78 channel=59
    -9, -11, -2, 8, 0, 4, -8, 1, 3,
    -- layer=1 filter=78 channel=60
    2, 0, 6, -5, 11, 3, 1, -1, -5,
    -- layer=1 filter=78 channel=61
    5, 5, -12, 0, -4, 3, -6, 3, 3,
    -- layer=1 filter=78 channel=62
    -27, -12, -36, -16, -61, -35, -9, -67, -27,
    -- layer=1 filter=78 channel=63
    -9, -1, 12, -6, -4, -2, -12, -6, 11,
    -- layer=1 filter=78 channel=64
    -11, -8, -3, 0, -7, 17, -18, 0, 13,
    -- layer=1 filter=78 channel=65
    -20, -4, 25, -22, 18, 32, -17, 17, 15,
    -- layer=1 filter=78 channel=66
    0, -10, -5, -7, -3, 0, -20, -1, 15,
    -- layer=1 filter=78 channel=67
    -7, 2, 38, -1, -1, 39, 27, 15, 45,
    -- layer=1 filter=78 channel=68
    0, 29, 8, 0, 17, 14, 40, -3, 35,
    -- layer=1 filter=78 channel=69
    5, -2, -18, -7, -38, -4, 24, -38, 18,
    -- layer=1 filter=78 channel=70
    20, -17, 6, -6, -10, 16, -5, 4, 5,
    -- layer=1 filter=78 channel=71
    -2, 5, 19, 17, 8, 35, -12, 21, 14,
    -- layer=1 filter=78 channel=72
    -8, -25, -12, 8, -19, -108, 7, -50, -19,
    -- layer=1 filter=78 channel=73
    -7, -10, -6, 1, -7, 3, -8, 1, -6,
    -- layer=1 filter=78 channel=74
    -8, 18, 15, 11, 14, -6, 32, -13, 35,
    -- layer=1 filter=78 channel=75
    -2, -9, -2, 34, -66, -39, -96, -31, -53,
    -- layer=1 filter=78 channel=76
    -5, -7, 5, -14, -35, -18, 8, -21, 9,
    -- layer=1 filter=78 channel=77
    -27, -1, 12, -18, 12, 31, -25, -19, 18,
    -- layer=1 filter=78 channel=78
    -8, 1, -20, -11, 7, -15, -24, -2, -3,
    -- layer=1 filter=78 channel=79
    14, -2, -21, -5, -57, -4, 16, -33, -1,
    -- layer=1 filter=78 channel=80
    -5, 1, 1, 3, -7, 5, 6, 1, 5,
    -- layer=1 filter=78 channel=81
    -5, -20, 3, -16, 6, 22, 0, -17, 19,
    -- layer=1 filter=78 channel=82
    -25, -2, 17, -11, 10, 33, -6, -4, 11,
    -- layer=1 filter=78 channel=83
    2, -9, -23, -18, -25, -14, 18, -36, -5,
    -- layer=1 filter=78 channel=84
    -25, -43, -33, -27, -57, -65, -49, -70, -81,
    -- layer=1 filter=78 channel=85
    70, 30, 30, 76, 39, 43, 52, 49, 49,
    -- layer=1 filter=78 channel=86
    5, 8, -4, 17, 2, 4, -9, 7, -2,
    -- layer=1 filter=78 channel=87
    -1, -92, 7, 24, -49, -89, 11, -78, -8,
    -- layer=1 filter=78 channel=88
    19, -7, 28, 7, 7, 18, 3, -6, 23,
    -- layer=1 filter=78 channel=89
    -27, -6, 13, -13, -22, 19, -28, -21, 13,
    -- layer=1 filter=78 channel=90
    0, 27, 0, -7, 8, 29, 53, 2, 30,
    -- layer=1 filter=78 channel=91
    11, 5, 0, 2, -1, -9, -6, 13, 0,
    -- layer=1 filter=78 channel=92
    -2, -1, -9, -37, -36, -29, -29, -25, 24,
    -- layer=1 filter=78 channel=93
    -5, -2, 13, -12, -2, 34, -14, 6, 25,
    -- layer=1 filter=78 channel=94
    18, 6, 0, -11, 5, -8, -18, -3, -1,
    -- layer=1 filter=78 channel=95
    -20, -70, -10, -12, -60, -92, -58, -75, -64,
    -- layer=1 filter=78 channel=96
    7, -22, -11, -2, -13, -10, -11, 0, -18,
    -- layer=1 filter=78 channel=97
    -4, -4, 2, -7, 1, 23, 0, 0, 9,
    -- layer=1 filter=78 channel=98
    -9, 18, -21, -4, -18, -5, 23, -21, -33,
    -- layer=1 filter=78 channel=99
    47, 58, 47, 13, 122, 33, 58, 68, 68,
    -- layer=1 filter=78 channel=100
    6, 12, 2, -4, 10, -4, -4, 10, 5,
    -- layer=1 filter=78 channel=101
    2, -2, 15, 0, -13, 9, -16, 0, 7,
    -- layer=1 filter=78 channel=102
    -1, 1, 1, -23, 5, -9, -35, -5, -11,
    -- layer=1 filter=78 channel=103
    8, -1, 3, -4, 5, 21, -21, 0, 7,
    -- layer=1 filter=78 channel=104
    25, 1, 25, 73, 23, 46, 31, 10, 22,
    -- layer=1 filter=78 channel=105
    -9, -1, 7, -7, 11, 13, -6, -1, 17,
    -- layer=1 filter=78 channel=106
    -25, -27, 4, -22, -41, 1, -1, -34, 8,
    -- layer=1 filter=78 channel=107
    -3, 3, 4, 3, -12, 2, -11, 4, 4,
    -- layer=1 filter=78 channel=108
    -2, -17, 9, -5, -7, 29, 19, -5, 11,
    -- layer=1 filter=78 channel=109
    3, -9, -7, 6, 6, -3, 3, 9, -8,
    -- layer=1 filter=78 channel=110
    2, 5, 13, -10, 9, -6, -2, -4, 10,
    -- layer=1 filter=78 channel=111
    29, -47, -1, -35, 14, -81, -50, -38, -44,
    -- layer=1 filter=78 channel=112
    9, -55, 1, 0, -47, -20, -80, -33, -7,
    -- layer=1 filter=78 channel=113
    39, 9, -31, 29, -12, -21, 14, 1, -1,
    -- layer=1 filter=78 channel=114
    17, -17, 0, -13, -44, -38, 11, -42, -11,
    -- layer=1 filter=78 channel=115
    29, 2, 5, 5, 24, -17, 9, 26, 12,
    -- layer=1 filter=78 channel=116
    -11, -3, -3, 5, 0, -4, -8, -1, -10,
    -- layer=1 filter=78 channel=117
    23, -79, -8, -86, -37, -51, -53, -75, -35,
    -- layer=1 filter=78 channel=118
    -16, -20, -17, -19, -6, -70, -33, -70, -53,
    -- layer=1 filter=78 channel=119
    -4, 14, 20, -8, -8, 26, 0, 5, 7,
    -- layer=1 filter=78 channel=120
    1, -1, -2, 0, 0, 4, -5, 12, -2,
    -- layer=1 filter=78 channel=121
    -2, -42, 24, 32, 11, -23, -12, 3, -13,
    -- layer=1 filter=78 channel=122
    -4, 2, -7, 10, -7, 0, -3, -8, 6,
    -- layer=1 filter=78 channel=123
    10, -15, 27, 27, -2, -2, 9, 21, 23,
    -- layer=1 filter=78 channel=124
    1, -2, -9, 14, -10, 0, 2, -2, -9,
    -- layer=1 filter=78 channel=125
    41, 13, 20, 14, 29, 15, 28, 32, 5,
    -- layer=1 filter=78 channel=126
    -73, -24, -30, -26, -29, 6, -22, -87, -56,
    -- layer=1 filter=78 channel=127
    -4, -22, -19, -1, -31, -74, -50, -71, -64,
    -- layer=1 filter=79 channel=0
    1, -6, -7, -5, 4, -6, -1, 0, -3,
    -- layer=1 filter=79 channel=1
    -11, 6, -11, 7, -8, -7, -6, -6, -11,
    -- layer=1 filter=79 channel=2
    6, -10, 5, 4, -10, -7, -10, 3, 4,
    -- layer=1 filter=79 channel=3
    1, 3, -3, -2, 7, -6, -6, -5, 9,
    -- layer=1 filter=79 channel=4
    4, 6, -2, -1, 3, -12, 6, -9, 3,
    -- layer=1 filter=79 channel=5
    0, 3, -1, 0, -5, 3, -1, 7, 8,
    -- layer=1 filter=79 channel=6
    -9, -8, 5, -11, 2, 9, -5, 3, -1,
    -- layer=1 filter=79 channel=7
    -7, -7, -3, -8, -6, 5, -10, -5, -8,
    -- layer=1 filter=79 channel=8
    -11, -2, 1, -10, -9, 5, -6, -8, -5,
    -- layer=1 filter=79 channel=9
    -2, -11, -4, -9, -4, -11, -5, -11, 1,
    -- layer=1 filter=79 channel=10
    -1, -11, 2, -4, -2, -8, 4, -4, 1,
    -- layer=1 filter=79 channel=11
    -1, -8, 6, 8, -8, -4, 2, -1, -12,
    -- layer=1 filter=79 channel=12
    -4, -9, -6, 8, 10, -7, 8, 5, -8,
    -- layer=1 filter=79 channel=13
    -1, 2, -2, -9, 4, -6, 8, 4, 7,
    -- layer=1 filter=79 channel=14
    0, -3, -1, 6, -12, 10, 1, 0, 6,
    -- layer=1 filter=79 channel=15
    -2, -6, -9, -11, 3, 5, -3, 7, -9,
    -- layer=1 filter=79 channel=16
    5, -11, 7, 0, 4, -11, -2, 0, 7,
    -- layer=1 filter=79 channel=17
    8, 1, 0, 5, -8, -12, -1, 6, -12,
    -- layer=1 filter=79 channel=18
    2, -12, -10, -9, -3, -3, -6, 1, -8,
    -- layer=1 filter=79 channel=19
    8, -3, 0, 4, -5, 0, 8, 5, 4,
    -- layer=1 filter=79 channel=20
    5, 7, -3, -10, -11, 3, -5, 0, 3,
    -- layer=1 filter=79 channel=21
    -9, -8, 5, 3, 6, -4, 1, 1, 0,
    -- layer=1 filter=79 channel=22
    -6, 2, -4, 5, 9, -6, 1, -7, 0,
    -- layer=1 filter=79 channel=23
    2, -5, -5, 5, 8, 8, -5, -5, -6,
    -- layer=1 filter=79 channel=24
    -8, -12, -12, -2, -8, 8, -9, 7, -11,
    -- layer=1 filter=79 channel=25
    2, 4, 2, -6, 2, -2, -8, 3, 2,
    -- layer=1 filter=79 channel=26
    1, 1, -7, -3, -10, -4, -4, 0, 6,
    -- layer=1 filter=79 channel=27
    -2, -9, -1, -8, 6, -7, 5, 0, 2,
    -- layer=1 filter=79 channel=28
    -2, -3, -9, -8, -2, -8, -11, 7, 2,
    -- layer=1 filter=79 channel=29
    -6, 6, -3, 3, 2, -6, -1, -5, -4,
    -- layer=1 filter=79 channel=30
    -8, 0, -1, -3, 0, 9, -8, 7, 5,
    -- layer=1 filter=79 channel=31
    -1, 0, 7, -10, -11, -3, -8, -2, -4,
    -- layer=1 filter=79 channel=32
    -2, 2, 6, -8, 6, 2, -3, 9, -4,
    -- layer=1 filter=79 channel=33
    -2, -6, -9, 0, -3, 6, 10, 4, -12,
    -- layer=1 filter=79 channel=34
    5, -4, 4, -10, -9, 2, 1, 2, -2,
    -- layer=1 filter=79 channel=35
    -8, -11, -6, -11, -9, -6, 7, 8, 0,
    -- layer=1 filter=79 channel=36
    7, 7, 7, 7, -10, -9, -10, -10, -6,
    -- layer=1 filter=79 channel=37
    -2, 3, 6, -5, -11, 3, 10, -11, 4,
    -- layer=1 filter=79 channel=38
    -3, -2, 0, 4, -10, 9, -2, -1, 2,
    -- layer=1 filter=79 channel=39
    -8, -6, -11, 4, -5, 5, 4, 8, 7,
    -- layer=1 filter=79 channel=40
    4, -13, 3, 0, 3, -5, -6, 1, -12,
    -- layer=1 filter=79 channel=41
    2, 8, 7, -1, -1, 8, -5, -3, -11,
    -- layer=1 filter=79 channel=42
    2, 6, 5, -2, -7, -11, -3, 5, -3,
    -- layer=1 filter=79 channel=43
    0, 2, -8, 3, 7, -2, 1, -4, -11,
    -- layer=1 filter=79 channel=44
    -2, -4, 6, 0, -2, -10, -10, -6, -10,
    -- layer=1 filter=79 channel=45
    4, 4, -7, -1, 8, 2, 6, -5, 7,
    -- layer=1 filter=79 channel=46
    -10, -8, -4, 7, 1, -10, 1, 8, 1,
    -- layer=1 filter=79 channel=47
    11, -3, -7, 4, 8, -11, 5, 4, 4,
    -- layer=1 filter=79 channel=48
    -5, -3, 0, -6, -1, -9, 3, -5, 1,
    -- layer=1 filter=79 channel=49
    -3, -11, 1, -2, 9, -4, -3, -6, 6,
    -- layer=1 filter=79 channel=50
    1, 3, 2, 0, 0, -5, -8, 0, -3,
    -- layer=1 filter=79 channel=51
    4, -3, 7, -6, -8, 5, 3, 8, 10,
    -- layer=1 filter=79 channel=52
    2, 4, 6, -7, -4, 1, 5, 10, 8,
    -- layer=1 filter=79 channel=53
    -1, -6, -3, -3, -7, -11, 4, 3, -6,
    -- layer=1 filter=79 channel=54
    -3, 8, 4, -4, -8, -2, -10, 8, -8,
    -- layer=1 filter=79 channel=55
    -8, -2, 6, -1, -5, -8, 1, -3, -6,
    -- layer=1 filter=79 channel=56
    3, -7, -4, -5, -8, 1, -9, 0, 3,
    -- layer=1 filter=79 channel=57
    -12, 7, -7, -9, 2, -5, -3, -2, -4,
    -- layer=1 filter=79 channel=58
    3, 4, 7, -3, -5, 9, -1, -2, -5,
    -- layer=1 filter=79 channel=59
    -11, -4, 7, -3, -7, -2, 4, -3, -11,
    -- layer=1 filter=79 channel=60
    -8, -8, -1, 4, 5, 6, 0, 2, 0,
    -- layer=1 filter=79 channel=61
    -9, 0, -2, 6, 0, 6, 8, -10, 3,
    -- layer=1 filter=79 channel=62
    0, 1, 5, 2, -2, -3, -7, -3, -7,
    -- layer=1 filter=79 channel=63
    -11, 2, 4, -11, 4, 6, 6, 0, -4,
    -- layer=1 filter=79 channel=64
    5, -5, 0, 0, -7, 6, -3, -5, 5,
    -- layer=1 filter=79 channel=65
    5, -11, -9, -5, 0, 6, -6, -6, 1,
    -- layer=1 filter=79 channel=66
    0, 7, 4, 0, -3, -10, -3, -5, -11,
    -- layer=1 filter=79 channel=67
    4, -4, 2, -9, 0, 5, 0, -9, 9,
    -- layer=1 filter=79 channel=68
    -7, -11, -10, 2, 0, -6, -8, -7, 7,
    -- layer=1 filter=79 channel=69
    5, -5, -12, -3, -3, 1, -2, -7, -5,
    -- layer=1 filter=79 channel=70
    -5, -9, -2, 3, 0, 11, -9, -2, -7,
    -- layer=1 filter=79 channel=71
    3, 8, -3, -2, -8, -11, -2, -11, -3,
    -- layer=1 filter=79 channel=72
    3, -4, -12, 6, -2, -1, -5, -11, -3,
    -- layer=1 filter=79 channel=73
    1, 6, 0, -5, -7, -11, -6, -5, -9,
    -- layer=1 filter=79 channel=74
    3, -7, 3, -11, -2, 2, -9, -1, 0,
    -- layer=1 filter=79 channel=75
    1, -12, -1, -10, 0, 8, 8, -8, 0,
    -- layer=1 filter=79 channel=76
    5, 2, 1, -8, -4, -1, 4, -11, -12,
    -- layer=1 filter=79 channel=77
    3, -7, -9, 8, -1, 7, 8, 1, 8,
    -- layer=1 filter=79 channel=78
    -10, 4, -3, -6, -2, 1, 1, -5, 4,
    -- layer=1 filter=79 channel=79
    8, -7, -6, 0, -2, 4, 6, 5, -2,
    -- layer=1 filter=79 channel=80
    -7, -9, -3, 2, 2, 1, -8, 3, 9,
    -- layer=1 filter=79 channel=81
    -2, -11, 5, -4, -12, -8, -7, -2, 4,
    -- layer=1 filter=79 channel=82
    -1, 2, -11, -12, -6, 7, 9, 1, 6,
    -- layer=1 filter=79 channel=83
    -5, 1, -5, 7, 7, 5, -5, 3, -3,
    -- layer=1 filter=79 channel=84
    3, 2, 4, 4, 1, -8, -1, -11, -9,
    -- layer=1 filter=79 channel=85
    -2, -7, 6, 7, -8, 5, -9, 4, -10,
    -- layer=1 filter=79 channel=86
    4, 7, -7, -10, -11, -1, -2, 5, -9,
    -- layer=1 filter=79 channel=87
    4, 1, 1, 0, 6, -3, -2, 1, -4,
    -- layer=1 filter=79 channel=88
    -12, 0, -9, -8, 2, 4, -4, -1, 0,
    -- layer=1 filter=79 channel=89
    6, -7, -11, -7, 9, -5, -6, -2, 1,
    -- layer=1 filter=79 channel=90
    7, -7, 0, 6, -2, 2, 1, 9, 6,
    -- layer=1 filter=79 channel=91
    0, -1, 2, 7, 8, 3, -9, -5, -1,
    -- layer=1 filter=79 channel=92
    -5, -5, 8, -3, -6, -11, 2, -4, -8,
    -- layer=1 filter=79 channel=93
    3, 2, 4, -2, -1, 7, 5, 8, -2,
    -- layer=1 filter=79 channel=94
    3, -2, 4, -3, -8, 0, -2, -3, -5,
    -- layer=1 filter=79 channel=95
    5, 1, 0, 6, -9, 4, 6, -7, 0,
    -- layer=1 filter=79 channel=96
    -4, 0, -5, 3, 0, 1, -9, -9, -6,
    -- layer=1 filter=79 channel=97
    -7, -5, 8, -5, 0, -10, -9, -6, 4,
    -- layer=1 filter=79 channel=98
    -3, 3, 4, -4, 4, -11, 2, 3, 4,
    -- layer=1 filter=79 channel=99
    -4, -2, 2, -8, 0, 2, 6, 3, 0,
    -- layer=1 filter=79 channel=100
    -7, 7, 5, 1, -8, -7, -5, 2, -1,
    -- layer=1 filter=79 channel=101
    -5, -8, -3, 2, 6, -4, 5, -7, -1,
    -- layer=1 filter=79 channel=102
    -10, 3, 0, -9, -8, -12, -11, 8, 1,
    -- layer=1 filter=79 channel=103
    -1, -10, 0, -9, 3, -1, -9, 6, 6,
    -- layer=1 filter=79 channel=104
    4, 1, 0, -5, 2, 5, 6, 3, -6,
    -- layer=1 filter=79 channel=105
    0, -5, 2, 4, -6, 0, 2, 4, 4,
    -- layer=1 filter=79 channel=106
    4, -7, 11, 2, -7, -10, 6, 0, 9,
    -- layer=1 filter=79 channel=107
    -4, 3, 4, 2, -1, 4, 0, -3, 8,
    -- layer=1 filter=79 channel=108
    -4, -4, -11, 0, 1, -2, -11, -11, -2,
    -- layer=1 filter=79 channel=109
    -10, 1, 7, -12, -4, 7, 8, 1, -1,
    -- layer=1 filter=79 channel=110
    8, 0, -4, 4, 3, 5, -11, -9, 0,
    -- layer=1 filter=79 channel=111
    2, 6, 5, -1, 6, -2, -2, 6, 5,
    -- layer=1 filter=79 channel=112
    4, 5, -1, -4, 5, -2, -9, -8, -2,
    -- layer=1 filter=79 channel=113
    -5, -2, 11, 6, -6, 9, -7, -6, 4,
    -- layer=1 filter=79 channel=114
    -1, -3, 0, -2, -2, -3, -5, -4, -3,
    -- layer=1 filter=79 channel=115
    0, -3, -5, 0, 3, -7, 5, 8, -3,
    -- layer=1 filter=79 channel=116
    -4, -7, 4, -7, -6, 2, 1, 9, -7,
    -- layer=1 filter=79 channel=117
    -9, -7, 0, 1, 4, 0, -1, -8, 0,
    -- layer=1 filter=79 channel=118
    7, 5, 1, -3, -10, -8, 6, 0, 8,
    -- layer=1 filter=79 channel=119
    -1, 4, -2, 3, 1, -7, -4, 6, -9,
    -- layer=1 filter=79 channel=120
    1, 5, 2, 3, -2, 2, 3, -5, -7,
    -- layer=1 filter=79 channel=121
    0, -3, -1, 3, 6, -1, 4, -10, -8,
    -- layer=1 filter=79 channel=122
    -2, -3, -2, 0, 10, -8, 6, 0, 7,
    -- layer=1 filter=79 channel=123
    5, -4, -3, 3, -3, 1, 6, 0, 2,
    -- layer=1 filter=79 channel=124
    -2, 0, 0, -5, -11, -12, -6, -3, -6,
    -- layer=1 filter=79 channel=125
    8, 9, -1, 7, 8, 5, 8, 4, 4,
    -- layer=1 filter=79 channel=126
    6, 6, 4, 1, -6, -7, 3, 8, -7,
    -- layer=1 filter=79 channel=127
    -10, 0, -2, 2, 0, -12, 0, 0, 4,
    -- layer=1 filter=80 channel=0
    4, -14, -9, 2, 1, -8, -1, -9, -7,
    -- layer=1 filter=80 channel=1
    -7, -5, -1, 5, 5, 1, 1, 7, 0,
    -- layer=1 filter=80 channel=2
    -6, -6, 3, -6, -3, 8, 0, 10, 1,
    -- layer=1 filter=80 channel=3
    4, -4, -5, -1, -8, -8, -6, 0, 9,
    -- layer=1 filter=80 channel=4
    -7, -9, -11, 0, -7, 2, 6, -10, -12,
    -- layer=1 filter=80 channel=5
    -11, 0, -8, -1, -1, -1, 0, -8, 0,
    -- layer=1 filter=80 channel=6
    0, -3, 0, 1, -13, -1, -15, -2, 0,
    -- layer=1 filter=80 channel=7
    9, 6, 5, -12, 1, -4, -13, 3, 0,
    -- layer=1 filter=80 channel=8
    -7, 2, -10, 3, -4, -12, -2, 1, -7,
    -- layer=1 filter=80 channel=9
    -9, 8, 6, 15, 5, 7, 7, -7, 0,
    -- layer=1 filter=80 channel=10
    5, -8, 0, -11, 7, 8, -4, -3, -13,
    -- layer=1 filter=80 channel=11
    -13, -4, -13, -3, -8, -9, -1, 4, -19,
    -- layer=1 filter=80 channel=12
    4, 6, -6, -3, -6, 11, -9, 10, -9,
    -- layer=1 filter=80 channel=13
    -1, -13, -7, -12, -4, 1, 3, 2, -13,
    -- layer=1 filter=80 channel=14
    13, -9, -11, 6, -5, 8, -11, 4, -8,
    -- layer=1 filter=80 channel=15
    4, -7, -11, -2, 1, 4, 0, -7, -2,
    -- layer=1 filter=80 channel=16
    -3, 0, -14, 0, -6, -7, -5, -8, -14,
    -- layer=1 filter=80 channel=17
    -11, -5, -11, -3, -3, 6, -11, 0, 2,
    -- layer=1 filter=80 channel=18
    -12, -5, 0, 12, -10, 2, -17, -3, 1,
    -- layer=1 filter=80 channel=19
    0, -10, 6, -8, -1, -10, 4, -8, -3,
    -- layer=1 filter=80 channel=20
    -1, -13, 2, -1, -8, -10, -5, -10, -3,
    -- layer=1 filter=80 channel=21
    2, 1, -3, 3, 1, 4, -7, -4, -12,
    -- layer=1 filter=80 channel=22
    -1, 5, 0, -5, 3, -4, 1, -10, -1,
    -- layer=1 filter=80 channel=23
    -13, 1, 3, -13, 7, -7, -8, 5, -8,
    -- layer=1 filter=80 channel=24
    -7, -2, -5, -4, -7, -6, -5, -1, -9,
    -- layer=1 filter=80 channel=25
    -9, 6, -7, 0, 0, 3, 1, -4, -8,
    -- layer=1 filter=80 channel=26
    6, -2, 0, 3, -5, 6, 4, 0, -9,
    -- layer=1 filter=80 channel=27
    -1, -8, 7, 2, 3, 2, -8, 0, 2,
    -- layer=1 filter=80 channel=28
    -12, -11, 0, -11, 3, -13, 0, -5, -4,
    -- layer=1 filter=80 channel=29
    -4, -10, 8, 4, -11, 2, 0, 4, -5,
    -- layer=1 filter=80 channel=30
    3, 4, 2, 1, 0, -2, 1, -5, -12,
    -- layer=1 filter=80 channel=31
    -3, -10, 3, -7, 4, -3, 0, -12, 3,
    -- layer=1 filter=80 channel=32
    7, 6, -7, -6, -9, -9, 5, 2, 0,
    -- layer=1 filter=80 channel=33
    -4, 1, 1, 6, -4, 1, 8, 3, -12,
    -- layer=1 filter=80 channel=34
    0, 3, 0, 0, -6, -3, 6, -8, -10,
    -- layer=1 filter=80 channel=35
    6, -5, 0, -8, -4, 0, 4, -9, -1,
    -- layer=1 filter=80 channel=36
    2, 0, -14, -5, -18, -10, 3, -9, -7,
    -- layer=1 filter=80 channel=37
    -10, 9, 7, -7, 9, 1, -11, -3, -10,
    -- layer=1 filter=80 channel=38
    1, -12, -6, -1, -12, -11, -16, -4, -12,
    -- layer=1 filter=80 channel=39
    4, 0, 1, -13, 4, 3, -8, -4, -8,
    -- layer=1 filter=80 channel=40
    -7, -8, -9, -2, -9, -11, -7, -1, 0,
    -- layer=1 filter=80 channel=41
    4, -14, 3, 2, -9, -5, -1, -5, -6,
    -- layer=1 filter=80 channel=42
    5, 8, -3, 2, -6, 8, -12, 11, 0,
    -- layer=1 filter=80 channel=43
    -1, -3, -5, -1, -12, 0, 5, -9, -17,
    -- layer=1 filter=80 channel=44
    0, -2, 2, -6, -5, 9, -8, -4, -10,
    -- layer=1 filter=80 channel=45
    -1, -6, -12, -5, -9, 6, -4, -5, -3,
    -- layer=1 filter=80 channel=46
    13, -1, -9, 0, 4, 6, -10, 3, 2,
    -- layer=1 filter=80 channel=47
    -8, -11, -3, -10, 7, 6, -6, -2, -6,
    -- layer=1 filter=80 channel=48
    2, 1, 1, -14, -8, 1, -5, 0, 3,
    -- layer=1 filter=80 channel=49
    -1, 5, 2, 1, -5, 5, -8, -8, 9,
    -- layer=1 filter=80 channel=50
    -6, 2, 1, 8, 4, -8, -2, 1, -9,
    -- layer=1 filter=80 channel=51
    2, 7, -8, -1, -9, -4, -8, -2, 3,
    -- layer=1 filter=80 channel=52
    -5, 1, 1, 11, -9, 0, 6, 0, -6,
    -- layer=1 filter=80 channel=53
    0, -4, -8, 8, -9, -3, 2, -7, -1,
    -- layer=1 filter=80 channel=54
    -8, -4, 0, 8, -4, 2, -11, -6, 0,
    -- layer=1 filter=80 channel=55
    5, -14, -13, 0, -10, -13, 8, -14, -6,
    -- layer=1 filter=80 channel=56
    5, 3, -3, -9, -6, 0, 3, 6, 0,
    -- layer=1 filter=80 channel=57
    -11, 1, -3, 0, 3, -3, -7, -14, -11,
    -- layer=1 filter=80 channel=58
    -2, 1, 4, 0, 1, -3, -1, -15, 10,
    -- layer=1 filter=80 channel=59
    0, -4, 0, -2, -8, 5, 5, 0, -5,
    -- layer=1 filter=80 channel=60
    6, 1, 9, 7, -3, 9, 10, 2, 6,
    -- layer=1 filter=80 channel=61
    -5, 8, -3, 9, 0, -9, 7, -11, 7,
    -- layer=1 filter=80 channel=62
    -9, 4, 3, 12, 0, -5, -4, -6, -2,
    -- layer=1 filter=80 channel=63
    -12, 0, -11, -8, -6, -15, -10, 1, -11,
    -- layer=1 filter=80 channel=64
    -11, 1, -4, -6, -13, -9, -11, -8, -4,
    -- layer=1 filter=80 channel=65
    -6, -9, -3, -10, 2, 0, -1, -5, -11,
    -- layer=1 filter=80 channel=66
    -18, -16, 0, -7, -4, 1, -4, 0, -3,
    -- layer=1 filter=80 channel=67
    6, 1, -1, 12, 5, -9, 4, -3, 0,
    -- layer=1 filter=80 channel=68
    -4, -8, -10, 2, 0, 7, 9, -7, -6,
    -- layer=1 filter=80 channel=69
    -6, -3, 1, 4, 14, -8, -5, 0, -12,
    -- layer=1 filter=80 channel=70
    10, 7, -3, 1, 0, 3, 3, 8, 5,
    -- layer=1 filter=80 channel=71
    -12, 0, -6, -2, 2, 3, -11, 1, -12,
    -- layer=1 filter=80 channel=72
    -7, -10, -2, -10, 7, -11, -17, -4, 5,
    -- layer=1 filter=80 channel=73
    -1, 0, -8, 6, -7, 1, -1, 4, 5,
    -- layer=1 filter=80 channel=74
    -1, -4, 3, -11, -11, -5, -11, 8, -4,
    -- layer=1 filter=80 channel=75
    9, -8, 4, 10, 13, 3, -15, -12, -5,
    -- layer=1 filter=80 channel=76
    -4, -14, -10, -6, -3, -9, -10, -8, 6,
    -- layer=1 filter=80 channel=77
    1, -2, -7, 0, 3, 2, -11, 1, 0,
    -- layer=1 filter=80 channel=78
    -9, -9, 4, -8, 1, -10, 0, -8, 1,
    -- layer=1 filter=80 channel=79
    -7, -11, 0, -10, 11, -10, 3, -10, -14,
    -- layer=1 filter=80 channel=80
    -4, 9, 2, 6, 8, -5, -2, 1, 1,
    -- layer=1 filter=80 channel=81
    1, 1, -12, -11, -7, -1, -4, -6, -7,
    -- layer=1 filter=80 channel=82
    -10, -7, -2, -11, -5, 0, -2, 6, 5,
    -- layer=1 filter=80 channel=83
    -8, 4, -1, 5, 4, -2, 0, -6, -2,
    -- layer=1 filter=80 channel=84
    2, -1, 7, -4, -6, -8, -2, 0, 0,
    -- layer=1 filter=80 channel=85
    3, -10, -2, 0, 6, 9, 2, 0, 3,
    -- layer=1 filter=80 channel=86
    -2, -8, -17, -10, -12, -13, 7, -1, -6,
    -- layer=1 filter=80 channel=87
    7, 1, -8, 5, 1, 6, 8, 0, -5,
    -- layer=1 filter=80 channel=88
    -5, 3, -1, 0, -10, -9, -11, -9, -7,
    -- layer=1 filter=80 channel=89
    -5, -10, 3, 5, -10, -10, -13, 0, 0,
    -- layer=1 filter=80 channel=90
    7, -1, -14, 6, 0, -9, -8, -5, -5,
    -- layer=1 filter=80 channel=91
    0, 0, -1, -6, 0, -13, -12, 4, -11,
    -- layer=1 filter=80 channel=92
    10, -12, -7, 4, -5, -5, 5, 7, -8,
    -- layer=1 filter=80 channel=93
    -10, 0, 4, -7, 0, 0, 5, -2, -9,
    -- layer=1 filter=80 channel=94
    0, -15, 0, -8, 2, 0, -3, -3, -14,
    -- layer=1 filter=80 channel=95
    -6, -13, 6, 3, -12, -13, -2, -1, -4,
    -- layer=1 filter=80 channel=96
    -14, 5, 2, -11, -2, -13, 2, 0, -5,
    -- layer=1 filter=80 channel=97
    2, 0, 1, -3, -7, 2, -14, -16, -9,
    -- layer=1 filter=80 channel=98
    -3, 6, 0, 2, 2, -9, 0, -6, -19,
    -- layer=1 filter=80 channel=99
    6, 1, -12, -2, 8, 1, 4, -7, -4,
    -- layer=1 filter=80 channel=100
    2, 0, -11, -2, 2, -7, 0, -12, 2,
    -- layer=1 filter=80 channel=101
    0, 5, 4, -12, 2, 2, -4, 1, -3,
    -- layer=1 filter=80 channel=102
    0, -11, 6, 5, -8, 4, -8, -10, -2,
    -- layer=1 filter=80 channel=103
    -3, -16, -14, 3, -8, -18, 3, -11, -17,
    -- layer=1 filter=80 channel=104
    -11, 3, -1, 2, -9, -7, -13, -12, -4,
    -- layer=1 filter=80 channel=105
    -7, -13, 2, 6, -7, -8, 6, -2, 3,
    -- layer=1 filter=80 channel=106
    2, -9, -7, 4, -13, -8, 0, 8, -12,
    -- layer=1 filter=80 channel=107
    4, 8, 7, 0, -2, -8, -11, -3, 8,
    -- layer=1 filter=80 channel=108
    3, 3, -11, -7, -4, 7, -9, -2, -4,
    -- layer=1 filter=80 channel=109
    6, -4, 0, 6, 3, -1, 0, -3, -4,
    -- layer=1 filter=80 channel=110
    -9, -3, -3, -9, -3, 8, 8, 2, 5,
    -- layer=1 filter=80 channel=111
    0, -3, -9, 8, -10, -2, -1, -4, -7,
    -- layer=1 filter=80 channel=112
    -7, 4, 4, -7, 4, -2, 4, -10, -7,
    -- layer=1 filter=80 channel=113
    8, 0, 0, -3, -9, -14, -3, -10, -11,
    -- layer=1 filter=80 channel=114
    -3, -6, -6, 6, -2, 0, -10, -9, -1,
    -- layer=1 filter=80 channel=115
    2, 4, -8, 2, 1, 4, 0, 1, -9,
    -- layer=1 filter=80 channel=116
    0, -7, 4, 5, -7, 5, -8, 5, -8,
    -- layer=1 filter=80 channel=117
    7, 3, -1, -4, -6, -14, 0, 3, -3,
    -- layer=1 filter=80 channel=118
    7, 0, 2, 4, -6, -11, -5, -10, -11,
    -- layer=1 filter=80 channel=119
    0, 4, -3, -8, 6, -3, -10, -8, -9,
    -- layer=1 filter=80 channel=120
    -8, -1, -2, -4, -8, -10, 0, -12, -10,
    -- layer=1 filter=80 channel=121
    6, 2, -6, 2, -1, -13, -4, -15, -7,
    -- layer=1 filter=80 channel=122
    -4, 1, 7, 0, -5, -5, -8, 8, 6,
    -- layer=1 filter=80 channel=123
    2, -1, -4, -9, 3, -11, -3, 2, 0,
    -- layer=1 filter=80 channel=124
    0, -2, -8, 5, 0, -1, -7, -7, 0,
    -- layer=1 filter=80 channel=125
    15, -5, -11, -12, 0, -11, 11, 4, -4,
    -- layer=1 filter=80 channel=126
    1, 5, -12, 11, -1, -4, 0, 0, -7,
    -- layer=1 filter=80 channel=127
    -8, 3, 1, 6, -11, -11, -5, -3, -8,
    -- layer=1 filter=81 channel=0
    -9, -7, 1, -2, 0, -5, -5, -7, 5,
    -- layer=1 filter=81 channel=1
    -4, 5, -8, -10, 6, 2, -5, 0, -8,
    -- layer=1 filter=81 channel=2
    2, -10, -7, 0, -13, 2, -11, 4, 8,
    -- layer=1 filter=81 channel=3
    7, 0, -7, 5, 0, -8, 9, -4, -6,
    -- layer=1 filter=81 channel=4
    4, -2, 1, -8, -3, -1, -1, 2, 8,
    -- layer=1 filter=81 channel=5
    -2, 6, -6, 8, -1, -7, 4, -2, -7,
    -- layer=1 filter=81 channel=6
    12, 7, 7, 6, 0, 0, -7, -2, 5,
    -- layer=1 filter=81 channel=7
    9, -8, -6, -6, 0, -11, 8, 4, -1,
    -- layer=1 filter=81 channel=8
    -5, 7, 3, 7, 5, -6, 0, -3, -6,
    -- layer=1 filter=81 channel=9
    0, -5, 0, -3, -1, -11, -6, -5, 1,
    -- layer=1 filter=81 channel=10
    -12, -13, -7, -5, 6, -5, -11, -10, -8,
    -- layer=1 filter=81 channel=11
    -6, -10, 0, -3, 7, -8, 1, -3, 2,
    -- layer=1 filter=81 channel=12
    -4, -7, 7, -7, -4, -9, -4, 5, -5,
    -- layer=1 filter=81 channel=13
    -10, -4, -7, -6, -7, 0, -6, 4, -5,
    -- layer=1 filter=81 channel=14
    1, -1, -1, -9, 0, -10, 0, -6, 7,
    -- layer=1 filter=81 channel=15
    4, 4, 0, 4, -6, 6, -6, -11, 0,
    -- layer=1 filter=81 channel=16
    8, -8, 4, 3, -6, 0, 5, 3, 4,
    -- layer=1 filter=81 channel=17
    -4, 3, 7, -2, 5, -12, -11, 0, 7,
    -- layer=1 filter=81 channel=18
    0, 6, 1, -9, 2, 4, 8, -8, -11,
    -- layer=1 filter=81 channel=19
    0, -2, -7, 3, -10, 8, 1, 1, 4,
    -- layer=1 filter=81 channel=20
    5, 4, -10, 0, -5, -10, 1, 6, -3,
    -- layer=1 filter=81 channel=21
    0, -10, -7, -6, -2, 6, 7, -10, -9,
    -- layer=1 filter=81 channel=22
    -4, 9, -10, -4, 0, -4, -7, -7, -6,
    -- layer=1 filter=81 channel=23
    -1, -11, -1, -3, 0, 0, -3, -6, 7,
    -- layer=1 filter=81 channel=24
    -12, -7, -11, -11, -3, 0, 0, -9, -1,
    -- layer=1 filter=81 channel=25
    5, -11, -2, -11, -1, -1, 3, 9, -1,
    -- layer=1 filter=81 channel=26
    -4, -4, -2, 0, -4, 8, -8, 0, -12,
    -- layer=1 filter=81 channel=27
    0, 0, 9, 1, -4, -6, -5, 11, -1,
    -- layer=1 filter=81 channel=28
    -1, -11, -10, 7, 3, 4, -3, -10, 4,
    -- layer=1 filter=81 channel=29
    3, -12, 8, 5, 2, 7, -5, 3, 4,
    -- layer=1 filter=81 channel=30
    0, 5, -9, -3, 2, -8, 0, 4, 0,
    -- layer=1 filter=81 channel=31
    -9, 8, -5, 4, 0, 7, -4, 6, -8,
    -- layer=1 filter=81 channel=32
    -10, -10, -10, -1, 8, 6, -2, 0, 5,
    -- layer=1 filter=81 channel=33
    8, 1, 8, -7, -11, -3, 0, -6, -4,
    -- layer=1 filter=81 channel=34
    -5, 2, -9, -1, -10, 2, 8, -6, 1,
    -- layer=1 filter=81 channel=35
    -7, 2, -3, 4, -11, -10, -5, -12, -4,
    -- layer=1 filter=81 channel=36
    5, 5, -4, -7, -7, 6, 0, 6, -8,
    -- layer=1 filter=81 channel=37
    -6, 3, -4, -9, -5, 5, -6, -7, 7,
    -- layer=1 filter=81 channel=38
    -9, 0, -7, 5, -7, 5, 9, -3, 5,
    -- layer=1 filter=81 channel=39
    -12, 6, -9, 5, -10, 0, 5, 7, 0,
    -- layer=1 filter=81 channel=40
    -7, 5, -3, 0, 1, -10, -4, -11, -3,
    -- layer=1 filter=81 channel=41
    -6, -5, 2, -2, 2, -12, -3, -6, 3,
    -- layer=1 filter=81 channel=42
    -10, -5, 4, 1, 2, -9, 0, 0, -18,
    -- layer=1 filter=81 channel=43
    -5, -5, -9, -6, 7, 0, -10, -4, 7,
    -- layer=1 filter=81 channel=44
    -1, 0, -2, 0, 5, 6, 0, 5, -7,
    -- layer=1 filter=81 channel=45
    -5, -3, 1, 1, 1, -9, 5, 0, -5,
    -- layer=1 filter=81 channel=46
    -11, 5, 6, 5, -3, 7, -1, -7, -18,
    -- layer=1 filter=81 channel=47
    -2, 3, 0, 8, 4, 8, 4, -4, 1,
    -- layer=1 filter=81 channel=48
    4, 5, -2, -7, -3, -6, 2, -4, 0,
    -- layer=1 filter=81 channel=49
    -9, -5, -1, -12, 1, 0, 8, 3, 0,
    -- layer=1 filter=81 channel=50
    -1, -4, 0, 6, -3, -9, -7, 6, -9,
    -- layer=1 filter=81 channel=51
    -10, -10, -8, 4, -1, -11, -10, 8, 8,
    -- layer=1 filter=81 channel=52
    3, -7, 3, -5, 3, 0, 2, -3, -3,
    -- layer=1 filter=81 channel=53
    3, 1, -8, 0, 4, 0, -4, -9, 5,
    -- layer=1 filter=81 channel=54
    8, 2, 2, 4, -11, 6, -3, -12, -4,
    -- layer=1 filter=81 channel=55
    4, 7, 4, 2, -7, 3, 6, -13, -12,
    -- layer=1 filter=81 channel=56
    -10, -5, -3, -4, -10, 5, -7, 4, 8,
    -- layer=1 filter=81 channel=57
    -4, 5, -7, 0, -6, -6, 2, -10, 2,
    -- layer=1 filter=81 channel=58
    0, 0, 5, -12, 3, 6, -7, -1, 1,
    -- layer=1 filter=81 channel=59
    -6, -10, -12, 8, -10, -11, -3, 7, -6,
    -- layer=1 filter=81 channel=60
    -4, -3, -3, 2, 2, 5, -8, 0, 9,
    -- layer=1 filter=81 channel=61
    -1, -5, -6, -9, 0, 6, 1, 2, -9,
    -- layer=1 filter=81 channel=62
    -7, 7, -1, -6, -12, 3, -9, -5, 2,
    -- layer=1 filter=81 channel=63
    -7, -12, -13, 2, -9, -10, -4, -1, 4,
    -- layer=1 filter=81 channel=64
    0, -1, 3, 6, -4, 6, -11, -1, 5,
    -- layer=1 filter=81 channel=65
    -5, -4, -9, -4, 0, 2, 8, 8, 0,
    -- layer=1 filter=81 channel=66
    -7, -6, -5, 7, -12, -5, 2, -4, 2,
    -- layer=1 filter=81 channel=67
    -8, -9, -2, 0, -9, -9, -4, -3, 11,
    -- layer=1 filter=81 channel=68
    -11, -3, 9, -3, -2, -1, -1, 3, -5,
    -- layer=1 filter=81 channel=69
    -5, 0, -5, 3, -7, 5, 0, 0, -10,
    -- layer=1 filter=81 channel=70
    0, -5, 5, 0, 10, -7, -7, -6, 4,
    -- layer=1 filter=81 channel=71
    -10, 7, -5, -11, -2, 8, -6, -7, 0,
    -- layer=1 filter=81 channel=72
    -6, -6, 1, -3, -4, 6, 4, 7, 6,
    -- layer=1 filter=81 channel=73
    -4, 4, -1, -6, 2, 5, 2, -1, 0,
    -- layer=1 filter=81 channel=74
    -9, -6, -3, 3, 1, -12, -5, 3, 0,
    -- layer=1 filter=81 channel=75
    -6, -9, -11, -3, 0, 4, -10, -12, 10,
    -- layer=1 filter=81 channel=76
    2, -12, -4, 5, 4, 7, -8, -10, 4,
    -- layer=1 filter=81 channel=77
    0, 3, 3, 1, -4, 4, 6, -11, -2,
    -- layer=1 filter=81 channel=78
    -12, 2, -6, -12, 5, -1, 3, 4, 5,
    -- layer=1 filter=81 channel=79
    -4, -2, -2, -5, -11, 0, 2, -6, 0,
    -- layer=1 filter=81 channel=80
    -3, -1, -8, -2, 5, 8, -9, 4, -1,
    -- layer=1 filter=81 channel=81
    -1, 4, -2, -4, -6, -3, -4, 3, -2,
    -- layer=1 filter=81 channel=82
    0, -4, -12, -4, -3, -11, -8, 1, 5,
    -- layer=1 filter=81 channel=83
    4, 5, -8, 3, -13, 6, 0, 0, 4,
    -- layer=1 filter=81 channel=84
    5, -3, -9, -3, -11, -6, 2, -9, -5,
    -- layer=1 filter=81 channel=85
    5, 4, 8, -11, 7, -11, 5, 0, 3,
    -- layer=1 filter=81 channel=86
    -12, -13, -4, -4, -13, -9, 1, -5, -7,
    -- layer=1 filter=81 channel=87
    -1, 5, -3, -1, 8, -8, 6, -2, -10,
    -- layer=1 filter=81 channel=88
    -2, 9, 0, -6, -5, 0, -9, 1, 5,
    -- layer=1 filter=81 channel=89
    1, -10, -8, -5, -13, 0, -12, 4, -1,
    -- layer=1 filter=81 channel=90
    -12, 7, 3, 0, -9, 4, 8, -12, -5,
    -- layer=1 filter=81 channel=91
    2, 3, 4, 5, 0, 2, -6, -8, -10,
    -- layer=1 filter=81 channel=92
    -5, 5, -4, 5, 7, -12, 2, 0, -11,
    -- layer=1 filter=81 channel=93
    -4, 6, 1, 1, -4, -10, 2, 3, -12,
    -- layer=1 filter=81 channel=94
    -13, -5, 3, 1, 6, -9, 1, 5, -5,
    -- layer=1 filter=81 channel=95
    -1, -8, -11, -11, 7, -4, -7, -11, -10,
    -- layer=1 filter=81 channel=96
    7, 0, -3, 6, 2, 5, -2, -6, 2,
    -- layer=1 filter=81 channel=97
    -7, -6, 3, 5, -8, -10, -8, 7, -6,
    -- layer=1 filter=81 channel=98
    -2, -8, 5, -10, -9, 1, -3, -9, -8,
    -- layer=1 filter=81 channel=99
    -3, -10, -6, 0, -9, 0, -7, -5, -6,
    -- layer=1 filter=81 channel=100
    1, -11, -8, -2, 0, 5, 1, -12, -7,
    -- layer=1 filter=81 channel=101
    -1, 2, 1, 7, -8, 4, 0, -5, 3,
    -- layer=1 filter=81 channel=102
    4, 5, 0, 3, -10, 7, 4, -9, 0,
    -- layer=1 filter=81 channel=103
    -4, 8, 0, 1, -4, 4, -6, -10, -1,
    -- layer=1 filter=81 channel=104
    6, -7, -4, -1, -11, 4, 5, -7, -3,
    -- layer=1 filter=81 channel=105
    0, -12, -2, 3, -7, -7, -7, -5, 7,
    -- layer=1 filter=81 channel=106
    -8, -6, 3, 3, -4, -7, 11, 4, -7,
    -- layer=1 filter=81 channel=107
    3, -10, 1, -7, 7, 6, 6, 5, 3,
    -- layer=1 filter=81 channel=108
    -3, -7, 2, 1, -6, -5, -4, 4, 10,
    -- layer=1 filter=81 channel=109
    0, -7, -4, -3, 6, 0, -5, -9, -6,
    -- layer=1 filter=81 channel=110
    3, -1, 8, 0, 0, -5, -7, 7, -7,
    -- layer=1 filter=81 channel=111
    3, 4, -6, 5, 5, 7, 7, -1, -10,
    -- layer=1 filter=81 channel=112
    4, -5, -1, 7, -4, -7, -5, 1, -2,
    -- layer=1 filter=81 channel=113
    9, 5, 9, 7, 7, -8, -2, 7, 0,
    -- layer=1 filter=81 channel=114
    -4, -6, -1, 1, 5, -4, 8, -4, 2,
    -- layer=1 filter=81 channel=115
    -10, 5, -7, 7, 7, 4, 2, 8, 5,
    -- layer=1 filter=81 channel=116
    -2, 1, -9, -1, 3, -3, -1, -9, 1,
    -- layer=1 filter=81 channel=117
    4, 7, -7, 5, -10, -3, 0, -7, -3,
    -- layer=1 filter=81 channel=118
    6, -1, 2, 6, 0, 4, -10, -7, 0,
    -- layer=1 filter=81 channel=119
    3, 1, -5, 0, 2, 1, 4, -4, 2,
    -- layer=1 filter=81 channel=120
    -2, 2, 3, -13, -8, -6, -10, -4, 0,
    -- layer=1 filter=81 channel=121
    -10, 1, -2, 5, 6, 1, -6, 5, -4,
    -- layer=1 filter=81 channel=122
    0, -3, 7, -5, -4, -5, 7, 7, -4,
    -- layer=1 filter=81 channel=123
    1, -6, 4, -2, -9, 3, -3, -11, -10,
    -- layer=1 filter=81 channel=124
    -5, 7, 0, 2, -6, 5, -7, 3, -3,
    -- layer=1 filter=81 channel=125
    -4, -2, 3, 4, 11, 6, 3, -2, -8,
    -- layer=1 filter=81 channel=126
    -5, 2, -12, -7, -1, -5, 7, -10, -7,
    -- layer=1 filter=81 channel=127
    10, 10, 4, 0, -7, -6, 6, -12, 6,
    -- layer=1 filter=82 channel=0
    -32, -37, -34, -12, -16, -37, 24, 31, 18,
    -- layer=1 filter=82 channel=1
    -40, -49, -71, 20, 31, 4, 27, 17, 20,
    -- layer=1 filter=82 channel=2
    30, 24, 9, 37, 27, 6, 48, 19, 12,
    -- layer=1 filter=82 channel=3
    0, -1, -4, 10, -9, -2, 8, 3, 4,
    -- layer=1 filter=82 channel=4
    -8, -2, -14, -19, 6, 3, -1, -20, 0,
    -- layer=1 filter=82 channel=5
    -44, -43, -60, 45, 53, 37, 8, 32, 3,
    -- layer=1 filter=82 channel=6
    13, 8, 18, -21, -29, -5, -82, -55, -36,
    -- layer=1 filter=82 channel=7
    16, -74, -92, 56, -74, -82, 59, 19, -19,
    -- layer=1 filter=82 channel=8
    -39, -36, -57, 30, 34, 15, 25, 30, 21,
    -- layer=1 filter=82 channel=9
    -47, -34, -26, -60, -19, -15, -11, -7, 13,
    -- layer=1 filter=82 channel=10
    28, -65, -86, 60, -46, -34, 79, 13, -12,
    -- layer=1 filter=82 channel=11
    -6, -7, -2, 9, 6, 0, 10, 25, 26,
    -- layer=1 filter=82 channel=12
    44, -4, -32, -1, 3, -57, 43, 18, -26,
    -- layer=1 filter=82 channel=13
    -15, -1, 14, -27, -31, 18, -32, -8, 20,
    -- layer=1 filter=82 channel=14
    3, -67, -77, 5, -28, -82, 51, 28, -14,
    -- layer=1 filter=82 channel=15
    26, -38, -17, 37, -3, 59, -7, 3, 4,
    -- layer=1 filter=82 channel=16
    -63, -40, -63, 52, 42, 30, 22, 25, 0,
    -- layer=1 filter=82 channel=17
    -6, -35, -42, -22, -21, -32, 22, 20, 47,
    -- layer=1 filter=82 channel=18
    -43, -59, -52, -43, -43, -75, -8, -12, -17,
    -- layer=1 filter=82 channel=19
    -48, -83, -78, 84, 67, 84, 35, -33, -34,
    -- layer=1 filter=82 channel=20
    11, 12, 12, -3, -9, 20, -21, -17, -3,
    -- layer=1 filter=82 channel=21
    -8, -19, -5, -3, 3, -15, 20, 4, -4,
    -- layer=1 filter=82 channel=22
    -18, -8, 6, -12, -5, -16, 0, 13, 23,
    -- layer=1 filter=82 channel=23
    -23, -63, -49, 44, -18, 0, 81, 59, 60,
    -- layer=1 filter=82 channel=24
    -43, -22, -35, -7, 29, 25, 12, 28, 29,
    -- layer=1 filter=82 channel=25
    -12, -62, -106, 62, -4, -24, 50, 19, -11,
    -- layer=1 filter=82 channel=26
    -44, -59, -30, -2, -42, -16, 1, 8, 25,
    -- layer=1 filter=82 channel=27
    46, 46, 40, 26, 67, 58, 64, 65, 57,
    -- layer=1 filter=82 channel=28
    -13, -94, -116, 30, -35, -82, 57, 1, -5,
    -- layer=1 filter=82 channel=29
    -1, 18, 16, 11, 37, 38, 29, 32, 23,
    -- layer=1 filter=82 channel=30
    -60, -69, -55, -41, -36, -37, -14, -34, -65,
    -- layer=1 filter=82 channel=31
    22, 7, -18, 10, 27, -7, -7, 0, -27,
    -- layer=1 filter=82 channel=32
    -45, -91, -46, 3, -83, -22, 42, 4, 6,
    -- layer=1 filter=82 channel=33
    -12, -29, 6, 3, -5, 2, -5, -2, 22,
    -- layer=1 filter=82 channel=34
    -20, 0, 8, -6, -35, 21, -2, 1, 12,
    -- layer=1 filter=82 channel=35
    26, -7, 13, 22, 12, 27, 2, 13, 0,
    -- layer=1 filter=82 channel=36
    -20, -12, -23, -14, -4, -5, 32, 20, 19,
    -- layer=1 filter=82 channel=37
    -31, -28, -43, 73, 60, 47, 22, 10, -4,
    -- layer=1 filter=82 channel=38
    5, 22, 21, -13, 13, 22, -36, -20, -10,
    -- layer=1 filter=82 channel=39
    -15, 0, -16, -2, 8, 3, 24, 30, 14,
    -- layer=1 filter=82 channel=40
    12, -3, 25, -21, 32, -15, -41, -23, 5,
    -- layer=1 filter=82 channel=41
    -13, -41, -20, 33, -19, -34, 47, 2, 29,
    -- layer=1 filter=82 channel=42
    46, 25, 12, 45, 24, 17, 58, 48, 29,
    -- layer=1 filter=82 channel=43
    -56, -66, -71, 66, 46, 0, 40, 26, 17,
    -- layer=1 filter=82 channel=44
    -54, -88, -51, -4, -48, 4, 34, 24, 20,
    -- layer=1 filter=82 channel=45
    -52, -19, 1, -8, 35, 16, 4, 31, 10,
    -- layer=1 filter=82 channel=46
    -21, -24, 6, 99, 104, 144, 24, 18, -8,
    -- layer=1 filter=82 channel=47
    5, -42, 6, 32, 11, 1, 67, 22, 58,
    -- layer=1 filter=82 channel=48
    0, 16, 8, -21, -30, -17, 11, 11, -4,
    -- layer=1 filter=82 channel=49
    18, 13, 27, -6, -19, 16, 17, -9, 17,
    -- layer=1 filter=82 channel=50
    -4, -19, 9, -8, -25, -6, -10, -23, 2,
    -- layer=1 filter=82 channel=51
    38, 16, -16, 0, -18, -46, 25, -18, -33,
    -- layer=1 filter=82 channel=52
    -8, 8, -26, -8, 1, -32, 18, 5, -11,
    -- layer=1 filter=82 channel=53
    5, 7, 9, 6, 18, 19, 9, 13, 18,
    -- layer=1 filter=82 channel=54
    -8, -54, -88, 84, 33, 29, 53, 19, -36,
    -- layer=1 filter=82 channel=55
    7, 0, 5, 19, 13, 5, 28, 27, 36,
    -- layer=1 filter=82 channel=56
    -4, 0, 3, 9, -2, -5, -2, -4, 3,
    -- layer=1 filter=82 channel=57
    31, -36, -47, 29, -41, -33, 43, -9, -3,
    -- layer=1 filter=82 channel=58
    27, -58, -60, 71, -25, -16, 83, 14, 41,
    -- layer=1 filter=82 channel=59
    1, 1, 16, 14, -6, -5, -1, -2, -6,
    -- layer=1 filter=82 channel=60
    -5, 6, 20, 15, 6, 5, 8, -12, -14,
    -- layer=1 filter=82 channel=61
    2, -2, -5, 5, 0, -2, -5, 4, 3,
    -- layer=1 filter=82 channel=62
    -70, -50, -60, 53, 50, 17, 35, 44, 6,
    -- layer=1 filter=82 channel=63
    -21, -23, -5, 1, -8, -10, 20, 15, 12,
    -- layer=1 filter=82 channel=64
    -18, -9, -2, -34, -7, -29, 9, 0, 9,
    -- layer=1 filter=82 channel=65
    -2, 12, 0, -22, 27, -26, -10, 16, -1,
    -- layer=1 filter=82 channel=66
    -27, -23, -28, -6, -8, 3, 34, 29, 34,
    -- layer=1 filter=82 channel=67
    0, 68, 56, -51, 9, -11, -57, -23, -39,
    -- layer=1 filter=82 channel=68
    -87, -79, -31, -11, -46, -11, 16, 42, 21,
    -- layer=1 filter=82 channel=69
    -43, -94, -49, 23, 36, 29, -1, 31, 3,
    -- layer=1 filter=82 channel=70
    36, 39, 41, 19, 33, 40, -30, -24, 29,
    -- layer=1 filter=82 channel=71
    -14, -21, -46, 22, 41, 5, 37, 21, -4,
    -- layer=1 filter=82 channel=72
    -65, -75, -53, 16, -30, -3, 29, -45, -48,
    -- layer=1 filter=82 channel=73
    10, -19, 11, 0, -12, -8, 3, -7, -9,
    -- layer=1 filter=82 channel=74
    -85, -22, -2, -2, -4, -38, -30, 6, -7,
    -- layer=1 filter=82 channel=75
    -37, -66, -50, -30, -39, -58, -4, 36, -13,
    -- layer=1 filter=82 channel=76
    -50, -47, -37, 13, -53, -44, -8, 4, -8,
    -- layer=1 filter=82 channel=77
    -53, -30, -15, -31, 10, -24, 2, 39, -1,
    -- layer=1 filter=82 channel=78
    -57, -38, -59, 6, -18, -39, 28, 6, -31,
    -- layer=1 filter=82 channel=79
    -29, -57, -53, 54, 39, 24, 38, 32, 34,
    -- layer=1 filter=82 channel=80
    7, 7, 33, 31, -11, -3, 19, 36, -1,
    -- layer=1 filter=82 channel=81
    -47, -38, -42, 4, 0, -11, 34, 28, 27,
    -- layer=1 filter=82 channel=82
    5, 11, 0, -23, -4, -19, -7, 15, 4,
    -- layer=1 filter=82 channel=83
    -27, -88, -58, -3, -5, 18, 2, 31, 33,
    -- layer=1 filter=82 channel=84
    -84, -69, -20, -30, -85, -123, -38, -27, -45,
    -- layer=1 filter=82 channel=85
    -15, -49, -29, 38, -24, -11, 77, 16, 27,
    -- layer=1 filter=82 channel=86
    -20, -15, -18, -14, -3, 0, 14, 9, -6,
    -- layer=1 filter=82 channel=87
    -27, 0, -18, 37, 57, 63, 38, 0, 15,
    -- layer=1 filter=82 channel=88
    -5, 25, 12, -14, 2, -4, 7, 20, -4,
    -- layer=1 filter=82 channel=89
    -20, -1, 13, -40, -8, -23, -39, 13, -9,
    -- layer=1 filter=82 channel=90
    -80, -83, -61, -19, -28, 8, 14, 28, 35,
    -- layer=1 filter=82 channel=91
    36, 27, 12, -12, -21, -1, -24, -36, -15,
    -- layer=1 filter=82 channel=92
    -9, -67, -33, 8, -50, -4, 12, 21, 18,
    -- layer=1 filter=82 channel=93
    -24, -19, -24, -11, -2, -5, 16, 17, 12,
    -- layer=1 filter=82 channel=94
    -42, -43, -48, -9, -31, -36, 27, 35, -3,
    -- layer=1 filter=82 channel=95
    -81, -97, -49, -45, -66, -87, -43, -2, -34,
    -- layer=1 filter=82 channel=96
    -25, -34, -26, -6, -8, -22, 5, -24, -13,
    -- layer=1 filter=82 channel=97
    -33, -31, -36, -17, -4, -19, 38, 29, 19,
    -- layer=1 filter=82 channel=98
    -83, -72, -75, 21, 14, -8, 41, 37, 44,
    -- layer=1 filter=82 channel=99
    -31, -70, -84, -15, -12, -56, 55, 48, 16,
    -- layer=1 filter=82 channel=100
    -21, -1, 14, 10, 19, 24, 17, 30, 21,
    -- layer=1 filter=82 channel=101
    9, 21, 33, -24, -2, 0, -18, -22, -11,
    -- layer=1 filter=82 channel=102
    -25, -36, -61, -46, -25, -56, -6, 8, -40,
    -- layer=1 filter=82 channel=103
    -3, -4, 5, 21, 20, 13, 22, 36, 55,
    -- layer=1 filter=82 channel=104
    2, -18, -28, 0, -8, -23, 47, 35, 26,
    -- layer=1 filter=82 channel=105
    -18, -19, -35, -13, -10, -42, 29, 38, 32,
    -- layer=1 filter=82 channel=106
    -32, -3, 24, -26, -51, -6, -51, -17, 5,
    -- layer=1 filter=82 channel=107
    14, -5, 4, -8, -2, 5, 19, 22, 25,
    -- layer=1 filter=82 channel=108
    -47, -90, -36, -15, -47, 15, 21, 50, 44,
    -- layer=1 filter=82 channel=109
    -8, -9, 3, 0, -5, -3, 0, -9, -4,
    -- layer=1 filter=82 channel=110
    -13, -35, -21, -14, -32, -44, 6, 13, -13,
    -- layer=1 filter=82 channel=111
    -58, -55, -49, -62, -26, -97, -48, -12, -11,
    -- layer=1 filter=82 channel=112
    -39, -43, -7, -80, -98, -77, -40, -2, -7,
    -- layer=1 filter=82 channel=113
    24, -4, -6, 25, -9, 0, -3, 10, 18,
    -- layer=1 filter=82 channel=114
    5, -7, -17, 42, 59, 49, 16, 26, 6,
    -- layer=1 filter=82 channel=115
    -2, -18, -62, 28, -31, -39, 37, -2, -10,
    -- layer=1 filter=82 channel=116
    1, -9, 1, 5, -4, 1, 0, 3, -4,
    -- layer=1 filter=82 channel=117
    10, -40, -15, -79, -51, -32, 4, 16, 25,
    -- layer=1 filter=82 channel=118
    -82, -26, -33, -22, 3, -25, -24, -12, -23,
    -- layer=1 filter=82 channel=119
    -53, -105, -48, -17, -91, -40, 15, 7, 19,
    -- layer=1 filter=82 channel=120
    -4, -23, -14, 19, -1, -22, 19, -2, -10,
    -- layer=1 filter=82 channel=121
    -33, -41, -44, -6, 52, 67, 15, 57, 17,
    -- layer=1 filter=82 channel=122
    0, -7, -6, -2, -5, -4, -6, 5, 1,
    -- layer=1 filter=82 channel=123
    -9, -17, -35, 2, 19, 37, 39, 31, 13,
    -- layer=1 filter=82 channel=124
    15, 0, 14, 32, 16, 7, 1, -8, 0,
    -- layer=1 filter=82 channel=125
    58, 37, 44, -17, 21, 29, -20, -38, 14,
    -- layer=1 filter=82 channel=126
    -113, -68, -82, 17, 30, -16, 56, 52, 64,
    -- layer=1 filter=82 channel=127
    -71, -49, -26, -31, -11, -58, -19, -15, -38,
    -- layer=1 filter=83 channel=0
    3, 0, -4, 1, 5, -1, -1, 0, 7,
    -- layer=1 filter=83 channel=1
    -3, -11, -6, -4, 8, 0, 0, 3, 4,
    -- layer=1 filter=83 channel=2
    0, 0, -2, -21, 7, -9, -4, -2, -4,
    -- layer=1 filter=83 channel=3
    3, -4, 3, -2, -6, 9, 6, 6, 0,
    -- layer=1 filter=83 channel=4
    -10, 2, 8, -2, 0, -6, -3, 2, -9,
    -- layer=1 filter=83 channel=5
    -18, -6, 15, -3, -8, 11, -1, -15, -9,
    -- layer=1 filter=83 channel=6
    -1, -11, -12, -2, -14, -16, -10, -16, -9,
    -- layer=1 filter=83 channel=7
    -20, -8, -18, -8, 3, -13, -11, -5, 0,
    -- layer=1 filter=83 channel=8
    -9, 3, -11, -4, -6, -9, -4, -6, -16,
    -- layer=1 filter=83 channel=9
    -14, -12, 5, 10, 0, -13, 10, -12, 1,
    -- layer=1 filter=83 channel=10
    -4, -9, 0, -11, 1, 0, 2, -16, -8,
    -- layer=1 filter=83 channel=11
    -6, 0, -14, -2, 0, -4, -11, -3, -16,
    -- layer=1 filter=83 channel=12
    -20, -8, -3, 1, -8, 2, -10, -16, 0,
    -- layer=1 filter=83 channel=13
    -13, -4, -7, 2, -12, -13, 1, 0, -19,
    -- layer=1 filter=83 channel=14
    -3, -6, -7, 13, 5, 4, -4, -2, 18,
    -- layer=1 filter=83 channel=15
    -10, -7, 4, -1, -4, -8, -4, 11, -18,
    -- layer=1 filter=83 channel=16
    -3, -6, 12, 1, -8, 14, -2, -1, -9,
    -- layer=1 filter=83 channel=17
    -11, -11, -13, -2, 4, -4, -8, -12, -7,
    -- layer=1 filter=83 channel=18
    0, -10, -6, -4, 7, 5, -7, -1, 6,
    -- layer=1 filter=83 channel=19
    -9, 2, 0, 1, 7, -4, 4, -10, 0,
    -- layer=1 filter=83 channel=20
    -10, -7, -3, 0, -9, -6, -13, -4, -7,
    -- layer=1 filter=83 channel=21
    1, 0, -14, -14, 0, -12, -5, 0, -12,
    -- layer=1 filter=83 channel=22
    -6, -7, 4, 0, -14, -4, 1, 2, -15,
    -- layer=1 filter=83 channel=23
    -8, -12, 0, -5, 5, 0, -14, -12, -4,
    -- layer=1 filter=83 channel=24
    -6, 10, 0, -6, 3, -4, 0, 0, -15,
    -- layer=1 filter=83 channel=25
    -5, -2, 5, 9, 0, -17, 0, -15, -12,
    -- layer=1 filter=83 channel=26
    -14, 6, 3, -10, -1, -17, -4, 0, -13,
    -- layer=1 filter=83 channel=27
    -7, -5, 5, 1, -6, -7, 0, 2, -14,
    -- layer=1 filter=83 channel=28
    0, -10, -5, -3, -7, -10, 4, -5, -7,
    -- layer=1 filter=83 channel=29
    0, 3, 0, 6, 3, 0, 4, -2, -2,
    -- layer=1 filter=83 channel=30
    -13, -9, -10, 0, 6, -13, -8, -5, 1,
    -- layer=1 filter=83 channel=31
    -6, -4, 6, 7, -4, -13, -8, -4, 1,
    -- layer=1 filter=83 channel=32
    -8, 0, -9, 1, -7, 1, -11, 0, -18,
    -- layer=1 filter=83 channel=33
    -2, 8, 8, 3, -3, -2, 0, 5, -14,
    -- layer=1 filter=83 channel=34
    1, -6, -7, -9, 8, -2, -2, 1, -6,
    -- layer=1 filter=83 channel=35
    -6, 9, -1, -1, -10, 5, 6, -6, -2,
    -- layer=1 filter=83 channel=36
    -1, 0, -3, -6, 0, -8, -10, 3, 4,
    -- layer=1 filter=83 channel=37
    -13, -12, 0, 5, -3, -6, 2, -5, -12,
    -- layer=1 filter=83 channel=38
    -1, 0, -7, -14, -13, -9, -16, -5, -1,
    -- layer=1 filter=83 channel=39
    3, -7, 6, 5, -3, -12, 3, 4, 3,
    -- layer=1 filter=83 channel=40
    3, -1, -3, 11, -6, 2, -4, 0, 5,
    -- layer=1 filter=83 channel=41
    -9, -17, -2, -4, 6, -2, -18, 4, 0,
    -- layer=1 filter=83 channel=42
    -1, 0, 0, -14, -10, -11, -14, 2, 9,
    -- layer=1 filter=83 channel=43
    -9, -15, 1, -2, -7, 2, 6, -11, -14,
    -- layer=1 filter=83 channel=44
    -1, 0, 4, -5, 1, 2, -11, -4, 5,
    -- layer=1 filter=83 channel=45
    1, -9, 0, -4, 0, 0, -7, -7, -14,
    -- layer=1 filter=83 channel=46
    -19, -5, 16, 2, -17, -7, -3, -7, 4,
    -- layer=1 filter=83 channel=47
    0, -15, 2, -9, 2, -8, -2, 2, -17,
    -- layer=1 filter=83 channel=48
    -13, 2, -4, 7, -6, -11, -3, -1, -7,
    -- layer=1 filter=83 channel=49
    -13, -5, 6, 6, 2, -9, -13, -6, 2,
    -- layer=1 filter=83 channel=50
    -11, 6, -7, 4, -9, 5, 6, -5, -4,
    -- layer=1 filter=83 channel=51
    -4, -3, -7, -10, -3, 1, -10, -16, -6,
    -- layer=1 filter=83 channel=52
    1, -9, 5, 2, 8, -7, 0, 1, 0,
    -- layer=1 filter=83 channel=53
    -6, -5, -7, 5, 1, 0, -3, 8, 1,
    -- layer=1 filter=83 channel=54
    0, 3, -2, -2, -12, -8, -2, -12, -6,
    -- layer=1 filter=83 channel=55
    -8, 4, -2, -12, -3, -2, -11, -13, -15,
    -- layer=1 filter=83 channel=56
    -6, 7, 8, -4, -2, 5, -1, -3, -1,
    -- layer=1 filter=83 channel=57
    -12, -3, -12, -16, 0, 2, 0, -2, 3,
    -- layer=1 filter=83 channel=58
    -16, 5, -24, 7, 2, -1, -1, -8, -13,
    -- layer=1 filter=83 channel=59
    5, -6, 0, -6, -1, 1, -4, -5, -9,
    -- layer=1 filter=83 channel=60
    10, -6, 2, -9, 0, 0, 8, -6, 0,
    -- layer=1 filter=83 channel=61
    -1, 10, -4, -6, 12, 6, -3, -2, -6,
    -- layer=1 filter=83 channel=62
    -15, 0, 8, 2, 0, 5, 1, -14, -19,
    -- layer=1 filter=83 channel=63
    -8, -8, -10, -1, 5, -1, -8, -10, 2,
    -- layer=1 filter=83 channel=64
    -2, -2, -4, 5, -5, 5, 0, 1, 6,
    -- layer=1 filter=83 channel=65
    7, -9, -4, 4, -6, -1, 5, 0, 3,
    -- layer=1 filter=83 channel=66
    0, -12, -4, 3, -2, 0, -1, 4, -11,
    -- layer=1 filter=83 channel=67
    3, -4, -5, -10, -8, -8, -14, -2, -2,
    -- layer=1 filter=83 channel=68
    -14, 9, -3, -7, -12, -15, -13, 5, 9,
    -- layer=1 filter=83 channel=69
    -14, 1, 5, -9, -17, 0, -1, -8, -10,
    -- layer=1 filter=83 channel=70
    0, -2, -7, 2, 3, -16, -15, -1, -1,
    -- layer=1 filter=83 channel=71
    -12, -2, -4, -10, -18, -17, -7, -6, -18,
    -- layer=1 filter=83 channel=72
    5, 5, 3, 6, 0, -2, 6, -2, -7,
    -- layer=1 filter=83 channel=73
    2, 5, -11, -8, -9, 3, -9, 5, -6,
    -- layer=1 filter=83 channel=74
    -2, -6, 2, 9, -1, -14, 4, -1, -13,
    -- layer=1 filter=83 channel=75
    -5, -11, 3, -7, 7, -9, -1, -11, 17,
    -- layer=1 filter=83 channel=76
    -9, 0, 3, -6, -5, -9, -12, -3, -1,
    -- layer=1 filter=83 channel=77
    2, 0, 3, -2, 2, -7, -3, -9, 6,
    -- layer=1 filter=83 channel=78
    4, 6, -6, -3, 0, 1, 8, -9, -2,
    -- layer=1 filter=83 channel=79
    -19, 7, 1, 0, -2, -5, -6, -7, -5,
    -- layer=1 filter=83 channel=80
    -2, -4, -4, -6, 5, 3, -8, -7, -5,
    -- layer=1 filter=83 channel=81
    -4, -11, -9, -10, -10, 2, 2, -15, -12,
    -- layer=1 filter=83 channel=82
    -10, 0, -8, -7, -15, -2, -12, 0, -17,
    -- layer=1 filter=83 channel=83
    -11, -7, -4, 4, 2, -10, -1, -11, -12,
    -- layer=1 filter=83 channel=84
    -11, -5, -4, -1, 4, -9, -17, -17, 0,
    -- layer=1 filter=83 channel=85
    0, 0, -6, 7, -8, 1, 0, 0, -17,
    -- layer=1 filter=83 channel=86
    -11, -16, 2, 0, 0, -17, -11, 0, -7,
    -- layer=1 filter=83 channel=87
    2, 2, -10, -8, -8, -9, -10, -12, -12,
    -- layer=1 filter=83 channel=88
    -8, -3, -9, -2, -5, 6, -10, -19, 0,
    -- layer=1 filter=83 channel=89
    -5, -9, -11, -7, -12, -10, -10, -7, -12,
    -- layer=1 filter=83 channel=90
    0, -9, -8, 0, 1, -4, -1, -6, 7,
    -- layer=1 filter=83 channel=91
    -2, 2, -6, -11, 2, -5, -16, -16, -3,
    -- layer=1 filter=83 channel=92
    -10, 4, -5, -6, -7, -6, -13, -1, 0,
    -- layer=1 filter=83 channel=93
    -13, -1, -2, 0, -6, 0, -14, -11, -12,
    -- layer=1 filter=83 channel=94
    0, -4, -8, -11, 0, -10, 0, -5, -12,
    -- layer=1 filter=83 channel=95
    -10, -9, -14, 13, 2, -4, -7, -19, 4,
    -- layer=1 filter=83 channel=96
    0, 0, -12, -6, 2, 7, 0, -4, -5,
    -- layer=1 filter=83 channel=97
    -10, 4, -2, 1, -9, -7, -1, -13, -1,
    -- layer=1 filter=83 channel=98
    -4, -4, 0, 1, 2, 4, -5, -2, -14,
    -- layer=1 filter=83 channel=99
    10, -4, 0, 2, -11, 0, -6, -11, 1,
    -- layer=1 filter=83 channel=100
    -10, -14, -2, -9, -3, -7, 4, -2, -10,
    -- layer=1 filter=83 channel=101
    -5, -8, -10, 5, -12, 0, -1, -7, -7,
    -- layer=1 filter=83 channel=102
    6, 3, -2, -4, 0, 3, 6, -5, -1,
    -- layer=1 filter=83 channel=103
    -13, -5, -4, 0, 2, -9, -7, -11, -6,
    -- layer=1 filter=83 channel=104
    -5, -11, 1, -4, 0, -4, 7, -10, 0,
    -- layer=1 filter=83 channel=105
    5, -15, -2, 0, -2, -4, -6, -1, -9,
    -- layer=1 filter=83 channel=106
    -17, -5, 0, 5, -18, -16, 0, -7, -23,
    -- layer=1 filter=83 channel=107
    -3, 1, 4, -4, 9, 9, -8, -5, -5,
    -- layer=1 filter=83 channel=108
    -9, -3, -5, -23, -15, 0, -8, -7, -7,
    -- layer=1 filter=83 channel=109
    -3, 3, 5, -7, 10, -5, -6, 9, 3,
    -- layer=1 filter=83 channel=110
    -11, -7, 1, 0, -3, -10, 8, -11, -2,
    -- layer=1 filter=83 channel=111
    -16, -14, -9, -2, 6, 0, -3, -4, 2,
    -- layer=1 filter=83 channel=112
    -11, -11, 0, 0, -9, -12, -7, 1, -2,
    -- layer=1 filter=83 channel=113
    -5, 0, -10, -7, -5, 3, 1, 0, 5,
    -- layer=1 filter=83 channel=114
    -8, 4, 21, -17, 2, 4, 1, -4, -5,
    -- layer=1 filter=83 channel=115
    -1, 0, -3, -15, -15, -2, 2, -3, 1,
    -- layer=1 filter=83 channel=116
    3, -5, -6, -7, 8, -6, -7, -9, -6,
    -- layer=1 filter=83 channel=117
    -13, -13, -7, 2, 0, -2, -5, -6, 0,
    -- layer=1 filter=83 channel=118
    -9, -10, -5, 5, -2, -3, 1, -5, 0,
    -- layer=1 filter=83 channel=119
    -21, -6, -1, 5, 5, 0, -14, -14, -9,
    -- layer=1 filter=83 channel=120
    2, 2, 1, -11, -11, -18, -4, 0, -1,
    -- layer=1 filter=83 channel=121
    -14, -8, -11, 7, 6, -7, -2, -8, -3,
    -- layer=1 filter=83 channel=122
    -2, -7, -2, -7, 0, -2, -10, 10, -7,
    -- layer=1 filter=83 channel=123
    -16, -7, -10, -13, 0, -5, -12, -3, -3,
    -- layer=1 filter=83 channel=124
    -4, -7, 7, 0, -1, 0, -9, 0, -3,
    -- layer=1 filter=83 channel=125
    -14, -4, -12, -9, -20, -10, -7, -10, 0,
    -- layer=1 filter=83 channel=126
    -10, 8, -1, -6, -7, -2, 9, 4, -9,
    -- layer=1 filter=83 channel=127
    -11, -8, -3, 1, 5, -10, -2, -20, 8,
    -- layer=1 filter=84 channel=0
    -20, -20, -6, -8, 4, -13, 12, 2, -2,
    -- layer=1 filter=84 channel=1
    11, -5, -1, 14, 2, -1, 24, -16, 30,
    -- layer=1 filter=84 channel=2
    -9, -10, -27, -11, 0, 2, -33, -12, -24,
    -- layer=1 filter=84 channel=3
    -3, -3, -3, -3, 0, 0, -5, -3, -14,
    -- layer=1 filter=84 channel=4
    -11, 1, -9, -10, -6, -6, -4, -12, 4,
    -- layer=1 filter=84 channel=5
    4, 7, 16, 22, -26, -17, 12, -23, 22,
    -- layer=1 filter=84 channel=6
    -26, -26, -25, -10, -21, 3, -36, -22, -15,
    -- layer=1 filter=84 channel=7
    -5, 7, 6, -23, 11, 19, -6, 10, 0,
    -- layer=1 filter=84 channel=8
    10, 0, 5, 18, -1, -9, 26, -3, 33,
    -- layer=1 filter=84 channel=9
    -3, -4, 3, 3, 13, -15, 8, 16, 12,
    -- layer=1 filter=84 channel=10
    -8, 16, 2, -18, 12, 1, -4, 15, 0,
    -- layer=1 filter=84 channel=11
    -47, -48, -49, -42, -41, -43, -34, -43, -53,
    -- layer=1 filter=84 channel=12
    53, 12, 18, -28, -40, -12, 21, 24, 2,
    -- layer=1 filter=84 channel=13
    -8, -20, -16, -6, 7, 1, 13, 21, -1,
    -- layer=1 filter=84 channel=14
    14, 24, 2, -14, 7, 8, 18, 17, 3,
    -- layer=1 filter=84 channel=15
    8, -13, -6, 20, -12, -18, -12, -48, 22,
    -- layer=1 filter=84 channel=16
    19, 28, 8, 25, -3, -19, 6, 1, 35,
    -- layer=1 filter=84 channel=17
    -18, -18, -40, 3, -21, -12, 15, -1, -23,
    -- layer=1 filter=84 channel=18
    -31, -29, -22, -27, -25, -1, -10, -28, -17,
    -- layer=1 filter=84 channel=19
    14, 9, 8, 18, 18, 39, 5, 36, 16,
    -- layer=1 filter=84 channel=20
    -1, -9, -10, -6, 1, -12, 2, -3, 14,
    -- layer=1 filter=84 channel=21
    -7, -7, -1, -11, 16, 1, -3, 12, 0,
    -- layer=1 filter=84 channel=22
    -3, -16, -15, 2, 2, 0, 2, 6, 18,
    -- layer=1 filter=84 channel=23
    45, -11, 41, 0, -11, 11, -10, -14, -7,
    -- layer=1 filter=84 channel=24
    3, 10, -5, 5, -7, 13, 11, 27, 14,
    -- layer=1 filter=84 channel=25
    -7, 0, -7, 1, 11, -3, -1, 7, 21,
    -- layer=1 filter=84 channel=26
    -5, 0, -8, 12, 1, 11, 22, 19, 16,
    -- layer=1 filter=84 channel=27
    0, -4, 4, -9, -1, 1, -25, -23, -14,
    -- layer=1 filter=84 channel=28
    -8, 1, -8, -4, 28, 1, -13, 3, 1,
    -- layer=1 filter=84 channel=29
    -1, 17, 21, 0, 14, 5, -16, 0, 8,
    -- layer=1 filter=84 channel=30
    -7, -6, 6, 9, 0, 33, 7, 4, 7,
    -- layer=1 filter=84 channel=31
    -24, -24, -17, -11, -29, -23, 2, -25, -12,
    -- layer=1 filter=84 channel=32
    0, -22, 15, 5, 18, 9, 7, -2, 28,
    -- layer=1 filter=84 channel=33
    3, -5, -8, -11, 7, -10, -16, -3, 1,
    -- layer=1 filter=84 channel=34
    -59, -43, -7, -22, -13, -22, -33, -32, -14,
    -- layer=1 filter=84 channel=35
    2, 6, 19, 21, 3, 6, 18, 10, 15,
    -- layer=1 filter=84 channel=36
    -41, -41, -42, -61, -52, -54, -55, -34, -61,
    -- layer=1 filter=84 channel=37
    8, 24, 26, 1, -23, -24, -15, -15, 3,
    -- layer=1 filter=84 channel=38
    0, -1, -4, -1, -7, -8, 12, 8, -2,
    -- layer=1 filter=84 channel=39
    -20, -11, -17, -4, -10, -25, -21, -5, 0,
    -- layer=1 filter=84 channel=40
    -8, -13, -2, -14, -8, 0, -12, -26, -29,
    -- layer=1 filter=84 channel=41
    -4, -12, 13, 7, 17, 1, 4, 11, 25,
    -- layer=1 filter=84 channel=42
    -22, -9, -14, -23, -19, 5, -21, -20, -27,
    -- layer=1 filter=84 channel=43
    7, 11, 20, 14, 4, 8, 14, 0, 12,
    -- layer=1 filter=84 channel=44
    3, 7, -7, 1, 26, 9, 13, 15, 27,
    -- layer=1 filter=84 channel=45
    1, 16, -1, -4, -4, 6, 2, 9, 8,
    -- layer=1 filter=84 channel=46
    0, 11, -3, 15, -13, -6, -17, -30, 11,
    -- layer=1 filter=84 channel=47
    8, -25, 20, -18, -11, 11, -27, -1, 6,
    -- layer=1 filter=84 channel=48
    -9, -1, -4, 4, 0, -4, -7, 19, -1,
    -- layer=1 filter=84 channel=49
    -12, -6, 8, -15, 1, 4, -11, 11, 6,
    -- layer=1 filter=84 channel=50
    0, 4, 9, -14, -4, 0, 2, 4, 5,
    -- layer=1 filter=84 channel=51
    -15, -8, -2, -1, 10, 5, 8, 7, -2,
    -- layer=1 filter=84 channel=52
    1, 0, 16, -13, 1, 5, -15, 8, -1,
    -- layer=1 filter=84 channel=53
    6, 12, 15, 11, 8, 13, 16, 0, -2,
    -- layer=1 filter=84 channel=54
    -14, 37, 13, -7, 0, 4, -4, 15, 21,
    -- layer=1 filter=84 channel=55
    -20, -23, -11, -43, -46, -34, -51, -31, -45,
    -- layer=1 filter=84 channel=56
    -3, -2, -3, -10, -6, 4, 3, -5, 6,
    -- layer=1 filter=84 channel=57
    -18, -11, -9, -6, -8, 3, -10, 7, -19,
    -- layer=1 filter=84 channel=58
    13, 29, 15, 10, -7, 26, -31, 10, -15,
    -- layer=1 filter=84 channel=59
    7, 4, -1, 7, 7, -3, 4, 2, 13,
    -- layer=1 filter=84 channel=60
    0, -3, 0, -9, 0, 6, -11, -1, 0,
    -- layer=1 filter=84 channel=61
    7, 5, 8, 1, 14, 3, -7, -10, 1,
    -- layer=1 filter=84 channel=62
    1, 17, 11, 31, -13, -6, 8, 2, 28,
    -- layer=1 filter=84 channel=63
    -8, -8, -5, -12, 6, -1, -7, -20, -16,
    -- layer=1 filter=84 channel=64
    -13, -6, 6, 1, -1, -1, 1, -3, 8,
    -- layer=1 filter=84 channel=65
    -15, 8, -9, 9, 2, -10, 11, 13, 16,
    -- layer=1 filter=84 channel=66
    -1, -6, -2, -13, -5, -9, 0, -20, -7,
    -- layer=1 filter=84 channel=67
    -26, -23, -9, -27, -35, -41, -53, -32, -31,
    -- layer=1 filter=84 channel=68
    5, 5, -16, 3, 29, 17, 16, 34, 19,
    -- layer=1 filter=84 channel=69
    29, 12, 8, 23, -4, -2, 2, -10, 32,
    -- layer=1 filter=84 channel=70
    -39, -30, 3, -32, -49, -24, -55, -46, -14,
    -- layer=1 filter=84 channel=71
    7, 13, -5, -1, 0, 1, 4, 5, 14,
    -- layer=1 filter=84 channel=72
    -15, -29, -3, 13, -4, 27, 6, -11, 6,
    -- layer=1 filter=84 channel=73
    0, -3, 10, 10, 0, 0, 14, 8, 11,
    -- layer=1 filter=84 channel=74
    -3, -7, -15, -4, 7, 16, -4, 0, 1,
    -- layer=1 filter=84 channel=75
    6, 0, -6, 5, -5, 6, -1, 0, -4,
    -- layer=1 filter=84 channel=76
    -9, -4, -3, 14, 2, 14, 22, 14, 8,
    -- layer=1 filter=84 channel=77
    -8, 1, -11, 0, 4, 1, -7, 1, -4,
    -- layer=1 filter=84 channel=78
    -5, -13, -12, -12, 7, -5, -8, 10, 2,
    -- layer=1 filter=84 channel=79
    23, 24, 21, 16, -11, 11, 11, 12, 19,
    -- layer=1 filter=84 channel=80
    -6, 0, 7, 6, 4, -3, 0, 0, -6,
    -- layer=1 filter=84 channel=81
    -3, 4, 0, 5, 0, 5, -10, 13, -1,
    -- layer=1 filter=84 channel=82
    13, 5, -9, -2, 2, 7, 9, 15, 6,
    -- layer=1 filter=84 channel=83
    17, -12, 5, 24, 13, 13, 12, 18, 4,
    -- layer=1 filter=84 channel=84
    -11, -12, -9, 6, -4, 20, 10, -6, 4,
    -- layer=1 filter=84 channel=85
    -17, -12, 7, -8, -8, 14, -29, 1, 2,
    -- layer=1 filter=84 channel=86
    -30, -31, -22, -42, -37, -46, -23, -44, -22,
    -- layer=1 filter=84 channel=87
    2, -22, -2, -22, -9, -6, 3, 7, 12,
    -- layer=1 filter=84 channel=88
    -24, -18, -7, -15, -17, -6, -12, 0, -15,
    -- layer=1 filter=84 channel=89
    -7, -2, -5, 0, 19, 3, -2, 20, 13,
    -- layer=1 filter=84 channel=90
    2, -8, -18, 6, 3, 2, 20, 33, 16,
    -- layer=1 filter=84 channel=91
    -17, -3, -9, -11, -2, -2, -12, 1, 4,
    -- layer=1 filter=84 channel=92
    0, -24, -8, -12, 18, -9, -3, 23, 37,
    -- layer=1 filter=84 channel=93
    14, 2, 12, 1, 22, 0, 18, 13, 2,
    -- layer=1 filter=84 channel=94
    -2, -27, -18, -15, -7, -26, 0, -13, -17,
    -- layer=1 filter=84 channel=95
    -3, -2, 6, 2, 18, 34, 22, -6, 13,
    -- layer=1 filter=84 channel=96
    -19, -14, -1, 0, -3, -18, -2, -10, 0,
    -- layer=1 filter=84 channel=97
    -5, -6, 0, 5, 10, -5, 14, 13, 7,
    -- layer=1 filter=84 channel=98
    12, 8, 0, 19, 1, 0, 18, 4, 3,
    -- layer=1 filter=84 channel=99
    11, 26, 4, -26, 14, 0, 19, 6, -4,
    -- layer=1 filter=84 channel=100
    -12, -37, -26, -33, -26, -15, -9, -14, 2,
    -- layer=1 filter=84 channel=101
    0, -18, -8, 0, 1, -10, 5, 6, 9,
    -- layer=1 filter=84 channel=102
    -6, -11, -18, 2, -7, -17, 16, 6, -6,
    -- layer=1 filter=84 channel=103
    -30, -25, -18, -15, -25, -25, -27, -13, -26,
    -- layer=1 filter=84 channel=104
    14, -22, -2, 9, -29, -7, -3, -19, -12,
    -- layer=1 filter=84 channel=105
    -11, -10, -2, -12, -4, 7, 7, 14, -9,
    -- layer=1 filter=84 channel=106
    -12, -13, -9, -7, 0, 5, 6, 4, 14,
    -- layer=1 filter=84 channel=107
    -6, -6, -4, 6, 2, -6, -7, 7, 8,
    -- layer=1 filter=84 channel=108
    19, -12, 23, 15, 9, 30, 14, 7, 34,
    -- layer=1 filter=84 channel=109
    5, 4, 0, 3, -6, 3, 0, 7, -10,
    -- layer=1 filter=84 channel=110
    -10, 4, -9, -5, 1, 8, -1, 3, -5,
    -- layer=1 filter=84 channel=111
    6, 11, -8, 7, 6, 40, 26, -8, 15,
    -- layer=1 filter=84 channel=112
    27, 18, 25, 18, 14, 33, 25, 18, 1,
    -- layer=1 filter=84 channel=113
    -23, -26, -16, -3, 0, 4, -20, 2, 6,
    -- layer=1 filter=84 channel=114
    -1, 6, 12, -5, -40, -60, -32, -49, -10,
    -- layer=1 filter=84 channel=115
    -29, -16, -25, -36, -10, -34, -25, -10, -34,
    -- layer=1 filter=84 channel=116
    0, 7, -5, 13, -4, 3, 4, -1, 7,
    -- layer=1 filter=84 channel=117
    15, 27, 31, 24, 13, 23, 50, 22, 18,
    -- layer=1 filter=84 channel=118
    -2, -2, -6, 5, 10, 19, -3, 1, -5,
    -- layer=1 filter=84 channel=119
    2, 14, 0, 8, 16, 14, 20, 28, 12,
    -- layer=1 filter=84 channel=120
    -12, -3, 7, -5, 0, 1, 5, 5, 14,
    -- layer=1 filter=84 channel=121
    -16, -9, -30, -7, -10, 14, 1, -18, -13,
    -- layer=1 filter=84 channel=122
    0, 0, 1, -9, -7, -4, -3, 7, -9,
    -- layer=1 filter=84 channel=123
    -19, -29, -28, -39, -26, -9, -41, -37, -43,
    -- layer=1 filter=84 channel=124
    0, 6, -4, 2, 3, 1, 3, -10, -5,
    -- layer=1 filter=84 channel=125
    -26, -35, 3, -18, -22, -15, -28, -24, -23,
    -- layer=1 filter=84 channel=126
    19, 15, 17, 19, 10, 23, 38, 15, 13,
    -- layer=1 filter=84 channel=127
    -4, 0, -3, -6, 4, 12, 10, -6, 12,
    -- layer=1 filter=85 channel=0
    -9, -4, -8, -8, -8, 0, -5, 1, -1,
    -- layer=1 filter=85 channel=1
    -3, -3, 1, -9, -10, -7, -2, -5, -7,
    -- layer=1 filter=85 channel=2
    -1, 6, -12, -2, -13, -5, -5, -3, 3,
    -- layer=1 filter=85 channel=3
    3, 7, 7, 1, 0, -2, 4, 4, -4,
    -- layer=1 filter=85 channel=4
    7, -3, 0, -7, -10, -2, 1, 7, -10,
    -- layer=1 filter=85 channel=5
    -4, -27, 1, -15, -5, -11, -10, -2, 7,
    -- layer=1 filter=85 channel=6
    -3, -10, 1, -8, -9, -2, 4, 3, 0,
    -- layer=1 filter=85 channel=7
    -6, -4, -16, -13, -6, -6, 0, 2, -11,
    -- layer=1 filter=85 channel=8
    -10, -9, -7, 4, -2, -9, 1, -4, -5,
    -- layer=1 filter=85 channel=9
    -4, -10, -8, 10, 7, -2, -1, -5, 12,
    -- layer=1 filter=85 channel=10
    11, -12, -1, -6, -8, -15, -7, -2, -14,
    -- layer=1 filter=85 channel=11
    3, 0, -12, -9, -4, -15, -16, -2, -5,
    -- layer=1 filter=85 channel=12
    -20, -6, -17, 0, -2, -10, 4, 9, 3,
    -- layer=1 filter=85 channel=13
    -7, -3, -5, -8, -3, -2, -10, 7, -3,
    -- layer=1 filter=85 channel=14
    -2, -9, -5, 12, 1, -10, 3, 12, 0,
    -- layer=1 filter=85 channel=15
    -8, -3, 4, 3, -3, 4, 7, -3, 7,
    -- layer=1 filter=85 channel=16
    -6, -11, -11, -17, -2, -2, 2, 5, -10,
    -- layer=1 filter=85 channel=17
    0, -12, -3, 2, -4, 0, -4, -1, 3,
    -- layer=1 filter=85 channel=18
    4, -10, 5, 10, 0, -9, -20, 0, -12,
    -- layer=1 filter=85 channel=19
    5, 4, 4, 6, 0, -6, -4, 5, -12,
    -- layer=1 filter=85 channel=20
    -12, 0, -7, -14, -5, -3, 9, 0, -10,
    -- layer=1 filter=85 channel=21
    -8, 2, -11, -12, 4, -1, -5, -8, 4,
    -- layer=1 filter=85 channel=22
    -17, -8, -4, -1, -6, -9, 7, -1, 9,
    -- layer=1 filter=85 channel=23
    -1, 4, 0, -4, -2, 9, 0, 9, 0,
    -- layer=1 filter=85 channel=24
    -2, 3, 5, -2, -5, -1, 0, -9, -10,
    -- layer=1 filter=85 channel=25
    0, -6, -5, 1, -13, -17, 3, -14, 1,
    -- layer=1 filter=85 channel=26
    1, -22, 5, -8, -14, -18, -1, -7, -1,
    -- layer=1 filter=85 channel=27
    7, 3, -5, -2, 2, -1, 6, -8, 0,
    -- layer=1 filter=85 channel=28
    -7, 0, -9, 9, 4, -3, 3, -5, -11,
    -- layer=1 filter=85 channel=29
    6, -4, -5, 0, -12, 0, -7, 5, -3,
    -- layer=1 filter=85 channel=30
    0, 4, 10, 6, -7, -24, -1, 1, -13,
    -- layer=1 filter=85 channel=31
    4, -9, -7, -2, 3, 3, -1, -2, 0,
    -- layer=1 filter=85 channel=32
    -12, -2, -9, 4, 3, 0, -5, -2, -7,
    -- layer=1 filter=85 channel=33
    -6, -1, 3, 5, 1, -11, 3, 4, -2,
    -- layer=1 filter=85 channel=34
    -10, 4, -2, 7, -4, 2, 0, 1, -9,
    -- layer=1 filter=85 channel=35
    -8, -4, -8, -3, -2, -1, 0, 0, -3,
    -- layer=1 filter=85 channel=36
    -1, -6, 1, -1, 0, -7, 0, -4, -3,
    -- layer=1 filter=85 channel=37
    -11, -16, 1, -4, -12, -11, -9, -4, 0,
    -- layer=1 filter=85 channel=38
    -2, -15, -5, -1, -4, -4, 3, -3, -14,
    -- layer=1 filter=85 channel=39
    0, 9, 1, 2, 5, 7, -5, -11, 8,
    -- layer=1 filter=85 channel=40
    -4, 0, -7, -7, -10, -12, -3, -5, -1,
    -- layer=1 filter=85 channel=41
    4, -1, -9, -9, -1, 0, -3, -10, -7,
    -- layer=1 filter=85 channel=42
    0, -9, -8, -7, -3, -19, 14, 18, -2,
    -- layer=1 filter=85 channel=43
    -5, 0, -9, 5, -10, -2, 7, -4, -8,
    -- layer=1 filter=85 channel=44
    3, -14, 1, -10, -3, -12, 6, 0, 6,
    -- layer=1 filter=85 channel=45
    -3, 4, 5, -4, -14, 3, 2, 1, -7,
    -- layer=1 filter=85 channel=46
    10, -7, -4, -7, 3, 0, 19, 19, -1,
    -- layer=1 filter=85 channel=47
    -18, 7, -13, 0, -12, -7, -3, -3, 0,
    -- layer=1 filter=85 channel=48
    -10, 4, -2, -8, -5, 5, -3, 0, -10,
    -- layer=1 filter=85 channel=49
    -10, -10, -4, -2, 4, 8, -11, -14, 0,
    -- layer=1 filter=85 channel=50
    0, 2, 3, 9, -2, 5, 5, 8, 6,
    -- layer=1 filter=85 channel=51
    -10, 0, 5, 0, -4, 7, -5, -5, -1,
    -- layer=1 filter=85 channel=52
    10, -2, 3, -12, 9, 2, -5, -7, 4,
    -- layer=1 filter=85 channel=53
    0, -5, 1, -1, 6, -1, 1, -6, -5,
    -- layer=1 filter=85 channel=54
    16, 5, -11, 5, -3, -8, 5, -6, -8,
    -- layer=1 filter=85 channel=55
    0, 2, -5, 4, -12, 1, -9, -2, -3,
    -- layer=1 filter=85 channel=56
    7, 2, -7, -8, 4, -10, 9, 7, 3,
    -- layer=1 filter=85 channel=57
    -5, -9, -8, 7, 3, -16, 3, 0, -11,
    -- layer=1 filter=85 channel=58
    0, -9, -8, 2, 13, 1, -12, -2, -1,
    -- layer=1 filter=85 channel=59
    -4, -3, -6, 1, 5, 0, -7, -3, 6,
    -- layer=1 filter=85 channel=60
    5, 5, 0, 2, -7, -9, -3, -6, 0,
    -- layer=1 filter=85 channel=61
    -3, 9, -10, -8, -2, -8, 11, -6, 3,
    -- layer=1 filter=85 channel=62
    -9, -26, -4, -4, -20, -12, 6, 6, -4,
    -- layer=1 filter=85 channel=63
    -3, -1, 0, -10, -6, -4, -16, 1, -16,
    -- layer=1 filter=85 channel=64
    5, -8, 4, 1, -10, -4, 4, -9, 2,
    -- layer=1 filter=85 channel=65
    1, 2, 3, 4, 8, 2, -5, -8, -7,
    -- layer=1 filter=85 channel=66
    0, -2, -4, -7, 5, -11, -4, 1, -6,
    -- layer=1 filter=85 channel=67
    -2, 3, -7, -3, 3, -1, 0, -4, -2,
    -- layer=1 filter=85 channel=68
    -6, -2, -5, -4, -14, -15, 0, 0, -2,
    -- layer=1 filter=85 channel=69
    10, -9, -1, -8, -18, -2, 9, -12, -12,
    -- layer=1 filter=85 channel=70
    -5, -7, -13, 3, 2, 7, -14, -5, -11,
    -- layer=1 filter=85 channel=71
    -1, -2, -11, -5, -8, 5, 1, -6, -8,
    -- layer=1 filter=85 channel=72
    0, -1, 8, -6, 5, -8, 0, -12, 5,
    -- layer=1 filter=85 channel=73
    -9, -6, 5, -12, -9, -2, -4, -10, 0,
    -- layer=1 filter=85 channel=74
    1, -3, -5, 3, 8, -5, 4, -6, -8,
    -- layer=1 filter=85 channel=75
    0, 3, -17, -7, 0, -2, 4, 8, -6,
    -- layer=1 filter=85 channel=76
    -3, 3, -3, -4, -1, 4, 0, 8, 6,
    -- layer=1 filter=85 channel=77
    7, 2, -4, -9, 4, -3, -9, -6, 2,
    -- layer=1 filter=85 channel=78
    4, 0, -11, 6, 0, -8, 5, 4, 5,
    -- layer=1 filter=85 channel=79
    -6, -2, -4, 0, -14, 5, -6, -8, -6,
    -- layer=1 filter=85 channel=80
    12, 8, 0, -12, -5, 11, 6, 0, -8,
    -- layer=1 filter=85 channel=81
    -3, -8, -10, -11, 0, -6, 4, -2, 5,
    -- layer=1 filter=85 channel=82
    -8, -6, 5, -4, -1, 0, -13, 3, 0,
    -- layer=1 filter=85 channel=83
    -4, -11, -9, -6, 6, 1, 1, -10, 4,
    -- layer=1 filter=85 channel=84
    -13, -6, 6, 0, -5, -10, -3, -12, 0,
    -- layer=1 filter=85 channel=85
    3, -4, 7, 7, -10, 3, 1, -6, 0,
    -- layer=1 filter=85 channel=86
    -15, -17, 0, 0, -4, -15, -8, 0, -4,
    -- layer=1 filter=85 channel=87
    8, 4, 4, 3, -5, -4, 5, -2, -4,
    -- layer=1 filter=85 channel=88
    0, -7, -12, -4, 1, -8, -8, -1, -9,
    -- layer=1 filter=85 channel=89
    -2, 6, -3, -6, -10, -10, 0, -8, 2,
    -- layer=1 filter=85 channel=90
    0, -8, -7, -3, -5, 1, 2, -7, -6,
    -- layer=1 filter=85 channel=91
    -12, 4, -4, -15, -12, -8, -4, 0, -8,
    -- layer=1 filter=85 channel=92
    5, -10, -4, 6, 3, -4, -4, -2, 2,
    -- layer=1 filter=85 channel=93
    -2, -12, -9, -13, -11, 1, -3, -9, 2,
    -- layer=1 filter=85 channel=94
    -5, -4, 2, -10, 4, 2, 0, -11, -3,
    -- layer=1 filter=85 channel=95
    -11, -3, -1, -1, -7, -4, -9, -1, -4,
    -- layer=1 filter=85 channel=96
    -1, 8, -5, 1, 5, -6, -6, -7, 8,
    -- layer=1 filter=85 channel=97
    -9, -8, 6, 0, 0, 6, -10, -3, -9,
    -- layer=1 filter=85 channel=98
    -10, -18, -10, -4, -4, -3, -8, 5, -10,
    -- layer=1 filter=85 channel=99
    0, 8, -6, 0, -2, -3, -1, -7, 3,
    -- layer=1 filter=85 channel=100
    9, 8, 7, -8, -1, 0, -4, 2, -8,
    -- layer=1 filter=85 channel=101
    -8, -1, 2, -1, -3, -2, -3, 0, -1,
    -- layer=1 filter=85 channel=102
    -8, -9, -2, 0, -6, 5, -12, 8, 1,
    -- layer=1 filter=85 channel=103
    -12, -10, -7, -1, -6, 0, -12, -4, 1,
    -- layer=1 filter=85 channel=104
    0, 2, 6, -3, -9, 8, 3, 2, 6,
    -- layer=1 filter=85 channel=105
    -1, -4, -10, 0, 2, -14, -2, -12, 2,
    -- layer=1 filter=85 channel=106
    -18, -4, -15, -14, -9, -11, -16, -9, -18,
    -- layer=1 filter=85 channel=107
    -4, 1, 1, -4, 4, 2, 5, -11, -4,
    -- layer=1 filter=85 channel=108
    -8, -10, 4, -17, -14, -14, -6, -2, -16,
    -- layer=1 filter=85 channel=109
    -10, 9, 6, 1, 1, 6, 4, 8, -2,
    -- layer=1 filter=85 channel=110
    3, -7, -2, -2, 5, 0, 7, -4, -9,
    -- layer=1 filter=85 channel=111
    4, -8, 8, -3, 3, -15, -19, -7, -14,
    -- layer=1 filter=85 channel=112
    -6, -10, -8, 7, 5, 6, -1, 1, -2,
    -- layer=1 filter=85 channel=113
    4, -6, 7, -8, -3, 9, -12, 0, -9,
    -- layer=1 filter=85 channel=114
    -11, -16, -10, -7, -13, -3, 2, 3, -7,
    -- layer=1 filter=85 channel=115
    -10, -4, -10, -3, 0, 0, -2, -4, 0,
    -- layer=1 filter=85 channel=116
    6, 8, -1, 5, -5, 1, 7, 6, -2,
    -- layer=1 filter=85 channel=117
    -2, 5, -1, 3, -7, -1, -10, -12, -6,
    -- layer=1 filter=85 channel=118
    -10, -1, 3, -2, -11, 0, -13, -3, -2,
    -- layer=1 filter=85 channel=119
    -12, -15, 10, -15, 0, 0, -7, -10, -17,
    -- layer=1 filter=85 channel=120
    0, -9, 0, -15, -12, -10, -4, -9, 3,
    -- layer=1 filter=85 channel=121
    2, -3, -6, 8, 2, -3, 10, -7, 0,
    -- layer=1 filter=85 channel=122
    -5, 4, -7, 7, -7, 7, 10, -10, 0,
    -- layer=1 filter=85 channel=123
    -6, 9, 2, -7, -11, 0, -6, 1, -5,
    -- layer=1 filter=85 channel=124
    7, -3, 2, -5, -7, -5, -2, -1, 0,
    -- layer=1 filter=85 channel=125
    0, -4, -3, 1, -8, -7, -14, 0, -10,
    -- layer=1 filter=85 channel=126
    -12, 0, -3, 0, 2, 5, 1, 8, 4,
    -- layer=1 filter=85 channel=127
    8, -1, 6, -6, -9, -9, 1, 4, -13,
    -- layer=1 filter=86 channel=0
    -87, -83, -56, -64, -52, -47, -61, -53, -21,
    -- layer=1 filter=86 channel=1
    -6, -28, -14, -9, 0, -5, -38, -4, -24,
    -- layer=1 filter=86 channel=2
    49, 64, 50, 50, 38, 38, 31, 8, 29,
    -- layer=1 filter=86 channel=3
    5, 8, -3, -9, 1, 0, 8, 2, 8,
    -- layer=1 filter=86 channel=4
    64, 14, 59, -36, 10, -6, -15, -9, -26,
    -- layer=1 filter=86 channel=5
    -12, -21, -16, 23, 23, 11, -15, -31, -32,
    -- layer=1 filter=86 channel=6
    -6, -75, -56, -38, -26, -42, -41, -36, -42,
    -- layer=1 filter=86 channel=7
    -9, -6, -27, -18, 12, -28, -31, -11, 2,
    -- layer=1 filter=86 channel=8
    -8, -30, -18, 25, 14, 21, -15, -13, -15,
    -- layer=1 filter=86 channel=9
    94, 52, 48, 0, -36, -3, -40, -34, 4,
    -- layer=1 filter=86 channel=10
    -1, -2, -24, -10, 19, -7, -12, 3, -17,
    -- layer=1 filter=86 channel=11
    32, 5, 37, 17, 15, 26, 8, 20, 28,
    -- layer=1 filter=86 channel=12
    48, -23, -2, -14, -24, -36, 10, 3, 28,
    -- layer=1 filter=86 channel=13
    0, -42, -37, -46, -46, -28, -64, -25, -23,
    -- layer=1 filter=86 channel=14
    -6, 22, 4, -11, -13, -54, 0, 48, 15,
    -- layer=1 filter=86 channel=15
    -53, -40, 0, 4, 33, 11, -36, -62, -15,
    -- layer=1 filter=86 channel=16
    -3, -26, -37, 23, 12, 11, -23, -29, -28,
    -- layer=1 filter=86 channel=17
    -43, -44, -69, -81, -59, -52, -53, -27, -46,
    -- layer=1 filter=86 channel=18
    59, 25, 19, 6, 2, -26, -14, -27, 13,
    -- layer=1 filter=86 channel=19
    73, 59, 59, -20, -5, 21, -72, -63, -39,
    -- layer=1 filter=86 channel=20
    -66, -89, -98, -56, -48, -52, -67, -50, -64,
    -- layer=1 filter=86 channel=21
    0, 0, -7, 22, 27, 8, 18, 18, -9,
    -- layer=1 filter=86 channel=22
    -40, -62, -65, -1, -3, -23, -31, -32, -24,
    -- layer=1 filter=86 channel=23
    20, 22, 52, -13, 23, 14, -34, -33, -1,
    -- layer=1 filter=86 channel=24
    19, 26, 18, 11, 13, 38, 26, 3, 25,
    -- layer=1 filter=86 channel=25
    36, -10, 2, 8, 20, 12, -30, -4, -24,
    -- layer=1 filter=86 channel=26
    43, 9, 22, -13, -38, 8, -41, -21, 0,
    -- layer=1 filter=86 channel=27
    -35, -23, 0, -2, 6, 13, 0, 0, -4,
    -- layer=1 filter=86 channel=28
    3, -17, -5, 1, 0, -21, -5, 10, -13,
    -- layer=1 filter=86 channel=29
    -44, -42, -27, -36, -33, -14, -46, -39, -48,
    -- layer=1 filter=86 channel=30
    49, 6, 8, -30, -22, -71, -63, -58, -22,
    -- layer=1 filter=86 channel=31
    72, 43, 10, 42, 8, -18, 23, 33, 21,
    -- layer=1 filter=86 channel=32
    55, -10, 43, -14, -34, 28, -48, 26, 7,
    -- layer=1 filter=86 channel=33
    17, 20, 3, 11, 24, 3, 9, 17, 7,
    -- layer=1 filter=86 channel=34
    37, -26, -37, 48, -17, -23, 24, -12, 7,
    -- layer=1 filter=86 channel=35
    -1, 8, 0, -17, 8, -3, -4, -39, -3,
    -- layer=1 filter=86 channel=36
    1, -4, 24, -20, -3, 5, -3, -7, 7,
    -- layer=1 filter=86 channel=37
    0, -18, -16, 23, 24, 23, -20, -29, -23,
    -- layer=1 filter=86 channel=38
    -12, -16, -35, 4, -14, -2, -8, -25, -9,
    -- layer=1 filter=86 channel=39
    -45, -58, -42, -34, -24, -5, -27, -24, -16,
    -- layer=1 filter=86 channel=40
    3, -3, -26, -13, -15, -64, -35, -46, -39,
    -- layer=1 filter=86 channel=41
    64, 34, 35, -27, -31, 38, -40, 43, 39,
    -- layer=1 filter=86 channel=42
    25, 64, 42, 34, 45, 21, 31, 28, 28,
    -- layer=1 filter=86 channel=43
    6, -45, -27, 26, 5, 9, -31, -33, -17,
    -- layer=1 filter=86 channel=44
    23, -23, 21, -45, -21, 0, -56, -24, -2,
    -- layer=1 filter=86 channel=45
    -24, -12, -16, 2, 9, 7, -24, -33, -10,
    -- layer=1 filter=86 channel=46
    32, 23, 36, -7, -21, -19, -48, -53, -50,
    -- layer=1 filter=86 channel=47
    -11, 31, 1, 6, 16, 27, -29, 14, 4,
    -- layer=1 filter=86 channel=48
    -24, -46, -37, -15, -4, -13, -8, -7, -2,
    -- layer=1 filter=86 channel=49
    7, 11, -9, 16, 9, 18, 12, 7, 25,
    -- layer=1 filter=86 channel=50
    65, 11, 24, -12, -9, 16, -27, -14, -19,
    -- layer=1 filter=86 channel=51
    -15, -8, -29, 7, 8, -21, -11, 15, -20,
    -- layer=1 filter=86 channel=52
    8, 25, 26, -8, -1, 16, -17, -15, 5,
    -- layer=1 filter=86 channel=53
    -8, 0, -2, -8, -14, -7, -4, 5, 0,
    -- layer=1 filter=86 channel=54
    47, 9, 28, 43, 35, 37, -15, 0, -16,
    -- layer=1 filter=86 channel=55
    44, 44, 49, 45, 49, 60, 34, 45, 51,
    -- layer=1 filter=86 channel=56
    -5, -4, -3, -7, -6, 1, 2, 2, 9,
    -- layer=1 filter=86 channel=57
    -1, 16, -27, 10, 26, -21, 17, 16, -5,
    -- layer=1 filter=86 channel=58
    -5, 0, -18, -20, 17, 6, -35, -29, -18,
    -- layer=1 filter=86 channel=59
    31, 4, 15, -4, 18, 6, -14, 0, -26,
    -- layer=1 filter=86 channel=60
    -44, -27, 7, -65, -16, -30, -25, -7, 1,
    -- layer=1 filter=86 channel=61
    2, -10, 11, 1, -7, -4, -3, -7, 2,
    -- layer=1 filter=86 channel=62
    -1, -26, -30, 13, 0, 11, -35, -38, -38,
    -- layer=1 filter=86 channel=63
    9, -1, 9, -24, -32, -23, -24, -20, 11,
    -- layer=1 filter=86 channel=64
    -28, -29, -13, -45, -48, -43, -27, 4, -17,
    -- layer=1 filter=86 channel=65
    -44, -41, -34, -6, -26, -14, -9, -24, -24,
    -- layer=1 filter=86 channel=66
    -60, -35, -36, -49, -36, -40, -29, -21, -5,
    -- layer=1 filter=86 channel=67
    -20, -16, -24, 32, 31, 3, 12, 29, 2,
    -- layer=1 filter=86 channel=68
    28, -21, -1, -46, -33, 11, -48, -47, 1,
    -- layer=1 filter=86 channel=69
    -2, 0, 3, 33, 26, 45, -6, -18, 6,
    -- layer=1 filter=86 channel=70
    -22, -69, -112, 31, -10, -64, -36, -15, -26,
    -- layer=1 filter=86 channel=71
    9, 14, 23, 29, 15, 28, 22, 0, 7,
    -- layer=1 filter=86 channel=72
    87, 48, 55, 2, 10, -33, -30, -15, 16,
    -- layer=1 filter=86 channel=73
    -11, 13, -8, 27, 0, 24, -22, -11, -8,
    -- layer=1 filter=86 channel=74
    44, -4, 8, -48, 41, -48, -93, -49, 5,
    -- layer=1 filter=86 channel=75
    45, 27, 46, 4, -12, -50, -11, 11, 25,
    -- layer=1 filter=86 channel=76
    13, -54, -13, -46, -42, -19, -91, -47, -51,
    -- layer=1 filter=86 channel=77
    -12, -9, -25, -11, -6, 0, 1, 2, 1,
    -- layer=1 filter=86 channel=78
    -15, -41, -13, 3, -2, -15, 5, -24, -5,
    -- layer=1 filter=86 channel=79
    0, -38, -47, 22, 7, 2, -14, -36, -27,
    -- layer=1 filter=86 channel=80
    8, 18, 44, -5, 15, 23, 6, -14, 4,
    -- layer=1 filter=86 channel=81
    -16, 11, 4, 23, 18, 32, 7, 9, 6,
    -- layer=1 filter=86 channel=82
    -2, -13, -20, -9, 4, 6, 8, -5, -4,
    -- layer=1 filter=86 channel=83
    -52, -97, -36, -65, -32, -37, -63, -38, -54,
    -- layer=1 filter=86 channel=84
    66, -5, 23, -18, -36, -14, -67, -52, 6,
    -- layer=1 filter=86 channel=85
    22, 30, -8, -29, 5, 10, -39, -55, 23,
    -- layer=1 filter=86 channel=86
    0, 16, 17, 18, 17, 0, 3, 26, 20,
    -- layer=1 filter=86 channel=87
    77, 42, 26, 18, 6, 31, -36, -28, 2,
    -- layer=1 filter=86 channel=88
    6, 8, 2, 12, 16, 21, 23, 7, 11,
    -- layer=1 filter=86 channel=89
    -15, -33, -5, -14, -8, -5, -8, -1, 2,
    -- layer=1 filter=86 channel=90
    37, -14, 1, -20, -35, -12, -61, -35, -25,
    -- layer=1 filter=86 channel=91
    -41, -51, -79, -47, -23, -62, -56, -30, -42,
    -- layer=1 filter=86 channel=92
    35, -24, 49, -14, -28, 45, -31, 9, 31,
    -- layer=1 filter=86 channel=93
    -14, -4, -10, 4, 0, -7, 5, -4, -9,
    -- layer=1 filter=86 channel=94
    -94, -60, -57, -65, -68, -48, -69, -57, -39,
    -- layer=1 filter=86 channel=95
    36, -9, 9, -48, -6, -68, -76, -53, -11,
    -- layer=1 filter=86 channel=96
    -19, 11, -5, -14, -46, -2, -38, -29, -6,
    -- layer=1 filter=86 channel=97
    -81, -60, -77, -41, -51, -35, -32, -27, -28,
    -- layer=1 filter=86 channel=98
    -10, -29, -57, 23, 24, 20, -13, -7, -16,
    -- layer=1 filter=86 channel=99
    -44, -40, -4, -21, -17, -19, 23, 0, -11,
    -- layer=1 filter=86 channel=100
    7, -2, 27, -11, -34, -33, -22, 0, -8,
    -- layer=1 filter=86 channel=101
    -30, -68, -61, -47, -16, -48, -26, -22, -28,
    -- layer=1 filter=86 channel=102
    -93, -101, -89, -38, -37, -3, -74, -79, -61,
    -- layer=1 filter=86 channel=103
    44, 10, 12, -9, -3, -4, -4, -8, 11,
    -- layer=1 filter=86 channel=104
    62, 37, 17, -26, -31, 10, -44, -71, -2,
    -- layer=1 filter=86 channel=105
    -75, -73, -60, -52, -56, -26, -33, -42, -4,
    -- layer=1 filter=86 channel=106
    -1, -61, -25, -35, -42, -10, -54, -3, -11,
    -- layer=1 filter=86 channel=107
    -2, -16, -7, -9, 0, -6, -10, -3, -8,
    -- layer=1 filter=86 channel=108
    39, 3, 24, -8, -10, 4, -26, -13, -10,
    -- layer=1 filter=86 channel=109
    4, 8, 4, 7, 0, -10, -2, 1, -6,
    -- layer=1 filter=86 channel=110
    9, -31, -35, -13, -28, -11, -8, -16, 1,
    -- layer=1 filter=86 channel=111
    23, -17, -26, -59, -35, -53, -47, -88, -7,
    -- layer=1 filter=86 channel=112
    17, -44, -32, -56, -13, -8, -85, -47, 18,
    -- layer=1 filter=86 channel=113
    -23, -21, -18, 32, 23, -6, 20, -11, -28,
    -- layer=1 filter=86 channel=114
    -26, -26, -41, 36, 34, 23, -16, -10, 0,
    -- layer=1 filter=86 channel=115
    -24, -14, -25, -15, -11, -23, 4, -22, -6,
    -- layer=1 filter=86 channel=116
    1, 4, 5, 6, 5, -5, -7, -7, 7,
    -- layer=1 filter=86 channel=117
    -14, -25, -42, -42, 6, -14, -48, -46, 2,
    -- layer=1 filter=86 channel=118
    42, 0, 16, -27, -34, -48, -61, -80, 1,
    -- layer=1 filter=86 channel=119
    50, -6, 5, -29, -47, -4, -43, -1, -5,
    -- layer=1 filter=86 channel=120
    1, 6, -20, 25, 29, 12, -6, 8, -9,
    -- layer=1 filter=86 channel=121
    54, 59, 65, 16, 4, 7, 23, 18, 21,
    -- layer=1 filter=86 channel=122
    0, -5, 8, 5, -10, -9, -9, 4, -7,
    -- layer=1 filter=86 channel=123
    54, 61, 70, 39, 12, 13, 20, 30, 34,
    -- layer=1 filter=86 channel=124
    -13, -5, -1, -5, -3, -1, -12, -13, -6,
    -- layer=1 filter=86 channel=125
    -20, -69, -127, -49, -27, -73, -17, -49, -65,
    -- layer=1 filter=86 channel=126
    -23, -30, -58, 5, -10, -13, -50, -30, -40,
    -- layer=1 filter=86 channel=127
    33, 6, 9, -34, -3, -79, -63, -53, 6,
    -- layer=1 filter=87 channel=0
    -10, -6, 8, 0, 3, -3, 0, 0, -5,
    -- layer=1 filter=87 channel=1
    8, -9, 0, 2, 0, 1, -1, -4, -8,
    -- layer=1 filter=87 channel=2
    3, -4, -5, 2, -1, -7, 0, -9, 0,
    -- layer=1 filter=87 channel=3
    -4, 5, 9, 5, 3, -8, -1, 7, -6,
    -- layer=1 filter=87 channel=4
    -5, -4, 9, 2, -7, 7, 0, -4, -10,
    -- layer=1 filter=87 channel=5
    5, -10, -14, 4, -6, -1, -2, -9, -4,
    -- layer=1 filter=87 channel=6
    -5, 7, 3, -7, 0, -2, -3, 9, 1,
    -- layer=1 filter=87 channel=7
    -3, -2, -6, 5, -1, 5, -2, -10, -8,
    -- layer=1 filter=87 channel=8
    -5, 6, 5, -8, 4, 2, 2, 3, -6,
    -- layer=1 filter=87 channel=9
    -7, 0, -10, -5, 7, -10, -7, -2, 7,
    -- layer=1 filter=87 channel=10
    0, -7, -6, 6, 0, -1, -5, -9, -2,
    -- layer=1 filter=87 channel=11
    -2, 3, -1, 9, -6, -7, 3, -12, 4,
    -- layer=1 filter=87 channel=12
    -4, 0, -8, -4, -1, 0, -3, -8, 2,
    -- layer=1 filter=87 channel=13
    2, -2, 6, -4, -9, 1, -5, -2, 2,
    -- layer=1 filter=87 channel=14
    -2, -9, -6, -5, 3, -2, 9, -7, -5,
    -- layer=1 filter=87 channel=15
    0, 3, 2, -7, 0, 2, -1, 5, 4,
    -- layer=1 filter=87 channel=16
    -9, 0, -4, -10, 0, 10, -7, -1, 0,
    -- layer=1 filter=87 channel=17
    8, -4, 4, -8, 0, 1, 4, -9, -4,
    -- layer=1 filter=87 channel=18
    -8, -13, -3, -4, 6, 5, 6, -8, -4,
    -- layer=1 filter=87 channel=19
    -3, 8, 6, -1, 2, -2, 2, 8, 1,
    -- layer=1 filter=87 channel=20
    -9, -2, 7, 0, -1, -1, 0, -3, -4,
    -- layer=1 filter=87 channel=21
    6, 1, 5, 7, -6, -8, -4, 1, 9,
    -- layer=1 filter=87 channel=22
    -1, 6, -8, 6, 2, -8, -2, 0, 0,
    -- layer=1 filter=87 channel=23
    -6, 0, -7, -5, 3, -8, 8, -3, -8,
    -- layer=1 filter=87 channel=24
    6, -4, -4, -2, 4, -8, -10, -7, -1,
    -- layer=1 filter=87 channel=25
    0, -14, 1, 2, -6, -9, -13, 3, -6,
    -- layer=1 filter=87 channel=26
    -6, 1, -16, 2, 5, 3, -5, -9, 1,
    -- layer=1 filter=87 channel=27
    2, -10, 9, -10, -4, -7, -5, 0, -8,
    -- layer=1 filter=87 channel=28
    4, 1, -5, -8, 8, -4, 1, 0, 4,
    -- layer=1 filter=87 channel=29
    -1, 0, -11, 4, -1, 2, 5, 9, -1,
    -- layer=1 filter=87 channel=30
    2, -13, -3, -9, 4, -8, 8, 1, -11,
    -- layer=1 filter=87 channel=31
    -2, 1, 7, -8, -11, 2, -6, 8, 1,
    -- layer=1 filter=87 channel=32
    3, 6, 0, 2, 0, -3, -10, 9, -6,
    -- layer=1 filter=87 channel=33
    0, -6, 4, 1, 2, 3, 0, -3, 1,
    -- layer=1 filter=87 channel=34
    0, 2, -6, -7, -8, -7, -7, 6, -4,
    -- layer=1 filter=87 channel=35
    -3, 1, -10, 5, 4, 4, -2, -1, 2,
    -- layer=1 filter=87 channel=36
    0, 4, 8, -5, 3, 0, -5, -2, -3,
    -- layer=1 filter=87 channel=37
    8, 3, -8, 7, 0, -10, -3, 3, -7,
    -- layer=1 filter=87 channel=38
    -4, 2, 2, 1, 0, -10, -5, -10, 3,
    -- layer=1 filter=87 channel=39
    -7, -2, -2, 1, -8, 4, -9, -11, -10,
    -- layer=1 filter=87 channel=40
    -4, -8, 1, 0, -15, 1, 7, 1, -3,
    -- layer=1 filter=87 channel=41
    2, 0, -8, 0, -7, 7, -3, -5, -4,
    -- layer=1 filter=87 channel=42
    1, 4, 0, -18, -15, -3, -3, -15, -9,
    -- layer=1 filter=87 channel=43
    5, 5, -4, 0, -10, 7, 8, 7, -6,
    -- layer=1 filter=87 channel=44
    0, -6, 5, 7, -6, 0, 7, 0, -9,
    -- layer=1 filter=87 channel=45
    -1, -4, -1, -1, -7, 0, -11, -2, -11,
    -- layer=1 filter=87 channel=46
    -11, -8, -5, 7, 2, -5, -7, 9, 5,
    -- layer=1 filter=87 channel=47
    -8, 9, -9, 2, 3, 5, 2, 1, 0,
    -- layer=1 filter=87 channel=48
    6, -5, -3, 1, 3, 3, -1, 0, 1,
    -- layer=1 filter=87 channel=49
    0, 4, -2, -2, 0, -9, 0, -9, -2,
    -- layer=1 filter=87 channel=50
    1, -3, -9, 2, -10, 7, -7, 3, 4,
    -- layer=1 filter=87 channel=51
    -12, 0, -3, 3, -6, 2, -3, -9, -8,
    -- layer=1 filter=87 channel=52
    -5, 0, 8, -4, 7, -1, -7, -6, 0,
    -- layer=1 filter=87 channel=53
    -4, -5, 1, 1, 3, -4, -2, -4, -7,
    -- layer=1 filter=87 channel=54
    -6, -6, 6, 6, -5, 7, -6, 7, 7,
    -- layer=1 filter=87 channel=55
    -2, -4, -4, 1, 2, -13, -4, -3, -15,
    -- layer=1 filter=87 channel=56
    -10, -8, 7, -4, 7, -3, -1, -7, 1,
    -- layer=1 filter=87 channel=57
    -4, 4, -4, 8, -10, 1, -5, -2, -3,
    -- layer=1 filter=87 channel=58
    -8, -2, 5, 10, -9, -5, -3, -6, 3,
    -- layer=1 filter=87 channel=59
    1, 1, 2, -7, 7, 5, 3, 0, 7,
    -- layer=1 filter=87 channel=60
    9, 2, -4, 8, 8, -6, 9, -1, 1,
    -- layer=1 filter=87 channel=61
    -5, -1, -1, 2, 2, 1, 3, 0, -8,
    -- layer=1 filter=87 channel=62
    3, -2, -8, -4, 7, 5, -8, -5, 7,
    -- layer=1 filter=87 channel=63
    4, -5, 7, 0, 3, 2, 4, 6, -11,
    -- layer=1 filter=87 channel=64
    -6, 4, 2, -5, 7, -11, -3, -3, 6,
    -- layer=1 filter=87 channel=65
    -3, -1, 4, 1, 0, 8, 5, 4, -1,
    -- layer=1 filter=87 channel=66
    1, -1, -6, -8, 0, 0, -10, 1, -7,
    -- layer=1 filter=87 channel=67
    -8, -11, -10, 10, -7, -4, -7, -2, 1,
    -- layer=1 filter=87 channel=68
    8, -1, -10, -4, 1, -10, 1, 2, -10,
    -- layer=1 filter=87 channel=69
    0, -8, -17, 2, -6, -8, 4, -7, 6,
    -- layer=1 filter=87 channel=70
    -4, -4, -6, 8, -8, 9, 4, 8, 6,
    -- layer=1 filter=87 channel=71
    2, 7, 6, -9, 0, -2, -9, 7, 5,
    -- layer=1 filter=87 channel=72
    0, 6, 6, -1, 1, -1, 0, -2, -6,
    -- layer=1 filter=87 channel=73
    4, -3, -5, -4, -8, 3, -10, 8, 2,
    -- layer=1 filter=87 channel=74
    2, -2, 0, -6, -8, -2, 1, -2, 3,
    -- layer=1 filter=87 channel=75
    -11, -8, 8, 2, 4, -9, -2, -1, -7,
    -- layer=1 filter=87 channel=76
    -3, 7, 0, 2, 2, -2, -10, -2, 6,
    -- layer=1 filter=87 channel=77
    5, 0, 1, -8, 6, 2, 8, -4, -10,
    -- layer=1 filter=87 channel=78
    1, -10, -5, -1, 1, 3, -1, -9, 3,
    -- layer=1 filter=87 channel=79
    9, -10, -4, 7, 0, -10, 4, -4, -10,
    -- layer=1 filter=87 channel=80
    -10, 1, -9, 0, -3, 5, 8, -4, 1,
    -- layer=1 filter=87 channel=81
    -3, 2, -11, -8, 8, -10, 2, -8, -2,
    -- layer=1 filter=87 channel=82
    -4, 6, 0, 0, -8, 6, 8, -1, -6,
    -- layer=1 filter=87 channel=83
    2, 1, 3, 3, 4, -10, -10, -2, 7,
    -- layer=1 filter=87 channel=84
    8, 7, -5, 6, 6, -4, -10, 7, -9,
    -- layer=1 filter=87 channel=85
    -6, -3, 0, 0, 7, -9, 9, -5, -10,
    -- layer=1 filter=87 channel=86
    6, 7, -2, 1, 8, -3, 5, -11, -12,
    -- layer=1 filter=87 channel=87
    -7, -5, 2, 2, 1, 3, 3, 5, 0,
    -- layer=1 filter=87 channel=88
    -4, 2, 7, 7, 4, 9, 6, -6, -5,
    -- layer=1 filter=87 channel=89
    4, 0, 0, 0, 2, 6, -6, -11, 7,
    -- layer=1 filter=87 channel=90
    -3, 0, -5, 5, -11, -9, -3, -9, -9,
    -- layer=1 filter=87 channel=91
    -7, -5, -8, -3, -4, 0, -9, 9, 2,
    -- layer=1 filter=87 channel=92
    -11, -3, 1, 8, -10, 2, -1, 4, 0,
    -- layer=1 filter=87 channel=93
    -8, 6, -9, -8, -8, -10, 8, -10, 5,
    -- layer=1 filter=87 channel=94
    6, -4, -9, -9, -5, 2, -4, -10, 0,
    -- layer=1 filter=87 channel=95
    -11, 1, -11, 3, -8, 7, -10, 0, 7,
    -- layer=1 filter=87 channel=96
    -4, 0, -6, 0, -6, 3, 1, 3, -6,
    -- layer=1 filter=87 channel=97
    -8, -5, -2, -3, -3, 5, -1, -7, 7,
    -- layer=1 filter=87 channel=98
    -1, -10, -7, 1, 2, -10, -10, -9, 2,
    -- layer=1 filter=87 channel=99
    -6, 0, 1, -10, 8, 7, -6, -3, 0,
    -- layer=1 filter=87 channel=100
    -5, -11, 0, -4, -11, -8, 7, 0, 5,
    -- layer=1 filter=87 channel=101
    0, -5, -11, -4, 6, 6, -10, -10, 3,
    -- layer=1 filter=87 channel=102
    1, 8, -5, -11, -4, -11, -4, -10, -1,
    -- layer=1 filter=87 channel=103
    -7, 0, 4, 5, -9, -7, -10, 0, 6,
    -- layer=1 filter=87 channel=104
    -9, -6, -8, -10, -7, -5, -8, -11, 8,
    -- layer=1 filter=87 channel=105
    -7, 2, -3, 3, -8, 4, -2, -2, -7,
    -- layer=1 filter=87 channel=106
    9, 3, 0, 4, 4, -8, 0, -8, 9,
    -- layer=1 filter=87 channel=107
    0, -9, 8, -4, -10, -2, 10, 7, 2,
    -- layer=1 filter=87 channel=108
    3, 8, 0, -9, -6, -6, -8, 0, -3,
    -- layer=1 filter=87 channel=109
    -10, -10, 6, 8, 4, -1, -5, -1, 9,
    -- layer=1 filter=87 channel=110
    -1, 2, 4, -3, 8, 4, -5, 6, -4,
    -- layer=1 filter=87 channel=111
    -1, 6, 4, 8, -9, -13, 1, -8, -2,
    -- layer=1 filter=87 channel=112
    7, -9, -1, -2, 1, -1, -8, 4, 8,
    -- layer=1 filter=87 channel=113
    1, 3, -10, -4, -1, 4, 10, -7, 9,
    -- layer=1 filter=87 channel=114
    5, -4, -1, 2, 2, -1, -7, -5, -8,
    -- layer=1 filter=87 channel=115
    0, 4, -9, -8, 0, 0, -7, -11, -4,
    -- layer=1 filter=87 channel=116
    10, 0, 0, 2, -9, -6, -2, 5, 5,
    -- layer=1 filter=87 channel=117
    -9, 5, -8, 3, 3, -6, 1, -8, 7,
    -- layer=1 filter=87 channel=118
    -3, -8, 0, 2, -5, -2, -7, -4, -7,
    -- layer=1 filter=87 channel=119
    -4, -2, -3, -3, -1, 0, -9, -6, 4,
    -- layer=1 filter=87 channel=120
    3, -6, -3, -10, 4, -5, 4, 6, 1,
    -- layer=1 filter=87 channel=121
    -8, -8, -10, 5, 2, -4, -13, 3, -8,
    -- layer=1 filter=87 channel=122
    -2, -9, -9, 0, 2, -7, 10, -3, -5,
    -- layer=1 filter=87 channel=123
    0, 0, -6, -6, -4, -4, 5, 7, -10,
    -- layer=1 filter=87 channel=124
    -5, -1, 1, -6, -3, 3, 0, -12, -6,
    -- layer=1 filter=87 channel=125
    -2, -6, 3, -5, 0, 9, -7, -10, 8,
    -- layer=1 filter=87 channel=126
    -3, -2, 8, 8, -11, -11, -11, 1, 3,
    -- layer=1 filter=87 channel=127
    5, -8, -8, -10, 3, -7, -1, 5, -3,
    -- layer=1 filter=88 channel=0
    -4, 4, 3, -3, 0, 0, -12, 4, -3,
    -- layer=1 filter=88 channel=1
    0, -5, 2, -1, -10, -3, -6, -5, -9,
    -- layer=1 filter=88 channel=2
    0, -11, 2, 6, 2, -1, -5, 0, 6,
    -- layer=1 filter=88 channel=3
    2, 0, 0, 8, 8, -9, -7, 4, -5,
    -- layer=1 filter=88 channel=4
    -1, -8, 6, -12, 4, -9, -5, 9, -10,
    -- layer=1 filter=88 channel=5
    -1, -9, -18, 6, -6, -16, -14, -3, 2,
    -- layer=1 filter=88 channel=6
    9, 9, 10, 2, 0, -2, -4, 1, 0,
    -- layer=1 filter=88 channel=7
    5, -11, -11, -9, -11, -10, -4, -10, -10,
    -- layer=1 filter=88 channel=8
    4, -9, -7, -7, -11, -7, 0, 0, -20,
    -- layer=1 filter=88 channel=9
    -11, -15, -2, -2, -16, -12, -7, 2, -13,
    -- layer=1 filter=88 channel=10
    -5, 1, -9, -16, -8, -19, -19, -9, -13,
    -- layer=1 filter=88 channel=11
    0, -5, 1, -3, -1, -12, -2, 0, -13,
    -- layer=1 filter=88 channel=12
    18, 17, 1, -10, -10, -1, -1, 1, -3,
    -- layer=1 filter=88 channel=13
    4, 0, 3, 3, 10, 2, -1, 1, -7,
    -- layer=1 filter=88 channel=14
    -3, 0, -17, -15, -11, -18, -8, -3, -3,
    -- layer=1 filter=88 channel=15
    -11, -11, -6, -5, -7, -4, 2, 2, -14,
    -- layer=1 filter=88 channel=16
    -16, -1, -14, 0, -3, 0, -2, -4, -8,
    -- layer=1 filter=88 channel=17
    1, -8, 3, -3, -10, 7, -10, -1, 6,
    -- layer=1 filter=88 channel=18
    0, -2, 2, -7, -17, 0, -7, -19, -7,
    -- layer=1 filter=88 channel=19
    -16, 1, 0, -2, -12, -10, 4, -12, 2,
    -- layer=1 filter=88 channel=20
    -2, -9, -8, -5, 6, -12, 3, 3, 1,
    -- layer=1 filter=88 channel=21
    0, -2, -1, 6, 2, 0, 7, 5, -3,
    -- layer=1 filter=88 channel=22
    -2, -12, -10, 0, -3, 2, -9, -1, -3,
    -- layer=1 filter=88 channel=23
    -1, -3, -1, -5, -2, -13, -1, 0, -7,
    -- layer=1 filter=88 channel=24
    0, -8, -4, 4, 2, -10, -11, -12, -4,
    -- layer=1 filter=88 channel=25
    -11, -7, -20, 4, -9, -17, 0, 0, -1,
    -- layer=1 filter=88 channel=26
    -11, -15, -7, 3, -13, -4, -8, -20, -2,
    -- layer=1 filter=88 channel=27
    0, 0, -5, 4, 2, -1, -3, 4, 3,
    -- layer=1 filter=88 channel=28
    -12, -1, -16, -2, -4, -5, -14, -16, -21,
    -- layer=1 filter=88 channel=29
    -9, 7, 11, 1, -3, 0, -8, 8, -8,
    -- layer=1 filter=88 channel=30
    -7, -8, -10, -13, -13, -4, -7, -11, 2,
    -- layer=1 filter=88 channel=31
    0, 5, -10, -6, -5, 1, -17, 7, -10,
    -- layer=1 filter=88 channel=32
    3, -27, -20, -1, -11, -7, 7, -7, -5,
    -- layer=1 filter=88 channel=33
    -5, -6, -7, 0, 2, -7, 6, -12, 1,
    -- layer=1 filter=88 channel=34
    -4, -10, 0, -4, 4, -1, 10, 4, -1,
    -- layer=1 filter=88 channel=35
    -3, -7, -8, -1, -1, 0, -8, 7, -12,
    -- layer=1 filter=88 channel=36
    -1, 1, -9, 4, 0, 1, 3, -15, -8,
    -- layer=1 filter=88 channel=37
    -5, -5, -20, -12, 0, -12, -12, -7, -1,
    -- layer=1 filter=88 channel=38
    0, 2, 0, 0, -7, -7, -7, 2, 3,
    -- layer=1 filter=88 channel=39
    -4, -4, 0, -1, -4, -2, 2, -12, -5,
    -- layer=1 filter=88 channel=40
    2, -2, -2, 2, -6, -7, -3, -6, 2,
    -- layer=1 filter=88 channel=41
    1, -15, 5, 8, -5, -2, 9, 5, -10,
    -- layer=1 filter=88 channel=42
    -5, 3, 2, -1, -5, -7, 4, -11, -6,
    -- layer=1 filter=88 channel=43
    0, -11, -12, -1, -6, -16, -12, -20, -9,
    -- layer=1 filter=88 channel=44
    -6, -4, -12, 5, -22, -4, 0, -8, -20,
    -- layer=1 filter=88 channel=45
    3, 3, -2, 7, -12, -2, -4, -12, 1,
    -- layer=1 filter=88 channel=46
    -19, -6, -20, -6, -4, 4, -13, -8, -20,
    -- layer=1 filter=88 channel=47
    -2, -13, -1, 7, -10, -18, 1, -12, -5,
    -- layer=1 filter=88 channel=48
    1, -1, -11, -9, -2, -10, 0, 3, -5,
    -- layer=1 filter=88 channel=49
    6, -11, -3, 1, 2, -3, 9, 0, -4,
    -- layer=1 filter=88 channel=50
    4, 0, 0, 0, 0, -10, -12, -11, -1,
    -- layer=1 filter=88 channel=51
    -14, -7, -8, -11, -12, -5, -6, -8, -2,
    -- layer=1 filter=88 channel=52
    1, -5, -11, -9, -11, -6, 6, 13, 0,
    -- layer=1 filter=88 channel=53
    -12, 4, -4, 8, 3, -7, -7, 3, -7,
    -- layer=1 filter=88 channel=54
    -26, -20, -11, -15, -17, -17, -15, -28, -15,
    -- layer=1 filter=88 channel=55
    -16, -19, -10, -18, -12, -6, -13, -20, -17,
    -- layer=1 filter=88 channel=56
    1, 1, -5, -6, -5, 2, 1, -10, -10,
    -- layer=1 filter=88 channel=57
    -5, 7, -8, -10, 8, -4, -12, 4, -7,
    -- layer=1 filter=88 channel=58
    -2, -15, -24, -15, -5, -23, -10, -16, -15,
    -- layer=1 filter=88 channel=59
    -8, 6, 0, 6, -9, -7, -7, -1, -10,
    -- layer=1 filter=88 channel=60
    -2, -5, 0, 2, -10, 9, -6, 0, -7,
    -- layer=1 filter=88 channel=61
    -2, -11, -10, -3, 3, 0, -3, 0, 7,
    -- layer=1 filter=88 channel=62
    -14, -7, -4, 3, -3, -15, -2, -4, -7,
    -- layer=1 filter=88 channel=63
    -16, -10, 0, -16, -13, -17, -17, -5, -13,
    -- layer=1 filter=88 channel=64
    1, -2, -3, -6, -5, -4, 0, -11, -4,
    -- layer=1 filter=88 channel=65
    0, -10, 1, -12, 0, -4, -2, 0, -11,
    -- layer=1 filter=88 channel=66
    -3, -6, 0, -4, -8, -15, -8, -2, 0,
    -- layer=1 filter=88 channel=67
    -1, -3, 8, 5, -10, 2, -5, 0, 7,
    -- layer=1 filter=88 channel=68
    0, -13, -13, -1, -7, -11, -4, -13, -10,
    -- layer=1 filter=88 channel=69
    0, -20, -7, 0, 0, 4, -15, -11, -1,
    -- layer=1 filter=88 channel=70
    2, 14, -7, -1, -2, 4, 10, 0, -1,
    -- layer=1 filter=88 channel=71
    0, -15, 7, -1, -5, -6, -14, -12, -10,
    -- layer=1 filter=88 channel=72
    -20, -9, -5, 0, -8, -8, -6, -6, -4,
    -- layer=1 filter=88 channel=73
    -8, 4, -13, -15, 0, 3, -12, 1, -9,
    -- layer=1 filter=88 channel=74
    -1, -10, 1, -3, -11, -1, 0, -9, -9,
    -- layer=1 filter=88 channel=75
    9, -1, -9, -8, -7, -15, 2, -12, -3,
    -- layer=1 filter=88 channel=76
    -7, 1, -3, 4, -5, 5, -3, -10, 0,
    -- layer=1 filter=88 channel=77
    -7, -13, 1, -18, -13, -8, -3, -6, -5,
    -- layer=1 filter=88 channel=78
    -10, -2, 4, 1, 4, 8, 6, -8, 3,
    -- layer=1 filter=88 channel=79
    -4, -9, -12, 2, 0, 1, -13, -10, 0,
    -- layer=1 filter=88 channel=80
    -12, -1, -4, 3, -8, 0, 0, 11, 6,
    -- layer=1 filter=88 channel=81
    -3, -16, -8, -22, -17, -23, -6, -19, -23,
    -- layer=1 filter=88 channel=82
    1, -6, -16, -3, -1, -7, -9, 3, -11,
    -- layer=1 filter=88 channel=83
    -4, -11, 0, -10, -9, -4, 1, 3, -12,
    -- layer=1 filter=88 channel=84
    -3, -3, -12, -8, -18, -12, -6, -26, -5,
    -- layer=1 filter=88 channel=85
    -1, -14, -12, -3, -17, -25, -6, -10, -16,
    -- layer=1 filter=88 channel=86
    -5, -19, -1, 2, -11, -1, -6, -3, -7,
    -- layer=1 filter=88 channel=87
    -16, -10, -1, -13, -1, 0, 2, -12, -3,
    -- layer=1 filter=88 channel=88
    4, 11, -1, 6, 6, 0, 6, 6, 7,
    -- layer=1 filter=88 channel=89
    -3, -12, -10, 2, -7, -16, -7, 0, -16,
    -- layer=1 filter=88 channel=90
    -2, -19, -14, -1, -20, 1, -13, -12, 1,
    -- layer=1 filter=88 channel=91
    -6, -6, -11, -7, -5, -1, -2, -3, 3,
    -- layer=1 filter=88 channel=92
    -6, -8, -17, 8, -9, -3, -12, 0, -1,
    -- layer=1 filter=88 channel=93
    -13, -17, -9, -2, 1, 1, -8, 1, -6,
    -- layer=1 filter=88 channel=94
    4, -8, -4, -6, 0, -6, -8, -11, -5,
    -- layer=1 filter=88 channel=95
    -19, -2, -15, -5, -22, -5, 0, -15, -12,
    -- layer=1 filter=88 channel=96
    -5, 0, 0, -13, -7, -4, -3, -8, -10,
    -- layer=1 filter=88 channel=97
    -5, -14, 2, -12, 0, -5, -13, -8, 3,
    -- layer=1 filter=88 channel=98
    -5, 4, -8, 10, -3, -8, -4, 0, -4,
    -- layer=1 filter=88 channel=99
    -7, -13, -5, 2, -12, -12, -7, -10, -2,
    -- layer=1 filter=88 channel=100
    -12, -14, -4, 7, 5, -5, -4, -5, -4,
    -- layer=1 filter=88 channel=101
    -10, -13, -6, 2, -3, -14, -3, 4, -5,
    -- layer=1 filter=88 channel=102
    -11, 6, 2, -5, -4, 2, 2, -1, 6,
    -- layer=1 filter=88 channel=103
    -1, -1, -14, -12, -4, -1, -6, -3, -8,
    -- layer=1 filter=88 channel=104
    8, -8, -10, -5, 5, -1, -5, -9, -13,
    -- layer=1 filter=88 channel=105
    0, -7, 3, 2, -6, 0, 2, 4, -12,
    -- layer=1 filter=88 channel=106
    0, 5, -9, 5, -3, 0, 6, 10, -6,
    -- layer=1 filter=88 channel=107
    -6, 2, 0, 5, -1, 1, 4, -5, -4,
    -- layer=1 filter=88 channel=108
    0, -7, -11, 10, -1, 4, 6, -16, -13,
    -- layer=1 filter=88 channel=109
    0, -1, 7, -4, -4, -10, 6, 6, 6,
    -- layer=1 filter=88 channel=110
    -11, -11, -9, -14, -5, -6, -15, -5, -4,
    -- layer=1 filter=88 channel=111
    -14, -8, -6, -13, -27, -18, -18, -3, -14,
    -- layer=1 filter=88 channel=112
    0, -4, -2, -5, -9, -9, 3, -9, 0,
    -- layer=1 filter=88 channel=113
    -2, 4, -7, -1, 0, 6, -6, -3, -6,
    -- layer=1 filter=88 channel=114
    -13, -12, -6, 8, -9, -7, -15, 1, -9,
    -- layer=1 filter=88 channel=115
    -5, 0, -18, 0, -4, -17, -12, -1, -3,
    -- layer=1 filter=88 channel=116
    -6, -5, -1, -6, -7, 1, 4, -7, -4,
    -- layer=1 filter=88 channel=117
    -16, -6, -23, 0, -7, -14, -6, 3, -8,
    -- layer=1 filter=88 channel=118
    -6, -18, -15, -5, -12, -4, -13, -8, -2,
    -- layer=1 filter=88 channel=119
    -10, -26, -24, 2, -13, 0, -13, -18, -15,
    -- layer=1 filter=88 channel=120
    -15, -9, -9, -8, -3, -5, 0, 9, 0,
    -- layer=1 filter=88 channel=121
    -13, -4, -7, -12, -15, 0, -1, -6, 1,
    -- layer=1 filter=88 channel=122
    5, -3, 3, 10, 0, -7, 1, 4, 8,
    -- layer=1 filter=88 channel=123
    -16, -11, -18, -11, -9, -11, 0, -12, -12,
    -- layer=1 filter=88 channel=124
    -4, 6, -4, -5, -5, -1, -4, 6, 6,
    -- layer=1 filter=88 channel=125
    4, 9, 3, -5, 0, 7, -3, 8, 5,
    -- layer=1 filter=88 channel=126
    -6, -2, 4, -13, -6, -14, 5, -7, -2,
    -- layer=1 filter=88 channel=127
    -8, 0, -17, -2, -12, -20, -6, -17, -11,
    -- layer=1 filter=89 channel=0
    -8, -16, -10, -22, -18, -18, 31, 39, 30,
    -- layer=1 filter=89 channel=1
    -24, 3, -32, 5, -8, 30, 45, 57, 42,
    -- layer=1 filter=89 channel=2
    -2, -9, 6, -7, -14, 6, -10, 3, -11,
    -- layer=1 filter=89 channel=3
    3, -1, -9, 9, -6, 7, 1, 2, -3,
    -- layer=1 filter=89 channel=4
    -22, -11, -21, -11, -10, 0, -1, 3, -7,
    -- layer=1 filter=89 channel=5
    -55, -39, -99, 11, 5, 45, 53, 51, 54,
    -- layer=1 filter=89 channel=6
    7, 0, -11, 51, 51, 38, -29, -43, -87,
    -- layer=1 filter=89 channel=7
    -75, -24, 12, -75, -25, -11, -7, 43, 4,
    -- layer=1 filter=89 channel=8
    -14, -42, -95, -14, -3, 24, 33, 40, 46,
    -- layer=1 filter=89 channel=9
    17, -35, -21, -86, -59, -18, -80, -19, -24,
    -- layer=1 filter=89 channel=10
    -59, -56, 9, -76, 1, -6, 40, 66, 13,
    -- layer=1 filter=89 channel=11
    -6, -39, -45, -73, -114, -83, -16, 6, 8,
    -- layer=1 filter=89 channel=12
    -31, -26, -29, -53, -56, -8, -43, 43, -22,
    -- layer=1 filter=89 channel=13
    27, 7, 1, 17, 6, 3, 0, -23, -20,
    -- layer=1 filter=89 channel=14
    -31, -50, 39, -82, -49, -37, -10, 20, -6,
    -- layer=1 filter=89 channel=15
    -14, 41, 15, -5, -27, 23, -13, -16, 0,
    -- layer=1 filter=89 channel=16
    -15, -31, -81, -6, 21, 25, 47, 52, 34,
    -- layer=1 filter=89 channel=17
    -8, -33, -5, -24, -10, -10, 24, 15, 42,
    -- layer=1 filter=89 channel=18
    12, -14, -14, -90, -89, -52, -2, -24, -50,
    -- layer=1 filter=89 channel=19
    4, -20, -58, -17, 11, 28, 56, 59, 36,
    -- layer=1 filter=89 channel=20
    21, 9, -6, 26, 18, 17, 21, 9, -6,
    -- layer=1 filter=89 channel=21
    -17, 1, 8, 8, 19, 3, 9, 25, -13,
    -- layer=1 filter=89 channel=22
    19, 20, 15, 22, 4, -11, 11, -1, -4,
    -- layer=1 filter=89 channel=23
    -35, -42, -53, -59, -81, -3, 21, 3, 62,
    -- layer=1 filter=89 channel=24
    -13, -28, -47, -9, 8, 11, 3, -2, 16,
    -- layer=1 filter=89 channel=25
    -40, -34, -5, -33, 4, 20, 46, 62, 31,
    -- layer=1 filter=89 channel=26
    45, 0, -8, -2, -27, -4, -6, -26, -29,
    -- layer=1 filter=89 channel=27
    -27, -22, -41, -33, -23, -11, 3, 11, -25,
    -- layer=1 filter=89 channel=28
    -76, -69, -5, -89, 7, -10, 17, 47, 7,
    -- layer=1 filter=89 channel=29
    0, -4, -9, 4, 21, 16, 13, 36, 35,
    -- layer=1 filter=89 channel=30
    19, -24, -4, -28, -49, -2, -46, -84, -98,
    -- layer=1 filter=89 channel=31
    8, -19, -16, 24, 5, 33, 0, -40, -6,
    -- layer=1 filter=89 channel=32
    12, -18, -32, -20, -46, 20, 22, -11, 4,
    -- layer=1 filter=89 channel=33
    15, -9, -2, 30, 19, 14, -10, 20, 16,
    -- layer=1 filter=89 channel=34
    -14, -16, -9, 18, -1, 3, -4, -7, -28,
    -- layer=1 filter=89 channel=35
    -7, -14, -3, -13, -6, 7, 6, 10, 28,
    -- layer=1 filter=89 channel=36
    -10, -45, -48, -88, -102, -72, 2, 10, 48,
    -- layer=1 filter=89 channel=37
    -46, -60, -95, 0, 33, 45, 67, 60, 52,
    -- layer=1 filter=89 channel=38
    4, 9, 11, 16, 25, 18, -3, -17, -49,
    -- layer=1 filter=89 channel=39
    -34, -62, -70, -30, -23, 19, -17, -16, -7,
    -- layer=1 filter=89 channel=40
    19, 20, 31, 42, 43, 26, -23, -54, -78,
    -- layer=1 filter=89 channel=41
    43, -20, -20, -29, -73, -20, 27, -16, 27,
    -- layer=1 filter=89 channel=42
    17, 8, 3, 19, 2, 18, 17, 22, 29,
    -- layer=1 filter=89 channel=43
    -36, -20, -75, -8, 12, -4, 10, 38, 25,
    -- layer=1 filter=89 channel=44
    -14, -40, -30, -12, -59, 0, 5, -8, 5,
    -- layer=1 filter=89 channel=45
    -16, -4, -18, -8, -3, -4, 15, 32, 12,
    -- layer=1 filter=89 channel=46
    -39, -11, -8, 24, 20, 70, 83, 83, 72,
    -- layer=1 filter=89 channel=47
    -9, -15, -6, -8, -10, 50, 78, 51, 87,
    -- layer=1 filter=89 channel=48
    15, 6, 10, -4, 29, -1, -1, -3, -36,
    -- layer=1 filter=89 channel=49
    6, 0, -1, 18, 28, 28, 7, -5, -26,
    -- layer=1 filter=89 channel=50
    27, 28, 17, 0, 12, 0, 10, 12, -1,
    -- layer=1 filter=89 channel=51
    -17, -1, 14, 13, 29, -14, -27, -16, -38,
    -- layer=1 filter=89 channel=52
    16, 29, -13, 10, 16, 1, 3, 7, -4,
    -- layer=1 filter=89 channel=53
    -5, -5, 3, -10, 4, 15, 9, 14, 4,
    -- layer=1 filter=89 channel=54
    -35, -71, -43, -35, 19, 2, 52, 74, 34,
    -- layer=1 filter=89 channel=55
    -73, -71, -57, -64, -75, -41, -22, 0, -7,
    -- layer=1 filter=89 channel=56
    -8, 6, 4, -11, -10, 6, 2, -8, 8,
    -- layer=1 filter=89 channel=57
    -8, -18, 27, -18, 9, -6, 13, 44, 8,
    -- layer=1 filter=89 channel=58
    -56, -21, -30, -34, -31, 17, 55, 55, 44,
    -- layer=1 filter=89 channel=59
    -5, -5, -10, -8, -12, -12, 0, -7, -32,
    -- layer=1 filter=89 channel=60
    -8, -32, 2, 20, 14, -31, 0, 17, -25,
    -- layer=1 filter=89 channel=61
    -9, -3, 11, -2, 6, 8, 4, 10, 8,
    -- layer=1 filter=89 channel=62
    -6, -32, -97, -1, 15, 41, 35, 48, 40,
    -- layer=1 filter=89 channel=63
    3, -27, -30, -64, -93, -57, -22, 39, 24,
    -- layer=1 filter=89 channel=64
    -15, -1, -4, 20, -3, -3, 8, 19, -3,
    -- layer=1 filter=89 channel=65
    16, 12, 10, 9, 6, -13, -15, -1, -46,
    -- layer=1 filter=89 channel=66
    -42, -42, -32, -57, -49, -15, 15, 42, 36,
    -- layer=1 filter=89 channel=67
    -68, -45, -42, -36, -12, -4, -76, -45, -64,
    -- layer=1 filter=89 channel=68
    -27, -51, -27, -27, -89, -29, -10, -16, -7,
    -- layer=1 filter=89 channel=69
    -38, -16, -84, -5, -21, 14, 22, 30, 29,
    -- layer=1 filter=89 channel=70
    -58, -34, -26, 23, 51, 28, -32, -10, 9,
    -- layer=1 filter=89 channel=71
    -37, -24, -34, -11, 11, -9, 8, 15, -1,
    -- layer=1 filter=89 channel=72
    37, -1, -25, -27, -60, 3, 27, -23, -2,
    -- layer=1 filter=89 channel=73
    -7, -12, 2, -20, -9, -2, -3, -8, 5,
    -- layer=1 filter=89 channel=74
    3, -50, -15, 19, -13, 5, 6, -60, -57,
    -- layer=1 filter=89 channel=75
    -3, -16, 9, -69, -86, -1, -82, -114, -58,
    -- layer=1 filter=89 channel=76
    28, -23, -32, -51, -50, -32, -18, -35, -19,
    -- layer=1 filter=89 channel=77
    -15, -10, -4, -18, 12, -21, -19, 23, 10,
    -- layer=1 filter=89 channel=78
    -35, -56, -19, -48, -32, -26, 41, 31, 17,
    -- layer=1 filter=89 channel=79
    -2, -7, -61, -2, 20, 32, 49, 49, 49,
    -- layer=1 filter=89 channel=80
    -22, 6, 5, -5, -23, -29, 39, -6, 8,
    -- layer=1 filter=89 channel=81
    -45, -35, -40, -39, 3, 4, -5, 16, 24,
    -- layer=1 filter=89 channel=82
    6, 6, -3, 22, 30, 2, -18, -4, -31,
    -- layer=1 filter=89 channel=83
    -29, -43, -17, -27, -30, 6, -5, 4, 31,
    -- layer=1 filter=89 channel=84
    14, -24, -5, -7, -29, -12, -21, -70, -99,
    -- layer=1 filter=89 channel=85
    -16, -29, -16, -29, -5, 19, 51, 40, 63,
    -- layer=1 filter=89 channel=86
    -53, -71, -58, -59, -82, 0, 14, 29, 31,
    -- layer=1 filter=89 channel=87
    6, -39, -38, -37, -42, 3, 48, 59, 88,
    -- layer=1 filter=89 channel=88
    -2, 4, 9, -8, 2, -12, -8, -9, -17,
    -- layer=1 filter=89 channel=89
    -2, 5, 1, 10, 0, 18, -33, -30, -50,
    -- layer=1 filter=89 channel=90
    -16, -68, -34, -13, -63, 0, 13, -11, 21,
    -- layer=1 filter=89 channel=91
    10, 7, 25, 16, 32, 14, -20, -6, -34,
    -- layer=1 filter=89 channel=92
    -11, -3, 28, -43, -66, 27, -10, -7, 36,
    -- layer=1 filter=89 channel=93
    -22, 3, -5, -8, -2, -19, 9, 5, 5,
    -- layer=1 filter=89 channel=94
    -22, -25, 7, -39, -50, -18, 14, 37, 21,
    -- layer=1 filter=89 channel=95
    29, -14, -13, -37, -63, -21, -39, -108, -107,
    -- layer=1 filter=89 channel=96
    -13, -46, -38, -28, -18, -29, 20, -1, 4,
    -- layer=1 filter=89 channel=97
    -7, -9, 0, -19, -12, -7, 8, 18, 30,
    -- layer=1 filter=89 channel=98
    2, -3, -47, -18, 1, -10, 42, 42, 33,
    -- layer=1 filter=89 channel=99
    -94, -103, -7, -91, -27, -56, -11, 47, 2,
    -- layer=1 filter=89 channel=100
    19, -37, -15, -75, -91, -54, 1, 38, 9,
    -- layer=1 filter=89 channel=101
    10, 5, 1, 20, 25, 13, -9, -24, -34,
    -- layer=1 filter=89 channel=102
    -4, -21, -1, 19, 15, 11, 1, 29, 11,
    -- layer=1 filter=89 channel=103
    3, -32, -18, -68, -92, -43, 19, 9, 16,
    -- layer=1 filter=89 channel=104
    17, 0, 3, -29, -24, -1, 26, 21, 46,
    -- layer=1 filter=89 channel=105
    -27, -19, -5, -43, -27, -30, 2, 20, 24,
    -- layer=1 filter=89 channel=106
    12, 1, -7, 19, 0, 2, -19, -43, -44,
    -- layer=1 filter=89 channel=107
    2, 10, 13, 17, 20, 12, 18, 23, 10,
    -- layer=1 filter=89 channel=108
    -2, -34, -51, -29, -58, 4, 25, 16, 20,
    -- layer=1 filter=89 channel=109
    -6, -1, -8, 2, -3, -9, 8, 6, -2,
    -- layer=1 filter=89 channel=110
    -19, -12, 7, -16, -22, -29, 4, -2, -37,
    -- layer=1 filter=89 channel=111
    24, -16, 9, -35, -32, -33, -60, -74, -87,
    -- layer=1 filter=89 channel=112
    6, -10, 0, -38, -42, -32, 8, 8, -16,
    -- layer=1 filter=89 channel=113
    15, 20, 11, 45, 25, 18, 35, 29, 6,
    -- layer=1 filter=89 channel=114
    -45, -61, -89, -5, -1, 38, 11, 16, -7,
    -- layer=1 filter=89 channel=115
    -75, -34, -18, -63, -33, -28, 5, 18, 13,
    -- layer=1 filter=89 channel=116
    -8, -6, 1, 0, -5, -8, 0, -7, -4,
    -- layer=1 filter=89 channel=117
    -12, -37, 5, -60, -52, -71, -16, 6, -9,
    -- layer=1 filter=89 channel=118
    10, -38, -22, 2, -12, 17, -53, -103, -103,
    -- layer=1 filter=89 channel=119
    2, -40, -53, -25, -57, -6, 0, -27, 9,
    -- layer=1 filter=89 channel=120
    -1, 13, 5, -21, 23, 0, 5, 25, 11,
    -- layer=1 filter=89 channel=121
    -1, -57, -47, -86, -52, 0, 40, 37, 19,
    -- layer=1 filter=89 channel=122
    -6, 5, 0, 7, -10, 6, 9, 7, -3,
    -- layer=1 filter=89 channel=123
    -2, -24, -26, -62, -79, -5, -3, 14, 9,
    -- layer=1 filter=89 channel=124
    -13, 5, 8, -10, 12, -8, 3, 9, 2,
    -- layer=1 filter=89 channel=125
    -36, -38, -28, 18, 45, 19, -3, 4, -6,
    -- layer=1 filter=89 channel=126
    -42, -60, -44, -42, 18, 22, 58, 62, 79,
    -- layer=1 filter=89 channel=127
    1, -33, -17, -29, -29, 14, -42, -126, -93,
    -- layer=1 filter=90 channel=0
    -7, 0, -9, -10, -1, -8, 8, 5, -6,
    -- layer=1 filter=90 channel=1
    -1, 4, -9, 7, 1, 1, -7, -2, 1,
    -- layer=1 filter=90 channel=2
    7, 0, -5, -4, -4, -4, 9, 1, 2,
    -- layer=1 filter=90 channel=3
    9, 1, 9, 0, 0, 5, -4, 6, 2,
    -- layer=1 filter=90 channel=4
    -7, -8, 6, 3, -1, 4, 0, 0, -1,
    -- layer=1 filter=90 channel=5
    4, 0, -6, -2, -7, 0, -5, -8, -10,
    -- layer=1 filter=90 channel=6
    10, -10, -8, -6, -3, 10, -10, 6, 4,
    -- layer=1 filter=90 channel=7
    -6, 7, 9, -8, -6, 10, 1, -6, 9,
    -- layer=1 filter=90 channel=8
    -11, 1, -3, -8, 4, 6, -3, -7, 6,
    -- layer=1 filter=90 channel=9
    -1, -2, 0, 1, 6, -7, -4, -10, 6,
    -- layer=1 filter=90 channel=10
    -3, 3, -3, -9, 6, 9, -9, -6, -7,
    -- layer=1 filter=90 channel=11
    -4, -6, -12, 1, -6, 2, 2, 8, 0,
    -- layer=1 filter=90 channel=12
    -3, 0, -10, -10, 5, -1, 7, 8, 10,
    -- layer=1 filter=90 channel=13
    -10, 6, 4, 5, 9, 2, -12, -11, -6,
    -- layer=1 filter=90 channel=14
    -8, 5, -5, 8, 2, 3, 1, 6, -3,
    -- layer=1 filter=90 channel=15
    6, 2, 10, 5, 2, -6, 8, 7, -1,
    -- layer=1 filter=90 channel=16
    3, -13, -4, -6, -5, 0, -5, 4, -7,
    -- layer=1 filter=90 channel=17
    -7, -8, -5, 0, 0, -8, 3, -10, -9,
    -- layer=1 filter=90 channel=18
    -6, -8, -7, 0, 3, -2, -5, -3, 2,
    -- layer=1 filter=90 channel=19
    -6, -8, 3, -7, 2, -11, -5, 7, 5,
    -- layer=1 filter=90 channel=20
    -11, 1, 0, 0, -1, -1, -1, 1, -5,
    -- layer=1 filter=90 channel=21
    2, -2, 3, 0, -5, -3, 2, 6, -4,
    -- layer=1 filter=90 channel=22
    3, 3, -3, 6, 5, 7, -4, -1, -1,
    -- layer=1 filter=90 channel=23
    -4, -2, 6, 5, 6, -5, -8, 9, -8,
    -- layer=1 filter=90 channel=24
    -12, -10, 0, 1, 3, -12, -11, -11, -9,
    -- layer=1 filter=90 channel=25
    -6, 4, 5, -1, 1, 3, 3, 9, -1,
    -- layer=1 filter=90 channel=26
    7, -1, 9, -5, -4, 4, -10, 0, -6,
    -- layer=1 filter=90 channel=27
    -5, -2, 8, -6, -4, 6, 5, 0, -6,
    -- layer=1 filter=90 channel=28
    -6, -14, -8, 0, 0, -6, 7, 1, 6,
    -- layer=1 filter=90 channel=29
    -7, -4, -1, -7, 1, 4, 1, 1, -9,
    -- layer=1 filter=90 channel=30
    8, 1, 8, 4, 4, 4, -8, 10, 4,
    -- layer=1 filter=90 channel=31
    10, -4, 6, -12, 0, -6, -6, -7, 0,
    -- layer=1 filter=90 channel=32
    -8, -7, 0, 1, 0, 0, -9, -8, -6,
    -- layer=1 filter=90 channel=33
    -9, 3, 9, 8, -1, -5, -5, -1, -3,
    -- layer=1 filter=90 channel=34
    0, 1, -8, -4, 6, 8, -10, 9, -7,
    -- layer=1 filter=90 channel=35
    3, -7, -4, -10, 4, 1, -2, -4, 10,
    -- layer=1 filter=90 channel=36
    4, 0, 2, 0, 2, 0, -2, -2, -4,
    -- layer=1 filter=90 channel=37
    -5, -1, -5, 0, 5, 7, 7, -9, -10,
    -- layer=1 filter=90 channel=38
    3, 3, 5, -13, 4, -12, -11, 7, -11,
    -- layer=1 filter=90 channel=39
    4, 0, -1, -1, 6, -5, 2, -9, -7,
    -- layer=1 filter=90 channel=40
    -4, 4, -7, -3, -9, 0, 4, -9, 2,
    -- layer=1 filter=90 channel=41
    1, 5, -3, 0, 10, -5, 5, 6, 0,
    -- layer=1 filter=90 channel=42
    8, 7, -6, 4, 1, 3, 3, -3, 4,
    -- layer=1 filter=90 channel=43
    6, 0, 0, -7, 10, -8, -8, -10, -4,
    -- layer=1 filter=90 channel=44
    0, 3, -11, -4, 9, -4, -6, 8, 4,
    -- layer=1 filter=90 channel=45
    0, 1, 4, 0, 1, 1, -5, -8, -5,
    -- layer=1 filter=90 channel=46
    -6, -5, 2, -3, 2, 7, 3, 8, -4,
    -- layer=1 filter=90 channel=47
    -7, -5, -9, -3, -10, -10, -1, 4, 6,
    -- layer=1 filter=90 channel=48
    4, 0, 3, 2, -3, -3, -11, -11, 3,
    -- layer=1 filter=90 channel=49
    0, -7, -7, -8, 5, 6, -4, 2, -2,
    -- layer=1 filter=90 channel=50
    9, 1, 0, -8, -9, 2, -6, -2, 2,
    -- layer=1 filter=90 channel=51
    -3, -3, -3, -8, -8, -2, 6, 2, 3,
    -- layer=1 filter=90 channel=52
    -9, 2, 2, 9, 8, -4, -5, 8, -6,
    -- layer=1 filter=90 channel=53
    6, -9, -3, 0, -7, 1, 7, -9, 1,
    -- layer=1 filter=90 channel=54
    -1, 0, 0, -5, 8, -5, 3, 6, 6,
    -- layer=1 filter=90 channel=55
    0, -8, 1, -5, 8, 4, 5, -7, -1,
    -- layer=1 filter=90 channel=56
    -10, 2, -4, 7, 9, 5, -6, -4, -10,
    -- layer=1 filter=90 channel=57
    0, -9, -1, -7, -3, 0, -4, 8, -10,
    -- layer=1 filter=90 channel=58
    -8, -5, 8, -8, -6, -9, 3, 1, -4,
    -- layer=1 filter=90 channel=59
    -3, -10, 6, -7, 1, 2, -9, -3, 0,
    -- layer=1 filter=90 channel=60
    0, 0, -4, -5, 0, -3, 1, 4, -1,
    -- layer=1 filter=90 channel=61
    8, 0, 3, -2, 7, -8, 8, -2, 8,
    -- layer=1 filter=90 channel=62
    4, 0, 0, 0, -1, 9, -1, -1, 8,
    -- layer=1 filter=90 channel=63
    -9, -9, -10, -10, 1, -8, -3, -6, 9,
    -- layer=1 filter=90 channel=64
    -6, -9, 5, -10, 0, -4, 8, -1, 9,
    -- layer=1 filter=90 channel=65
    -8, 5, 4, -10, -13, -10, 9, -6, -7,
    -- layer=1 filter=90 channel=66
    3, -12, -3, -7, 2, -8, -2, -6, -10,
    -- layer=1 filter=90 channel=67
    -7, 0, 2, 2, 6, -2, -6, 2, -8,
    -- layer=1 filter=90 channel=68
    -4, 4, 4, -3, -7, -11, 6, 0, -9,
    -- layer=1 filter=90 channel=69
    -5, 2, -7, -2, -6, 4, -4, -4, 3,
    -- layer=1 filter=90 channel=70
    2, -9, -11, -7, -6, 1, -10, 2, 9,
    -- layer=1 filter=90 channel=71
    6, -1, -4, 5, -10, -9, -3, -6, -7,
    -- layer=1 filter=90 channel=72
    -8, -5, -2, 2, 4, -6, 4, 7, -10,
    -- layer=1 filter=90 channel=73
    -6, -6, -3, -9, 2, 3, 1, 0, -10,
    -- layer=1 filter=90 channel=74
    7, 0, 2, -4, 2, 6, 2, -4, -10,
    -- layer=1 filter=90 channel=75
    -4, 0, -4, -6, -2, 4, 1, -8, -9,
    -- layer=1 filter=90 channel=76
    0, -1, -6, -7, -11, 4, -3, -2, 0,
    -- layer=1 filter=90 channel=77
    1, 6, -11, -3, -7, 1, -8, -7, 0,
    -- layer=1 filter=90 channel=78
    5, 2, 8, 0, 6, 4, -1, 8, -7,
    -- layer=1 filter=90 channel=79
    -9, 7, -4, -6, 2, 1, 9, 0, 7,
    -- layer=1 filter=90 channel=80
    7, -7, -5, 7, -6, -8, 9, -2, -9,
    -- layer=1 filter=90 channel=81
    -5, 1, 8, -1, -3, 7, -3, 3, -8,
    -- layer=1 filter=90 channel=82
    0, -8, -11, 7, -1, -5, 4, 0, -10,
    -- layer=1 filter=90 channel=83
    -6, -8, -4, 2, -8, -2, 0, -7, -4,
    -- layer=1 filter=90 channel=84
    -10, -9, -6, -7, -6, 0, -12, 1, 2,
    -- layer=1 filter=90 channel=85
    -2, 4, -8, -9, 6, -10, 2, -1, -2,
    -- layer=1 filter=90 channel=86
    -4, 1, -10, 0, 4, -2, 5, 0, -9,
    -- layer=1 filter=90 channel=87
    -9, 6, 8, 8, 0, 6, 3, -1, -5,
    -- layer=1 filter=90 channel=88
    -1, -2, 1, -3, -1, 2, -9, -11, -2,
    -- layer=1 filter=90 channel=89
    1, -12, 4, -5, -12, 4, 0, 3, 6,
    -- layer=1 filter=90 channel=90
    0, -1, -5, -7, 1, 3, 4, -2, 9,
    -- layer=1 filter=90 channel=91
    -8, 8, 2, -2, 1, -10, -11, -8, 4,
    -- layer=1 filter=90 channel=92
    6, -3, -10, 2, 8, -2, 0, -1, -8,
    -- layer=1 filter=90 channel=93
    -12, 4, -7, -8, 7, 4, -11, -3, 0,
    -- layer=1 filter=90 channel=94
    4, -12, -14, 1, 0, 6, -10, -3, -10,
    -- layer=1 filter=90 channel=95
    3, 5, -5, -3, -10, -3, -5, -4, 10,
    -- layer=1 filter=90 channel=96
    -6, 2, 2, -7, 0, -7, -9, 9, 6,
    -- layer=1 filter=90 channel=97
    -9, 2, -11, 5, -6, 0, -2, -7, -3,
    -- layer=1 filter=90 channel=98
    -9, 8, -3, -4, -3, -7, -2, -4, 1,
    -- layer=1 filter=90 channel=99
    -10, 6, 8, 4, 9, -3, -5, -9, -10,
    -- layer=1 filter=90 channel=100
    0, -2, -9, -10, -7, 5, 1, -1, 10,
    -- layer=1 filter=90 channel=101
    5, -8, -5, -6, -10, -4, -8, -5, -10,
    -- layer=1 filter=90 channel=102
    5, -11, 7, 1, 1, -4, 2, -2, 5,
    -- layer=1 filter=90 channel=103
    -3, -1, -2, 2, 5, -5, -11, -4, -1,
    -- layer=1 filter=90 channel=104
    1, -1, -6, 5, 0, 6, 9, 8, 5,
    -- layer=1 filter=90 channel=105
    -8, 3, 5, -5, -5, -5, 2, -4, -8,
    -- layer=1 filter=90 channel=106
    6, 2, -7, 3, 1, -4, 1, -2, -6,
    -- layer=1 filter=90 channel=107
    -4, -2, 7, -5, 6, -5, -10, -8, 10,
    -- layer=1 filter=90 channel=108
    -2, 5, 0, -8, -3, -7, 6, -6, -5,
    -- layer=1 filter=90 channel=109
    -8, 0, 9, -7, -8, 0, -2, 10, 7,
    -- layer=1 filter=90 channel=110
    5, -7, -11, 5, -2, -8, 4, 1, 8,
    -- layer=1 filter=90 channel=111
    -8, 6, 4, 5, -6, -12, -13, 10, 3,
    -- layer=1 filter=90 channel=112
    -10, 7, 6, -2, -3, 2, -8, 8, 8,
    -- layer=1 filter=90 channel=113
    -5, 6, 6, -5, 0, -10, 7, -10, 2,
    -- layer=1 filter=90 channel=114
    -6, 5, -8, -8, -5, 8, -8, 6, 0,
    -- layer=1 filter=90 channel=115
    -5, -10, -10, -7, -4, -9, 0, -5, 3,
    -- layer=1 filter=90 channel=116
    -2, 0, -8, -2, 0, 3, 5, 10, 7,
    -- layer=1 filter=90 channel=117
    5, 2, -5, 5, -8, 6, 1, 9, -5,
    -- layer=1 filter=90 channel=118
    -5, -5, -8, -8, -3, -14, 5, 3, 3,
    -- layer=1 filter=90 channel=119
    2, 5, 7, -9, -11, -2, 5, 0, -3,
    -- layer=1 filter=90 channel=120
    1, -10, 0, 1, -1, 0, -5, -8, -10,
    -- layer=1 filter=90 channel=121
    -1, 2, 0, 3, 6, -9, -2, -10, -10,
    -- layer=1 filter=90 channel=122
    -5, 9, 1, -5, 0, 1, 10, 0, 6,
    -- layer=1 filter=90 channel=123
    -1, -5, -7, 0, 4, -2, 0, -6, -9,
    -- layer=1 filter=90 channel=124
    10, 1, -1, 5, 0, -7, 3, 0, 2,
    -- layer=1 filter=90 channel=125
    5, 2, -8, 9, -8, 1, 0, 7, -1,
    -- layer=1 filter=90 channel=126
    0, -2, -1, -1, 10, -6, 0, -9, 9,
    -- layer=1 filter=90 channel=127
    -6, -3, -7, -11, -5, -12, 0, -6, -6,
    -- layer=1 filter=91 channel=0
    -43, -51, -23, -25, -34, -22, -9, -30, -16,
    -- layer=1 filter=91 channel=1
    -3, -13, -32, -6, 0, 31, -5, 13, 13,
    -- layer=1 filter=91 channel=2
    30, 56, 29, 42, 35, 36, 59, 53, 9,
    -- layer=1 filter=91 channel=3
    2, 0, 0, 6, -9, -12, 0, 0, -4,
    -- layer=1 filter=91 channel=4
    -15, -17, -15, 13, -14, -10, -21, -9, -13,
    -- layer=1 filter=91 channel=5
    19, -26, -41, 8, 13, 44, -11, 22, 3,
    -- layer=1 filter=91 channel=6
    9, 18, 7, -9, 16, 2, 0, 16, 19,
    -- layer=1 filter=91 channel=7
    7, 14, 9, -18, 41, 40, -6, 87, 19,
    -- layer=1 filter=91 channel=8
    13, -41, -59, -3, 23, 47, 6, 24, 0,
    -- layer=1 filter=91 channel=9
    -5, -1, -26, 13, -25, 0, -28, -4, -13,
    -- layer=1 filter=91 channel=10
    -13, 0, 42, 3, 66, 46, -15, 74, 33,
    -- layer=1 filter=91 channel=11
    15, -16, -46, 15, -4, -48, -21, -22, -26,
    -- layer=1 filter=91 channel=12
    -22, -33, 5, 11, -25, -41, -37, 41, -74,
    -- layer=1 filter=91 channel=13
    7, 17, 1, 5, 2, 4, 12, 0, 16,
    -- layer=1 filter=91 channel=14
    -23, 22, 26, -30, 0, -17, -20, 48, -25,
    -- layer=1 filter=91 channel=15
    28, 4, -28, 14, 1, 20, 0, 8, -24,
    -- layer=1 filter=91 channel=16
    15, -32, -6, 2, 35, 57, 13, 30, 7,
    -- layer=1 filter=91 channel=17
    -60, -90, -51, -47, -48, -54, -27, -33, -13,
    -- layer=1 filter=91 channel=18
    -23, 20, 6, -43, -14, -55, -64, -16, -22,
    -- layer=1 filter=91 channel=19
    -31, -36, 5, 0, 25, 36, 26, 4, -8,
    -- layer=1 filter=91 channel=20
    14, 6, -2, 7, 15, 24, -4, -1, 26,
    -- layer=1 filter=91 channel=21
    -7, -8, -16, -14, -1, 26, 11, 19, 35,
    -- layer=1 filter=91 channel=22
    12, -3, -4, 0, 0, 21, 8, 9, 18,
    -- layer=1 filter=91 channel=23
    -35, -30, -85, -40, 20, -61, 11, 48, -14,
    -- layer=1 filter=91 channel=24
    -21, -50, -24, 8, 5, -6, 21, 0, -14,
    -- layer=1 filter=91 channel=25
    9, -9, 16, 11, 54, 58, -5, 82, 7,
    -- layer=1 filter=91 channel=26
    -1, 3, -9, 10, 10, -19, 41, 3, 3,
    -- layer=1 filter=91 channel=27
    -35, -51, -36, -30, -56, -24, -12, -10, 9,
    -- layer=1 filter=91 channel=28
    -18, -13, -7, -25, -5, 30, -36, 75, 28,
    -- layer=1 filter=91 channel=29
    -11, 14, 41, 11, 16, 43, 16, 5, 29,
    -- layer=1 filter=91 channel=30
    -58, -28, -5, -31, -26, -47, -82, -17, -28,
    -- layer=1 filter=91 channel=31
    -15, 7, -21, -17, -40, -41, -21, 1, -20,
    -- layer=1 filter=91 channel=32
    4, 16, -34, 35, 30, -1, 32, 37, 10,
    -- layer=1 filter=91 channel=33
    -15, -17, -8, -14, 6, 18, 7, 8, 26,
    -- layer=1 filter=91 channel=34
    -9, -33, -9, -35, -42, -13, -24, -25, 1,
    -- layer=1 filter=91 channel=35
    5, 8, 14, 4, 4, 11, 24, -3, 15,
    -- layer=1 filter=91 channel=36
    -9, -41, -49, -14, -99, -77, -11, -42, -26,
    -- layer=1 filter=91 channel=37
    17, -35, 4, 12, 39, 42, -3, 38, -3,
    -- layer=1 filter=91 channel=38
    -6, 14, 8, 3, 14, 21, 5, 0, 15,
    -- layer=1 filter=91 channel=39
    -40, -62, -37, -28, -37, -35, -1, -14, -19,
    -- layer=1 filter=91 channel=40
    5, 25, 40, -16, 10, -4, -21, 18, 28,
    -- layer=1 filter=91 channel=41
    -9, 14, -21, 7, 28, 14, 22, 60, 53,
    -- layer=1 filter=91 channel=42
    52, 66, 55, 47, 63, 41, 50, 60, 16,
    -- layer=1 filter=91 channel=43
    1, -23, -36, -1, 23, 57, -11, 29, 0,
    -- layer=1 filter=91 channel=44
    9, -2, -31, 17, 30, -9, 35, 11, -9,
    -- layer=1 filter=91 channel=45
    -4, -16, -7, 12, 1, 17, 10, 10, -2,
    -- layer=1 filter=91 channel=46
    28, 6, 18, 45, 26, 24, 11, 6, -7,
    -- layer=1 filter=91 channel=47
    -19, 13, -50, 8, 58, -2, 20, 34, 11,
    -- layer=1 filter=91 channel=48
    -27, -30, -26, -18, -6, 6, 0, 24, 18,
    -- layer=1 filter=91 channel=49
    4, 27, 5, 15, 16, -1, 12, 28, 6,
    -- layer=1 filter=91 channel=50
    -23, -15, -22, -15, -29, -21, -9, -13, -4,
    -- layer=1 filter=91 channel=51
    0, 1, 9, -13, 21, 17, -25, 43, 36,
    -- layer=1 filter=91 channel=52
    -2, -16, 3, 10, 11, 4, 1, 5, 5,
    -- layer=1 filter=91 channel=53
    9, -16, 14, -13, 4, 22, 11, 20, 4,
    -- layer=1 filter=91 channel=54
    21, -19, 19, 18, 81, 73, 13, 84, -3,
    -- layer=1 filter=91 channel=55
    11, -16, -30, -21, -24, -13, -5, 0, -17,
    -- layer=1 filter=91 channel=56
    6, 10, 6, -2, -1, 8, 0, 10, -9,
    -- layer=1 filter=91 channel=57
    -2, 7, 27, -24, 47, 43, -15, 68, 21,
    -- layer=1 filter=91 channel=58
    -17, 8, 4, -22, 71, 14, 26, 86, 1,
    -- layer=1 filter=91 channel=59
    -10, -3, 5, 10, -2, -10, -23, 26, -1,
    -- layer=1 filter=91 channel=60
    -24, 4, 19, -8, 25, 10, -28, 3, -10,
    -- layer=1 filter=91 channel=61
    -11, -9, 4, -13, -10, -19, -3, -4, -10,
    -- layer=1 filter=91 channel=62
    0, -26, -3, -12, 35, 47, 12, 29, -2,
    -- layer=1 filter=91 channel=63
    -34, -44, -45, -24, -55, -48, -11, -24, -5,
    -- layer=1 filter=91 channel=64
    -11, -19, -4, -15, -14, 7, -3, -3, 21,
    -- layer=1 filter=91 channel=65
    -42, -25, -22, -25, -2, 13, 2, 13, 30,
    -- layer=1 filter=91 channel=66
    -24, -55, -52, -30, -62, -20, -14, 0, 4,
    -- layer=1 filter=91 channel=67
    -24, -28, -39, -11, -17, -23, -15, -3, 14,
    -- layer=1 filter=91 channel=68
    9, -6, -26, 29, 2, 21, 46, 29, 10,
    -- layer=1 filter=91 channel=69
    29, -9, -15, 13, 27, 15, 28, -9, -21,
    -- layer=1 filter=91 channel=70
    8, 8, 5, -21, 5, -13, -10, 18, 24,
    -- layer=1 filter=91 channel=71
    -74, -75, -48, -43, -36, 11, -12, 30, 16,
    -- layer=1 filter=91 channel=72
    -16, -23, -32, -21, 4, 19, -26, -36, -6,
    -- layer=1 filter=91 channel=73
    -4, -21, -9, 0, -24, -3, 0, -2, 0,
    -- layer=1 filter=91 channel=74
    -9, 17, -40, -37, -19, -19, 23, 6, 21,
    -- layer=1 filter=91 channel=75
    -15, 1, -16, -32, -36, -52, -46, 11, -71,
    -- layer=1 filter=91 channel=76
    -33, -63, -56, -4, -6, -40, -6, 8, -9,
    -- layer=1 filter=91 channel=77
    -48, -60, -37, -18, -27, 19, -2, 10, 39,
    -- layer=1 filter=91 channel=78
    -64, -31, 3, -41, 3, 18, -21, 17, 5,
    -- layer=1 filter=91 channel=79
    7, -26, -20, -12, 37, 47, 6, 36, -3,
    -- layer=1 filter=91 channel=80
    9, 9, -28, -1, 6, 5, 6, 27, -7,
    -- layer=1 filter=91 channel=81
    -76, -119, -93, -34, -37, 10, -14, 15, 0,
    -- layer=1 filter=91 channel=82
    -14, -11, -22, -4, 7, 6, 12, 21, 24,
    -- layer=1 filter=91 channel=83
    -34, -29, -80, -14, -15, 6, 1, -11, -26,
    -- layer=1 filter=91 channel=84
    -27, -1, -37, 5, -10, -33, -21, 8, -34,
    -- layer=1 filter=91 channel=85
    -35, -14, -36, -42, 38, -19, 38, 65, -12,
    -- layer=1 filter=91 channel=86
    -10, -43, -49, -39, -78, -42, -23, -15, -4,
    -- layer=1 filter=91 channel=87
    4, 11, 0, -33, 6, -1, 7, -6, -30,
    -- layer=1 filter=91 channel=88
    -3, -2, -12, 2, 16, 0, 10, 7, 23,
    -- layer=1 filter=91 channel=89
    -23, -19, -33, 0, -14, -1, 21, -2, 15,
    -- layer=1 filter=91 channel=90
    2, -26, -34, 1, 8, -16, 25, -2, -12,
    -- layer=1 filter=91 channel=91
    7, 15, 16, -4, -3, 4, -8, 0, 11,
    -- layer=1 filter=91 channel=92
    13, 27, 2, 31, 45, 6, 51, -7, 8,
    -- layer=1 filter=91 channel=93
    -42, -34, -46, -22, -20, -6, -8, 14, 11,
    -- layer=1 filter=91 channel=94
    -60, -66, -19, -41, -56, -13, -20, -19, -13,
    -- layer=1 filter=91 channel=95
    -40, -11, -25, -31, -34, -66, -36, -40, -47,
    -- layer=1 filter=91 channel=96
    -16, -44, -47, -8, -12, -22, 23, 1, -35,
    -- layer=1 filter=91 channel=97
    -54, -74, -51, -49, -57, -13, -18, -11, -3,
    -- layer=1 filter=91 channel=98
    -4, -39, -31, -20, 36, 67, -4, 33, -7,
    -- layer=1 filter=91 channel=99
    -30, -5, -8, -19, 5, 2, -42, 29, 23,
    -- layer=1 filter=91 channel=100
    -12, -18, -97, -43, -10, -65, -6, -12, -11,
    -- layer=1 filter=91 channel=101
    -2, 12, -8, -2, -1, -1, 4, 9, 25,
    -- layer=1 filter=91 channel=102
    -55, -70, -17, -55, -52, -32, -48, -36, -25,
    -- layer=1 filter=91 channel=103
    0, -46, -17, 16, -51, -44, 20, -9, 17,
    -- layer=1 filter=91 channel=104
    -19, 17, -26, -10, 4, -46, -23, 70, -18,
    -- layer=1 filter=91 channel=105
    -52, -62, -22, -33, -42, -13, -21, -9, 0,
    -- layer=1 filter=91 channel=106
    2, 10, -10, 25, 0, 4, 19, 0, 4,
    -- layer=1 filter=91 channel=107
    5, 20, 3, 11, 3, 12, 29, 22, 19,
    -- layer=1 filter=91 channel=108
    1, -3, -42, 8, 35, -12, 43, 20, -3,
    -- layer=1 filter=91 channel=109
    -2, -9, 5, -1, 3, 1, 7, -1, -3,
    -- layer=1 filter=91 channel=110
    -24, -15, -17, -27, -25, -2, -6, 0, 18,
    -- layer=1 filter=91 channel=111
    -40, -5, -12, -63, -33, -59, -65, -32, -9,
    -- layer=1 filter=91 channel=112
    -20, -36, -7, -31, -23, -41, -41, -7, -35,
    -- layer=1 filter=91 channel=113
    18, 29, 29, 4, 25, 38, 7, 49, 29,
    -- layer=1 filter=91 channel=114
    48, -3, 0, -8, -2, 20, -10, -10, 0,
    -- layer=1 filter=91 channel=115
    -61, -37, -5, -39, -17, 8, -53, 36, 10,
    -- layer=1 filter=91 channel=116
    -4, -4, -10, 9, 3, 8, -7, 2, 4,
    -- layer=1 filter=91 channel=117
    -46, -29, 27, -31, -31, -41, -54, -39, -8,
    -- layer=1 filter=91 channel=118
    -26, 0, -31, -2, -33, -50, -25, -7, -12,
    -- layer=1 filter=91 channel=119
    -4, -10, -28, 11, 14, -22, 31, 58, 7,
    -- layer=1 filter=91 channel=120
    -14, -25, -13, -21, 30, 27, -10, 32, 16,
    -- layer=1 filter=91 channel=121
    -49, -35, -26, -23, -41, -51, -40, -8, -52,
    -- layer=1 filter=91 channel=122
    9, -1, 6, -9, -9, 10, 4, -3, 0,
    -- layer=1 filter=91 channel=123
    -34, -32, -24, -37, -10, -46, -46, 6, -41,
    -- layer=1 filter=91 channel=124
    25, -12, 28, 17, -2, 26, -10, 9, -11,
    -- layer=1 filter=91 channel=125
    18, 26, 9, 0, 9, 22, 5, 38, 44,
    -- layer=1 filter=91 channel=126
    -48, -91, -37, -40, 0, 48, -13, 35, 3,
    -- layer=1 filter=91 channel=127
    -35, 9, -14, -30, -28, -47, -27, -27, -35,
    -- layer=1 filter=92 channel=0
    5, 2, -7, 6, 1, 4, -1, 2, -7,
    -- layer=1 filter=92 channel=1
    1, 6, 0, -12, -1, -4, -12, 2, -10,
    -- layer=1 filter=92 channel=2
    -6, -3, -6, 3, -4, -3, 1, 7, -9,
    -- layer=1 filter=92 channel=3
    9, 6, -1, 6, -5, -7, -9, 4, 4,
    -- layer=1 filter=92 channel=4
    0, -1, 1, 6, -2, 5, 1, 0, -8,
    -- layer=1 filter=92 channel=5
    -3, -3, -9, -3, 8, 6, -1, -2, -11,
    -- layer=1 filter=92 channel=6
    -10, -6, -10, -3, 5, 2, -9, -1, 1,
    -- layer=1 filter=92 channel=7
    -9, 5, -8, 7, -7, -2, -4, -8, 4,
    -- layer=1 filter=92 channel=8
    0, -11, 3, 7, -1, 0, 0, -7, 3,
    -- layer=1 filter=92 channel=9
    7, -6, 0, -5, 4, 5, 11, 0, 11,
    -- layer=1 filter=92 channel=10
    -5, 2, 7, -6, 1, -1, 3, -10, -6,
    -- layer=1 filter=92 channel=11
    -2, 0, -1, -6, 0, -9, 7, 3, -4,
    -- layer=1 filter=92 channel=12
    4, -9, 4, 8, 6, -3, 3, 0, 9,
    -- layer=1 filter=92 channel=13
    1, -5, -1, -4, -1, 7, -12, -11, 1,
    -- layer=1 filter=92 channel=14
    -1, -8, -5, 2, 6, -10, 3, 2, 7,
    -- layer=1 filter=92 channel=15
    0, -4, -11, -9, 7, 9, 7, -11, 4,
    -- layer=1 filter=92 channel=16
    1, -3, 4, -10, -1, -9, -3, -1, -2,
    -- layer=1 filter=92 channel=17
    0, 0, -11, 2, -2, -5, -8, -8, 5,
    -- layer=1 filter=92 channel=18
    -6, -7, -9, 4, 0, -7, 11, 0, -2,
    -- layer=1 filter=92 channel=19
    1, -1, -3, 3, -4, 3, -8, -3, 4,
    -- layer=1 filter=92 channel=20
    0, -4, -4, 3, 4, 7, -12, 0, -2,
    -- layer=1 filter=92 channel=21
    0, 10, 6, 0, -5, -6, -9, -8, -6,
    -- layer=1 filter=92 channel=22
    5, -10, 1, -5, 0, 4, -12, -8, 1,
    -- layer=1 filter=92 channel=23
    -3, 2, 6, 1, 5, 1, 3, 7, 1,
    -- layer=1 filter=92 channel=24
    -5, 6, -5, 8, -1, -4, 8, 0, 3,
    -- layer=1 filter=92 channel=25
    5, -2, 2, -2, 3, -10, -5, 1, 0,
    -- layer=1 filter=92 channel=26
    6, 7, 0, 5, 6, 0, 1, 0, 4,
    -- layer=1 filter=92 channel=27
    6, -2, -4, -6, -2, -9, -7, 3, 7,
    -- layer=1 filter=92 channel=28
    2, -8, 0, 3, -5, -4, -11, -4, 4,
    -- layer=1 filter=92 channel=29
    -6, 9, 9, 3, -6, 5, 3, -3, -6,
    -- layer=1 filter=92 channel=30
    -5, -2, 4, 5, -10, -3, -11, -7, -2,
    -- layer=1 filter=92 channel=31
    -3, -10, 0, 0, -12, 0, 4, -11, -9,
    -- layer=1 filter=92 channel=32
    3, 1, 0, -5, 4, 0, -6, 0, -7,
    -- layer=1 filter=92 channel=33
    5, -4, 11, -5, 2, -6, 10, 3, 1,
    -- layer=1 filter=92 channel=34
    -5, 0, -8, 1, -4, 1, 8, 6, 1,
    -- layer=1 filter=92 channel=35
    -10, -11, -10, 8, -4, -6, -8, 1, -1,
    -- layer=1 filter=92 channel=36
    -8, 6, -7, 5, -2, -7, 0, 8, -5,
    -- layer=1 filter=92 channel=37
    0, -9, -8, 0, -7, -3, -2, -11, -2,
    -- layer=1 filter=92 channel=38
    0, 0, 1, -3, -6, 0, 5, -2, 1,
    -- layer=1 filter=92 channel=39
    -3, -10, 0, -1, 1, 0, -11, -12, 0,
    -- layer=1 filter=92 channel=40
    2, -7, -3, -8, -7, -8, 3, -8, -1,
    -- layer=1 filter=92 channel=41
    -8, 4, -7, -1, -11, -6, 1, -1, -3,
    -- layer=1 filter=92 channel=42
    1, 9, -1, -9, 2, 5, 6, -8, 4,
    -- layer=1 filter=92 channel=43
    -4, 0, 0, -1, 6, -1, 4, 2, 6,
    -- layer=1 filter=92 channel=44
    -3, -6, 2, -11, -9, 3, 6, -6, -7,
    -- layer=1 filter=92 channel=45
    4, 2, -10, -5, 2, 3, 2, 8, 2,
    -- layer=1 filter=92 channel=46
    7, 8, 9, 3, -2, -1, 10, 4, 10,
    -- layer=1 filter=92 channel=47
    -5, -10, -6, -2, -8, -6, -12, -1, 7,
    -- layer=1 filter=92 channel=48
    -1, 0, 0, -9, -3, 1, 0, 7, 1,
    -- layer=1 filter=92 channel=49
    -12, 8, 0, 0, 4, -9, 1, -9, -1,
    -- layer=1 filter=92 channel=50
    3, -9, -8, 7, -7, 0, -8, -6, -5,
    -- layer=1 filter=92 channel=51
    0, -8, 2, -7, 0, 1, -11, 2, 9,
    -- layer=1 filter=92 channel=52
    -5, -7, -2, 11, 3, -2, 2, 0, -6,
    -- layer=1 filter=92 channel=53
    -3, -12, -4, 0, -1, 2, -8, -10, -4,
    -- layer=1 filter=92 channel=54
    -5, -7, 7, 0, -6, -11, -7, 0, -2,
    -- layer=1 filter=92 channel=55
    -1, -11, -11, 4, -9, -4, 0, 3, -6,
    -- layer=1 filter=92 channel=56
    0, 0, -10, -4, -1, 2, -10, 4, -2,
    -- layer=1 filter=92 channel=57
    2, -1, -6, 5, 0, -6, 0, 2, 3,
    -- layer=1 filter=92 channel=58
    6, -1, -1, -7, -9, -4, 4, -9, 0,
    -- layer=1 filter=92 channel=59
    -5, -7, -1, -5, -5, -9, 2, -4, 5,
    -- layer=1 filter=92 channel=60
    5, 0, 2, -11, -7, 0, 4, -8, -5,
    -- layer=1 filter=92 channel=61
    -11, 2, 0, -10, 4, 5, -2, -5, 6,
    -- layer=1 filter=92 channel=62
    -2, -5, -12, 9, 2, -5, 8, 2, 7,
    -- layer=1 filter=92 channel=63
    -7, -3, -10, 4, 4, -5, -4, 5, 1,
    -- layer=1 filter=92 channel=64
    -6, 7, 1, -9, 1, -8, 0, -11, 7,
    -- layer=1 filter=92 channel=65
    -12, 7, 1, -8, -6, -3, -7, -11, 1,
    -- layer=1 filter=92 channel=66
    -4, -2, -1, -2, -5, -8, -11, -6, 0,
    -- layer=1 filter=92 channel=67
    1, -8, 8, 7, -4, 8, 9, -3, 3,
    -- layer=1 filter=92 channel=68
    1, -11, -7, -11, 5, 0, 0, -11, -3,
    -- layer=1 filter=92 channel=69
    7, 6, 8, 3, 0, -8, 9, -3, 7,
    -- layer=1 filter=92 channel=70
    0, 1, 0, -7, -1, 5, 9, -1, -2,
    -- layer=1 filter=92 channel=71
    3, 4, 1, -10, -8, 2, -9, -9, 0,
    -- layer=1 filter=92 channel=72
    5, -8, 3, -3, 3, -12, -6, 5, 3,
    -- layer=1 filter=92 channel=73
    -2, 1, 0, -9, 2, -1, 6, 8, -8,
    -- layer=1 filter=92 channel=74
    4, 7, 0, -5, 6, 0, 2, -2, 7,
    -- layer=1 filter=92 channel=75
    1, -6, -8, -7, -10, -5, -6, 8, 8,
    -- layer=1 filter=92 channel=76
    2, 1, -2, 4, 2, 6, 7, 7, 6,
    -- layer=1 filter=92 channel=77
    -9, -7, 4, -1, 5, -4, -6, -8, 2,
    -- layer=1 filter=92 channel=78
    -5, -1, 2, 7, 0, -11, -10, -2, -9,
    -- layer=1 filter=92 channel=79
    -9, -9, -7, -5, -8, 0, -9, -5, 7,
    -- layer=1 filter=92 channel=80
    7, -5, -9, -6, 1, 0, -2, 0, 3,
    -- layer=1 filter=92 channel=81
    1, -5, 8, -10, -10, 2, -5, -8, -9,
    -- layer=1 filter=92 channel=82
    -7, 6, 0, -6, -1, 0, -3, 0, 3,
    -- layer=1 filter=92 channel=83
    6, 0, 2, 6, 0, 7, -5, -10, 0,
    -- layer=1 filter=92 channel=84
    6, -10, 2, -5, -5, 1, 6, 6, -2,
    -- layer=1 filter=92 channel=85
    0, -6, 2, -7, 0, 7, -3, 0, -4,
    -- layer=1 filter=92 channel=86
    0, 8, 8, -8, 0, -10, 0, 0, -2,
    -- layer=1 filter=92 channel=87
    -5, 2, 6, -3, -5, -4, 2, -7, 0,
    -- layer=1 filter=92 channel=88
    5, 4, 6, 5, 6, 11, -4, 1, -4,
    -- layer=1 filter=92 channel=89
    1, -3, 4, -4, -2, -10, 5, -5, -7,
    -- layer=1 filter=92 channel=90
    -8, -1, -11, 6, -4, 6, 4, 1, 4,
    -- layer=1 filter=92 channel=91
    4, -9, -8, -11, -5, -7, -10, 1, -4,
    -- layer=1 filter=92 channel=92
    -4, 3, 1, 7, -10, 0, 1, -9, 3,
    -- layer=1 filter=92 channel=93
    -1, -9, -1, -8, 4, 0, -2, -11, 8,
    -- layer=1 filter=92 channel=94
    -1, -7, -7, -1, -2, 0, -4, 2, 4,
    -- layer=1 filter=92 channel=95
    -7, -4, 3, -5, -11, -10, 11, -5, 0,
    -- layer=1 filter=92 channel=96
    -8, -10, 0, 7, -7, -2, 6, 0, 4,
    -- layer=1 filter=92 channel=97
    7, 1, -7, 4, -6, -5, 1, -9, 2,
    -- layer=1 filter=92 channel=98
    -2, 3, -7, 0, 8, -8, -1, 6, 0,
    -- layer=1 filter=92 channel=99
    -5, -9, -12, 5, -3, -1, -4, 7, 6,
    -- layer=1 filter=92 channel=100
    -2, -2, 6, 2, -1, -12, 5, -5, 1,
    -- layer=1 filter=92 channel=101
    -1, -10, 3, 1, -12, 7, 1, -9, 5,
    -- layer=1 filter=92 channel=102
    -9, -3, -5, 7, -3, 7, -6, 0, -6,
    -- layer=1 filter=92 channel=103
    2, -6, 6, -3, -7, 2, 0, 7, -6,
    -- layer=1 filter=92 channel=104
    -5, 2, -3, -5, 6, 3, -4, -8, -4,
    -- layer=1 filter=92 channel=105
    -8, 1, -11, -11, 7, 6, 1, -11, -13,
    -- layer=1 filter=92 channel=106
    2, 6, -4, -9, 7, -7, -4, -12, -7,
    -- layer=1 filter=92 channel=107
    2, -2, -4, -3, 7, -10, 2, -3, -8,
    -- layer=1 filter=92 channel=108
    6, -7, 8, 5, -9, 0, -6, -7, -10,
    -- layer=1 filter=92 channel=109
    4, -3, -6, -2, 5, 6, -6, -8, 0,
    -- layer=1 filter=92 channel=110
    7, -8, -3, 4, 4, 0, -12, 1, -11,
    -- layer=1 filter=92 channel=111
    7, 5, -6, 3, 5, -2, 1, -6, 0,
    -- layer=1 filter=92 channel=112
    -4, -10, -9, -9, 0, -4, -10, -1, -10,
    -- layer=1 filter=92 channel=113
    -7, 0, -1, 6, -4, 0, 4, 3, -11,
    -- layer=1 filter=92 channel=114
    3, -10, -9, 2, -8, -4, 2, 1, -3,
    -- layer=1 filter=92 channel=115
    -8, -1, -7, 2, -12, 1, 1, -3, 0,
    -- layer=1 filter=92 channel=116
    -5, 0, -5, 2, -2, -7, 4, -10, 6,
    -- layer=1 filter=92 channel=117
    -1, 4, -2, 5, -7, 6, 10, 1, 2,
    -- layer=1 filter=92 channel=118
    0, 0, 0, 6, -6, -2, -7, 0, 6,
    -- layer=1 filter=92 channel=119
    -2, 5, -1, 0, -1, 0, 0, -9, 0,
    -- layer=1 filter=92 channel=120
    -8, 3, -6, 8, -1, -8, 1, -8, 5,
    -- layer=1 filter=92 channel=121
    -5, 5, 9, 7, -2, -9, -6, 5, -6,
    -- layer=1 filter=92 channel=122
    6, 0, 2, 4, -3, 10, 7, 9, -7,
    -- layer=1 filter=92 channel=123
    -8, -10, 2, 5, 0, 0, 7, 2, 4,
    -- layer=1 filter=92 channel=124
    8, -10, -1, -5, -2, -5, -8, -3, -4,
    -- layer=1 filter=92 channel=125
    -4, 10, 6, 8, 2, -8, 7, -1, 0,
    -- layer=1 filter=92 channel=126
    -6, 0, -9, -5, 2, 8, 2, -7, 1,
    -- layer=1 filter=92 channel=127
    -5, -4, -8, -6, -7, -2, -2, -12, 8,
    -- layer=1 filter=93 channel=0
    -10, 5, -3, 1, 3, -6, -9, -2, 1,
    -- layer=1 filter=93 channel=1
    2, 5, -6, -3, -2, -7, 0, 3, -3,
    -- layer=1 filter=93 channel=2
    8, 7, 3, -6, 4, 2, 7, -8, -6,
    -- layer=1 filter=93 channel=3
    3, -3, 4, -8, 2, -1, -10, -6, -9,
    -- layer=1 filter=93 channel=4
    -10, -10, -9, 4, -10, 0, 1, -1, 4,
    -- layer=1 filter=93 channel=5
    5, -3, -3, 6, 3, 4, 0, -1, -7,
    -- layer=1 filter=93 channel=6
    -7, -3, 8, 0, -8, 0, -8, 5, -5,
    -- layer=1 filter=93 channel=7
    -8, 6, -2, 6, 4, -13, -7, 0, 4,
    -- layer=1 filter=93 channel=8
    -6, -8, 1, -3, -2, -7, -5, 2, 6,
    -- layer=1 filter=93 channel=9
    -11, -14, -7, -5, -2, -11, -1, -6, -9,
    -- layer=1 filter=93 channel=10
    7, 4, -9, -10, -9, -4, 6, 0, -11,
    -- layer=1 filter=93 channel=11
    -2, 1, -5, -8, 2, 6, 2, -1, -5,
    -- layer=1 filter=93 channel=12
    2, 1, -8, -1, 5, 6, -7, 4, -7,
    -- layer=1 filter=93 channel=13
    4, 8, 4, -4, 7, -6, -7, 0, 0,
    -- layer=1 filter=93 channel=14
    4, 8, -8, -10, -10, -2, 8, 0, -8,
    -- layer=1 filter=93 channel=15
    -11, -5, 8, 4, -9, -8, -3, 2, -5,
    -- layer=1 filter=93 channel=16
    8, -3, -9, -8, 4, 7, 8, -6, 0,
    -- layer=1 filter=93 channel=17
    6, 3, -2, 0, 3, 5, 2, 3, 4,
    -- layer=1 filter=93 channel=18
    -3, 2, 4, 7, 6, -1, 8, -8, 5,
    -- layer=1 filter=93 channel=19
    7, 0, 5, -2, -7, 1, 1, 6, -6,
    -- layer=1 filter=93 channel=20
    6, 0, 2, -3, -2, 0, 6, 2, 8,
    -- layer=1 filter=93 channel=21
    4, -8, -7, -12, -4, -10, 7, -9, -10,
    -- layer=1 filter=93 channel=22
    5, -10, 8, 0, -5, 0, -3, 7, -10,
    -- layer=1 filter=93 channel=23
    -2, 0, 0, 2, -7, 8, -6, -5, -2,
    -- layer=1 filter=93 channel=24
    1, -3, -6, -8, 0, -6, -7, 0, 5,
    -- layer=1 filter=93 channel=25
    5, -3, 0, -11, 10, -2, -4, -5, 0,
    -- layer=1 filter=93 channel=26
    -5, -10, -12, -5, 6, -4, -2, -10, -6,
    -- layer=1 filter=93 channel=27
    -3, -7, 0, 0, -4, -3, -1, 4, -11,
    -- layer=1 filter=93 channel=28
    3, 0, -11, 5, 0, -8, 8, 0, 6,
    -- layer=1 filter=93 channel=29
    2, 2, -5, 1, -6, -9, -4, 5, 2,
    -- layer=1 filter=93 channel=30
    -7, 4, -5, 6, -2, -7, -7, 8, 6,
    -- layer=1 filter=93 channel=31
    -11, 6, -11, -4, 7, -6, 5, -11, -5,
    -- layer=1 filter=93 channel=32
    -6, 2, 9, 3, -3, 5, -6, 5, -6,
    -- layer=1 filter=93 channel=33
    0, 9, -9, 8, -4, 3, 1, 3, 3,
    -- layer=1 filter=93 channel=34
    -11, -3, 8, 3, -2, 0, 7, -6, 3,
    -- layer=1 filter=93 channel=35
    -8, 1, -7, 2, -9, 4, -8, -3, 5,
    -- layer=1 filter=93 channel=36
    2, 5, -7, 1, -3, -5, -5, -2, 7,
    -- layer=1 filter=93 channel=37
    -5, 7, -11, 1, -12, -8, 3, -12, 3,
    -- layer=1 filter=93 channel=38
    -6, 0, -6, -11, -1, -12, -11, -12, -7,
    -- layer=1 filter=93 channel=39
    8, 8, 1, -1, 8, -5, 6, -1, 0,
    -- layer=1 filter=93 channel=40
    -5, -8, -2, 3, -4, 8, -8, -2, 0,
    -- layer=1 filter=93 channel=41
    9, -6, 1, -10, 7, 9, 7, 0, 5,
    -- layer=1 filter=93 channel=42
    -5, 6, 3, 0, 9, 3, 8, 0, 6,
    -- layer=1 filter=93 channel=43
    -5, 7, -6, 8, -7, -2, -9, 9, 3,
    -- layer=1 filter=93 channel=44
    -9, -9, -6, 3, -7, 9, 6, -4, 5,
    -- layer=1 filter=93 channel=45
    -3, 7, 0, -9, 5, 0, 4, -1, 6,
    -- layer=1 filter=93 channel=46
    -4, 9, 1, 4, -10, 7, 2, 9, 8,
    -- layer=1 filter=93 channel=47
    -6, 3, -9, -11, -5, -4, -13, -4, -7,
    -- layer=1 filter=93 channel=48
    3, -1, -8, -11, -3, -8, 7, -7, 2,
    -- layer=1 filter=93 channel=49
    7, -7, -4, -10, -11, 4, 2, 6, 3,
    -- layer=1 filter=93 channel=50
    -3, -4, 6, -1, -2, -6, 0, 4, -2,
    -- layer=1 filter=93 channel=51
    -1, 7, -4, -11, -2, 7, -1, 4, 0,
    -- layer=1 filter=93 channel=52
    1, 0, 0, 9, 2, 0, 8, -5, 6,
    -- layer=1 filter=93 channel=53
    5, 0, -4, -10, -4, 2, -2, -3, 7,
    -- layer=1 filter=93 channel=54
    4, -3, 8, 0, 9, -4, -4, 6, 1,
    -- layer=1 filter=93 channel=55
    -6, 2, 7, -2, -2, -5, -10, 1, -2,
    -- layer=1 filter=93 channel=56
    6, -11, 8, 1, 1, -2, 7, -8, -9,
    -- layer=1 filter=93 channel=57
    5, 3, -8, 2, -7, 0, -7, 0, -8,
    -- layer=1 filter=93 channel=58
    -9, -12, 7, -9, -8, -5, -4, 0, 6,
    -- layer=1 filter=93 channel=59
    8, 2, -7, -4, -5, -6, -11, 8, 10,
    -- layer=1 filter=93 channel=60
    1, -7, 8, -10, 1, 2, 7, -4, 1,
    -- layer=1 filter=93 channel=61
    4, -5, 1, -10, -3, -5, -10, -4, -8,
    -- layer=1 filter=93 channel=62
    0, 0, -3, 5, 7, -1, -5, -10, -12,
    -- layer=1 filter=93 channel=63
    -11, 5, 1, -8, 2, 5, 3, -1, 7,
    -- layer=1 filter=93 channel=64
    3, 2, -1, 0, -4, 0, 3, 6, 6,
    -- layer=1 filter=93 channel=65
    -4, 3, 7, 0, 0, -3, 1, 6, 1,
    -- layer=1 filter=93 channel=66
    7, 6, -4, -5, -5, 5, -4, -8, 7,
    -- layer=1 filter=93 channel=67
    9, 6, -7, -5, -6, 8, 1, -3, -6,
    -- layer=1 filter=93 channel=68
    -7, 0, -1, -9, -2, 4, 5, -5, 9,
    -- layer=1 filter=93 channel=69
    -1, 2, -10, -7, 3, -2, -12, -7, -7,
    -- layer=1 filter=93 channel=70
    -7, -8, 3, -7, -7, 3, 4, -9, 1,
    -- layer=1 filter=93 channel=71
    6, -4, 5, 4, -13, -6, 5, 2, -9,
    -- layer=1 filter=93 channel=72
    3, -10, -13, 4, 6, 7, 6, -5, -7,
    -- layer=1 filter=93 channel=73
    0, -9, -4, 0, -10, 3, -5, -6, 6,
    -- layer=1 filter=93 channel=74
    9, -3, 0, -3, -1, -1, 4, 7, 2,
    -- layer=1 filter=93 channel=75
    -6, 4, 1, 2, 5, -10, 1, 7, 15,
    -- layer=1 filter=93 channel=76
    4, -1, -1, 1, -2, -9, 4, 1, 4,
    -- layer=1 filter=93 channel=77
    -11, -11, 4, -4, -2, -8, -3, -12, -7,
    -- layer=1 filter=93 channel=78
    -7, -8, -10, 8, 0, -2, -9, -6, 4,
    -- layer=1 filter=93 channel=79
    -3, -12, 7, 7, -2, -7, 3, -3, -9,
    -- layer=1 filter=93 channel=80
    -10, -3, 7, -9, -2, 6, -1, 0, -8,
    -- layer=1 filter=93 channel=81
    5, -10, 5, 2, -7, -4, 0, 6, 6,
    -- layer=1 filter=93 channel=82
    0, 3, 4, -10, -10, -6, -3, 7, -6,
    -- layer=1 filter=93 channel=83
    -3, -7, 6, -5, 9, -2, 4, 3, 8,
    -- layer=1 filter=93 channel=84
    8, -1, -13, -5, 6, -8, -6, 9, -2,
    -- layer=1 filter=93 channel=85
    -3, 3, 7, -6, 4, -9, -1, 7, 10,
    -- layer=1 filter=93 channel=86
    -9, -12, 4, 8, -11, 0, -8, -3, 3,
    -- layer=1 filter=93 channel=87
    -2, 10, 7, -9, -5, -7, 2, 0, 1,
    -- layer=1 filter=93 channel=88
    -12, -5, -4, -3, -3, 4, -2, 4, 3,
    -- layer=1 filter=93 channel=89
    -8, -9, -2, -6, 0, -4, -4, -7, -8,
    -- layer=1 filter=93 channel=90
    -9, -3, 0, -1, 3, -10, 1, -11, -7,
    -- layer=1 filter=93 channel=91
    -3, -12, -6, -8, 5, 2, -9, 4, -3,
    -- layer=1 filter=93 channel=92
    5, 4, -9, -2, -4, 2, 8, -7, -2,
    -- layer=1 filter=93 channel=93
    -10, -8, 0, -1, 0, 1, 0, -7, -1,
    -- layer=1 filter=93 channel=94
    -8, 0, -1, -6, 3, 1, 5, -10, 8,
    -- layer=1 filter=93 channel=95
    -3, 4, -12, 0, 5, -8, -3, 7, 0,
    -- layer=1 filter=93 channel=96
    -5, 7, -7, 0, 1, -11, -11, -6, -4,
    -- layer=1 filter=93 channel=97
    -9, -12, 0, 0, 7, 4, -12, 3, 1,
    -- layer=1 filter=93 channel=98
    0, -7, 2, -2, -6, 6, 0, 0, 0,
    -- layer=1 filter=93 channel=99
    6, 2, -6, -6, 0, 3, -10, 0, 0,
    -- layer=1 filter=93 channel=100
    -9, -7, 4, -7, -9, 5, -1, -10, 3,
    -- layer=1 filter=93 channel=101
    -10, -7, -7, 0, -1, -2, 3, -11, -9,
    -- layer=1 filter=93 channel=102
    -8, -5, 1, -9, -6, 5, -7, -7, -4,
    -- layer=1 filter=93 channel=103
    7, 7, 8, 4, 5, 0, 9, -6, -9,
    -- layer=1 filter=93 channel=104
    -4, 0, -1, 8, -10, -8, 1, -3, 0,
    -- layer=1 filter=93 channel=105
    -9, 5, -9, 8, -1, -11, -8, 1, -6,
    -- layer=1 filter=93 channel=106
    -11, -6, 0, -8, 9, -11, 0, -7, -2,
    -- layer=1 filter=93 channel=107
    5, -6, 0, -10, -4, 6, -7, -4, 8,
    -- layer=1 filter=93 channel=108
    -3, -6, -6, -7, -1, 8, -2, 6, 3,
    -- layer=1 filter=93 channel=109
    -4, -1, 8, -7, -8, 7, 7, 2, -6,
    -- layer=1 filter=93 channel=110
    -2, -6, -10, -10, 1, -3, -5, -9, 5,
    -- layer=1 filter=93 channel=111
    8, -2, -8, 1, -6, -7, -7, -4, 4,
    -- layer=1 filter=93 channel=112
    -6, 3, 8, 0, -1, -5, -5, 1, -8,
    -- layer=1 filter=93 channel=113
    -5, 6, -7, 5, -8, -9, -10, -9, 0,
    -- layer=1 filter=93 channel=114
    -14, 0, -16, -13, 0, -9, -3, 0, -17,
    -- layer=1 filter=93 channel=115
    -5, 6, 4, 3, -3, -8, -3, 6, -11,
    -- layer=1 filter=93 channel=116
    -1, -6, 8, -1, 7, 2, -4, 3, -1,
    -- layer=1 filter=93 channel=117
    -3, 3, -1, -7, 2, -9, 3, 0, 10,
    -- layer=1 filter=93 channel=118
    -5, -5, 7, -9, -8, -6, -4, -7, 8,
    -- layer=1 filter=93 channel=119
    -8, 5, 0, -6, 1, -2, -3, 3, -10,
    -- layer=1 filter=93 channel=120
    4, -3, -10, 4, 0, 7, 0, -5, 4,
    -- layer=1 filter=93 channel=121
    5, 5, 0, -1, -7, -6, 1, -1, -2,
    -- layer=1 filter=93 channel=122
    0, 4, 7, -3, 4, 10, 5, 8, 3,
    -- layer=1 filter=93 channel=123
    -3, 5, -8, 4, 6, -12, 5, 0, -1,
    -- layer=1 filter=93 channel=124
    -8, -8, 0, 0, 5, -3, 7, 4, -7,
    -- layer=1 filter=93 channel=125
    -7, 3, 8, -5, 7, -3, 4, -3, -9,
    -- layer=1 filter=93 channel=126
    -8, -8, -7, -6, 4, 8, 0, 9, -4,
    -- layer=1 filter=93 channel=127
    4, -3, 3, -3, -12, -13, -4, -4, 2,
    -- layer=1 filter=94 channel=0
    1, 6, 5, 3, 4, 5, -8, -2, -8,
    -- layer=1 filter=94 channel=1
    3, -2, 3, -6, -8, 0, -5, -5, -4,
    -- layer=1 filter=94 channel=2
    -12, 2, -6, -14, -4, -12, -5, -7, 2,
    -- layer=1 filter=94 channel=3
    0, -2, -7, -10, 5, -5, 9, -7, 0,
    -- layer=1 filter=94 channel=4
    -5, 3, 3, 5, 0, -1, -1, 9, 5,
    -- layer=1 filter=94 channel=5
    7, 1, 6, -7, -10, -2, -1, 5, 1,
    -- layer=1 filter=94 channel=6
    -1, 9, -6, -9, 0, -5, 8, -4, -6,
    -- layer=1 filter=94 channel=7
    0, 2, -9, -11, 0, -8, 3, -9, 0,
    -- layer=1 filter=94 channel=8
    9, -9, 4, -3, 1, -1, -4, -8, 1,
    -- layer=1 filter=94 channel=9
    0, 1, -4, -3, 5, 5, 9, -3, 5,
    -- layer=1 filter=94 channel=10
    8, -2, 1, -6, -7, 2, -12, 2, -5,
    -- layer=1 filter=94 channel=11
    -7, -4, -5, 0, -7, -13, 2, 2, -12,
    -- layer=1 filter=94 channel=12
    7, -8, 0, 10, -5, -5, 2, 7, 7,
    -- layer=1 filter=94 channel=13
    -11, 3, -8, -3, 0, -1, 3, 2, -7,
    -- layer=1 filter=94 channel=14
    5, -12, 0, -9, -2, -12, -5, 5, -11,
    -- layer=1 filter=94 channel=15
    4, 4, 9, -10, -2, -9, 6, -11, 0,
    -- layer=1 filter=94 channel=16
    -2, -7, -10, -4, 0, 0, 0, 3, -7,
    -- layer=1 filter=94 channel=17
    -8, 0, 6, -10, 0, -4, 0, 2, -7,
    -- layer=1 filter=94 channel=18
    -14, 0, 1, 3, -4, 2, -7, 0, -1,
    -- layer=1 filter=94 channel=19
    2, 3, -6, 7, 8, -8, -1, 3, -10,
    -- layer=1 filter=94 channel=20
    4, -8, -2, -2, 6, -1, -8, 3, -4,
    -- layer=1 filter=94 channel=21
    -5, 6, -6, 4, 0, -9, -13, 2, -5,
    -- layer=1 filter=94 channel=22
    2, 0, 9, -7, 2, 7, 4, 1, 9,
    -- layer=1 filter=94 channel=23
    -5, 2, 2, -7, 0, -1, -3, -3, -7,
    -- layer=1 filter=94 channel=24
    0, -12, -8, -14, 4, 3, -6, 0, 3,
    -- layer=1 filter=94 channel=25
    -2, 4, 4, -7, 0, -11, -5, -5, -4,
    -- layer=1 filter=94 channel=26
    -2, 4, 0, 0, -14, 2, -13, 1, -3,
    -- layer=1 filter=94 channel=27
    -4, 2, -8, -14, -10, -2, 3, -4, -2,
    -- layer=1 filter=94 channel=28
    -2, -8, -7, -4, 0, -2, -8, -1, 7,
    -- layer=1 filter=94 channel=29
    -4, 3, -9, -8, -5, 9, -1, 2, -2,
    -- layer=1 filter=94 channel=30
    -7, -7, 1, -4, 3, -6, 9, -6, -3,
    -- layer=1 filter=94 channel=31
    -14, 3, -7, -14, -13, -14, -8, -14, -10,
    -- layer=1 filter=94 channel=32
    2, -1, -7, -2, -1, 4, 5, 7, 1,
    -- layer=1 filter=94 channel=33
    2, 10, 1, 5, 9, -1, -3, 8, -2,
    -- layer=1 filter=94 channel=34
    7, -4, 4, 2, 3, -7, -9, 2, 0,
    -- layer=1 filter=94 channel=35
    0, 2, -4, 1, 0, 1, 0, 4, 6,
    -- layer=1 filter=94 channel=36
    -10, 0, 1, -11, -3, 0, -10, -13, -16,
    -- layer=1 filter=94 channel=37
    1, -1, -7, -4, -9, 5, 1, 2, -8,
    -- layer=1 filter=94 channel=38
    -1, -6, -5, -3, 2, -11, 0, -11, -6,
    -- layer=1 filter=94 channel=39
    3, -11, -5, 0, -4, 0, 2, -6, -2,
    -- layer=1 filter=94 channel=40
    3, -4, 5, 0, 6, -8, -2, 3, 1,
    -- layer=1 filter=94 channel=41
    0, -8, -12, -11, 6, 6, -2, 4, 0,
    -- layer=1 filter=94 channel=42
    0, -4, 2, -1, -1, 0, -2, -4, -11,
    -- layer=1 filter=94 channel=43
    8, 2, 10, 0, 2, 0, -3, -1, 7,
    -- layer=1 filter=94 channel=44
    -4, 6, -6, -5, -10, -10, -6, -1, 1,
    -- layer=1 filter=94 channel=45
    4, -8, -5, -4, 3, 0, -5, 7, -9,
    -- layer=1 filter=94 channel=46
    -4, 4, -5, 0, -5, -6, -4, 5, -3,
    -- layer=1 filter=94 channel=47
    -1, -10, 9, 5, -3, -9, -2, 4, -8,
    -- layer=1 filter=94 channel=48
    6, -6, 4, 8, -9, 3, -9, -10, -3,
    -- layer=1 filter=94 channel=49
    1, -3, 0, 2, -8, 8, 0, -1, 2,
    -- layer=1 filter=94 channel=50
    -4, 3, 2, -6, 0, 2, -6, 10, -9,
    -- layer=1 filter=94 channel=51
    -3, 10, 7, -11, -1, -4, -5, -9, -3,
    -- layer=1 filter=94 channel=52
    4, 7, 1, -7, 0, -8, 4, 0, 4,
    -- layer=1 filter=94 channel=53
    0, 5, 10, 9, 0, -1, 0, 1, -10,
    -- layer=1 filter=94 channel=54
    -11, -1, -7, -3, -6, -2, -11, -15, 2,
    -- layer=1 filter=94 channel=55
    -6, -8, 2, -2, -2, 2, 3, -17, -1,
    -- layer=1 filter=94 channel=56
    -10, 3, -4, -4, -3, -7, 2, 3, -6,
    -- layer=1 filter=94 channel=57
    -11, 0, -8, 1, -4, 0, 2, -14, 3,
    -- layer=1 filter=94 channel=58
    1, -12, -4, 7, 6, -4, -3, -3, -7,
    -- layer=1 filter=94 channel=59
    -10, 3, 8, 7, -4, 2, 1, -9, 3,
    -- layer=1 filter=94 channel=60
    -4, 1, 1, 10, 4, 4, 3, -5, 1,
    -- layer=1 filter=94 channel=61
    -10, 1, 6, -5, -8, -8, 5, 3, -8,
    -- layer=1 filter=94 channel=62
    1, -9, -2, -6, -2, 6, 6, 2, 8,
    -- layer=1 filter=94 channel=63
    2, -17, -16, 3, 0, -2, -1, 3, 4,
    -- layer=1 filter=94 channel=64
    0, -1, 8, 5, -3, 5, 4, 4, 1,
    -- layer=1 filter=94 channel=65
    5, -1, 2, 0, -1, 0, 3, 3, 3,
    -- layer=1 filter=94 channel=66
    -2, -8, -5, 0, -7, -14, 5, 0, -4,
    -- layer=1 filter=94 channel=67
    3, 0, 4, -1, 5, -9, -7, -10, 10,
    -- layer=1 filter=94 channel=68
    -9, -3, -4, -1, -2, 2, -2, 6, -4,
    -- layer=1 filter=94 channel=69
    -11, 6, -11, -1, -12, 0, -2, -8, -7,
    -- layer=1 filter=94 channel=70
    -4, 0, 9, 4, 0, 6, 4, 3, 0,
    -- layer=1 filter=94 channel=71
    -8, -10, 0, 5, 5, 9, 1, -5, -5,
    -- layer=1 filter=94 channel=72
    0, -6, -12, -10, -7, -4, 0, 6, 7,
    -- layer=1 filter=94 channel=73
    -8, -5, 1, 4, 4, 3, 0, 1, -4,
    -- layer=1 filter=94 channel=74
    -3, -5, -4, -9, 5, -8, 5, 7, -2,
    -- layer=1 filter=94 channel=75
    -6, -5, 1, 1, -8, -1, -2, -2, 4,
    -- layer=1 filter=94 channel=76
    8, -6, -1, -8, -4, -1, -7, 10, -2,
    -- layer=1 filter=94 channel=77
    8, -5, 5, -1, -4, -3, 3, 8, 4,
    -- layer=1 filter=94 channel=78
    0, -4, -1, -2, -9, -6, 7, 3, -6,
    -- layer=1 filter=94 channel=79
    -6, 6, 8, -4, 4, -7, -11, 0, -5,
    -- layer=1 filter=94 channel=80
    -10, 7, 5, -4, 0, 5, 7, 1, 9,
    -- layer=1 filter=94 channel=81
    -8, -8, -10, -5, -11, -3, 0, 0, 4,
    -- layer=1 filter=94 channel=82
    -1, 10, 7, 5, -5, -9, 4, 1, -9,
    -- layer=1 filter=94 channel=83
    -3, 3, 0, -3, -7, 5, 3, -8, -1,
    -- layer=1 filter=94 channel=84
    -12, -5, 3, -10, -7, -7, 6, -13, -7,
    -- layer=1 filter=94 channel=85
    3, -2, 0, 3, -3, -10, -8, -1, -11,
    -- layer=1 filter=94 channel=86
    2, -13, 2, -6, -10, -11, -10, 1, 2,
    -- layer=1 filter=94 channel=87
    1, -7, 3, -6, 1, 5, 5, 4, 3,
    -- layer=1 filter=94 channel=88
    9, -8, -3, -9, -2, 6, 1, -1, -4,
    -- layer=1 filter=94 channel=89
    -4, -1, -9, 8, 0, 8, -9, 0, 7,
    -- layer=1 filter=94 channel=90
    -1, -5, -2, -2, -6, -6, 0, -5, 6,
    -- layer=1 filter=94 channel=91
    1, -1, -9, -4, -9, -2, 9, -9, 0,
    -- layer=1 filter=94 channel=92
    -2, 2, -5, 3, -9, -11, 4, 1, -6,
    -- layer=1 filter=94 channel=93
    -6, -4, 6, -5, 0, -6, 4, 9, 0,
    -- layer=1 filter=94 channel=94
    3, -2, -4, -10, -7, 6, 6, -6, 0,
    -- layer=1 filter=94 channel=95
    4, -12, 8, 0, -2, 3, -9, -1, 1,
    -- layer=1 filter=94 channel=96
    4, -3, -4, -5, 6, 4, 6, 6, -6,
    -- layer=1 filter=94 channel=97
    -9, -7, -6, 0, 1, 0, -8, -11, 5,
    -- layer=1 filter=94 channel=98
    8, -7, 2, 5, 4, -2, -3, -7, -5,
    -- layer=1 filter=94 channel=99
    5, -5, -1, 2, 3, -9, 4, -7, -9,
    -- layer=1 filter=94 channel=100
    -11, 1, 1, -4, -13, -11, -2, -7, 3,
    -- layer=1 filter=94 channel=101
    -6, -3, -8, 3, -7, -3, 3, 1, -3,
    -- layer=1 filter=94 channel=102
    5, 0, -7, -3, 8, 10, 0, -8, -4,
    -- layer=1 filter=94 channel=103
    -13, 3, -3, -15, -5, -5, -1, 1, -13,
    -- layer=1 filter=94 channel=104
    5, -4, -9, 7, 7, 10, -9, 1, -8,
    -- layer=1 filter=94 channel=105
    -6, -13, -13, -9, -5, -3, -2, -1, 0,
    -- layer=1 filter=94 channel=106
    6, 3, 2, -4, -5, 5, -8, -7, -10,
    -- layer=1 filter=94 channel=107
    0, 3, -5, 3, 9, 5, -4, 8, 2,
    -- layer=1 filter=94 channel=108
    -8, -1, 6, 3, 0, -6, -10, 9, 7,
    -- layer=1 filter=94 channel=109
    4, -6, -8, -4, 7, 6, -4, -2, -6,
    -- layer=1 filter=94 channel=110
    2, -8, 2, 7, -7, 1, -5, 0, -5,
    -- layer=1 filter=94 channel=111
    -9, -6, 9, 2, 6, -2, 6, -3, 9,
    -- layer=1 filter=94 channel=112
    -4, -2, -9, -4, -1, 7, -1, -5, -9,
    -- layer=1 filter=94 channel=113
    -2, -7, 0, 6, -5, -10, -14, 0, -12,
    -- layer=1 filter=94 channel=114
    -4, -6, 4, -6, 0, -7, 2, 6, 2,
    -- layer=1 filter=94 channel=115
    -8, 0, -13, 1, -15, -12, -11, 6, -1,
    -- layer=1 filter=94 channel=116
    4, 9, -7, 10, 4, -8, -5, 8, -4,
    -- layer=1 filter=94 channel=117
    5, 4, -3, -4, -4, 4, -2, 5, -5,
    -- layer=1 filter=94 channel=118
    -4, 6, 1, -7, -2, -2, 8, -5, 5,
    -- layer=1 filter=94 channel=119
    -7, -3, -3, -1, 4, -9, 5, -9, 0,
    -- layer=1 filter=94 channel=120
    -2, -7, -8, -2, 8, 7, -9, 0, 0,
    -- layer=1 filter=94 channel=121
    2, -14, -9, 1, -11, -10, -12, -8, -6,
    -- layer=1 filter=94 channel=122
    7, 4, -8, 7, -9, 0, 7, 8, 0,
    -- layer=1 filter=94 channel=123
    -3, 0, -7, 1, -6, -2, -12, -11, -12,
    -- layer=1 filter=94 channel=124
    -6, 3, 7, 7, -4, 1, 1, 2, 9,
    -- layer=1 filter=94 channel=125
    3, 9, -4, 6, 5, -8, -3, 5, 0,
    -- layer=1 filter=94 channel=126
    -9, -1, 10, 1, -2, 6, 2, 4, 9,
    -- layer=1 filter=94 channel=127
    2, -2, -11, 4, -7, -9, 10, -2, -8,
    -- layer=1 filter=95 channel=0
    5, -3, -10, -2, 5, 7, -12, 5, -3,
    -- layer=1 filter=95 channel=1
    -8, 0, -8, -12, 0, -7, -11, -9, -8,
    -- layer=1 filter=95 channel=2
    -4, -1, -8, -7, 0, -5, 1, -2, 9,
    -- layer=1 filter=95 channel=3
    4, -7, 8, -2, 6, 6, 1, -4, 1,
    -- layer=1 filter=95 channel=4
    -7, 3, 8, 7, -1, -6, 1, 3, -3,
    -- layer=1 filter=95 channel=5
    -3, 7, -9, 9, 7, 8, -5, -7, 2,
    -- layer=1 filter=95 channel=6
    1, -8, -7, 0, 8, 7, 2, -2, 7,
    -- layer=1 filter=95 channel=7
    10, 6, 5, 1, -2, -12, -3, 8, -5,
    -- layer=1 filter=95 channel=8
    -7, 6, -1, -2, -2, -7, 0, 0, -5,
    -- layer=1 filter=95 channel=9
    -1, -9, 0, -9, 2, -5, 2, -7, -7,
    -- layer=1 filter=95 channel=10
    -10, -3, 0, 8, -14, 6, -10, 0, -13,
    -- layer=1 filter=95 channel=11
    0, -4, -6, -2, -2, -3, -8, -5, -10,
    -- layer=1 filter=95 channel=12
    -8, -3, -5, 0, -4, 0, 5, -3, 6,
    -- layer=1 filter=95 channel=13
    8, 7, 5, -10, -9, -9, 1, -10, -2,
    -- layer=1 filter=95 channel=14
    1, 2, -7, 4, 8, 0, -11, 3, 8,
    -- layer=1 filter=95 channel=15
    1, 4, -5, 6, -8, 0, -6, -4, -11,
    -- layer=1 filter=95 channel=16
    -5, 0, -8, 1, 1, 4, -6, -8, -10,
    -- layer=1 filter=95 channel=17
    -11, 2, -7, -3, 0, 5, 0, -5, -4,
    -- layer=1 filter=95 channel=18
    11, 7, 1, 1, 0, 0, -1, -1, 6,
    -- layer=1 filter=95 channel=19
    -10, 0, -5, -11, -6, 2, -1, -9, -4,
    -- layer=1 filter=95 channel=20
    -8, -11, -11, -6, -4, 5, 3, -11, 7,
    -- layer=1 filter=95 channel=21
    -5, -4, 0, 8, -5, -5, 6, -10, -3,
    -- layer=1 filter=95 channel=22
    10, 9, -3, 5, 6, -8, -2, -1, 5,
    -- layer=1 filter=95 channel=23
    -6, 8, 2, -11, -5, -6, -5, -9, 5,
    -- layer=1 filter=95 channel=24
    6, 3, -5, -1, 0, 3, -6, 4, 0,
    -- layer=1 filter=95 channel=25
    -12, -4, 5, 5, 1, 4, 1, 6, -12,
    -- layer=1 filter=95 channel=26
    -10, -2, -6, -7, -2, 6, -8, 1, 7,
    -- layer=1 filter=95 channel=27
    -8, -6, -5, 9, 6, -7, 9, -5, 5,
    -- layer=1 filter=95 channel=28
    3, 4, 6, -10, -5, -8, -9, -7, 5,
    -- layer=1 filter=95 channel=29
    9, -8, 2, 6, 3, -6, 4, 7, -6,
    -- layer=1 filter=95 channel=30
    -4, -4, 0, -7, 6, -6, -2, -1, -11,
    -- layer=1 filter=95 channel=31
    0, -3, 0, 4, 7, -11, 7, 8, -1,
    -- layer=1 filter=95 channel=32
    7, 3, 8, -8, -10, -2, 0, -1, 6,
    -- layer=1 filter=95 channel=33
    2, 2, -1, -4, 5, -10, -6, -8, 2,
    -- layer=1 filter=95 channel=34
    -9, 8, 8, -9, 1, 4, 7, -3, -3,
    -- layer=1 filter=95 channel=35
    -1, -8, -6, 5, 5, 0, 7, -6, 0,
    -- layer=1 filter=95 channel=36
    4, 4, -6, -3, 7, -7, -5, -11, -3,
    -- layer=1 filter=95 channel=37
    -12, 4, -2, -4, 0, 8, -2, 9, 0,
    -- layer=1 filter=95 channel=38
    5, -5, -3, -1, 5, -7, -8, -6, -4,
    -- layer=1 filter=95 channel=39
    -11, -4, 1, -1, 6, 0, -5, -9, -3,
    -- layer=1 filter=95 channel=40
    3, -10, 8, -6, 8, 3, 0, -4, -4,
    -- layer=1 filter=95 channel=41
    0, 4, 6, -10, 0, -8, 6, -5, -4,
    -- layer=1 filter=95 channel=42
    -1, 5, 4, 9, -5, 7, -7, -5, 6,
    -- layer=1 filter=95 channel=43
    -6, -2, 3, -4, -5, 8, -10, -9, 9,
    -- layer=1 filter=95 channel=44
    -4, 3, 1, -10, 3, 4, -2, -1, 2,
    -- layer=1 filter=95 channel=45
    7, 0, 7, -11, 4, -1, -3, -2, -7,
    -- layer=1 filter=95 channel=46
    -7, 2, 4, 3, 9, -8, 7, 0, 6,
    -- layer=1 filter=95 channel=47
    0, -6, -10, 3, 0, 6, 4, 2, 4,
    -- layer=1 filter=95 channel=48
    -7, 6, -1, -5, -2, -2, -8, 3, -11,
    -- layer=1 filter=95 channel=49
    11, 8, 5, -5, 5, 1, -3, 4, -5,
    -- layer=1 filter=95 channel=50
    5, 5, 1, 8, 1, 6, -11, 8, 6,
    -- layer=1 filter=95 channel=51
    2, 0, -7, 4, 4, 8, 5, -10, -5,
    -- layer=1 filter=95 channel=52
    -7, 2, 0, 2, 3, -3, 1, 8, -7,
    -- layer=1 filter=95 channel=53
    6, -3, -4, -1, 1, -9, -2, 2, 4,
    -- layer=1 filter=95 channel=54
    -1, -5, -10, -5, -9, -11, 5, -7, -2,
    -- layer=1 filter=95 channel=55
    0, -7, 0, 8, 7, -6, 4, 5, 9,
    -- layer=1 filter=95 channel=56
    2, 2, 9, 5, -4, 8, -10, 3, 5,
    -- layer=1 filter=95 channel=57
    6, 3, -1, -5, 7, 1, 3, 2, 4,
    -- layer=1 filter=95 channel=58
    -1, 5, -7, 4, 1, -7, 10, -9, -10,
    -- layer=1 filter=95 channel=59
    -5, 3, -10, -10, -6, 1, -7, 3, -7,
    -- layer=1 filter=95 channel=60
    -10, -4, -6, -7, 0, -3, 5, -7, 12,
    -- layer=1 filter=95 channel=61
    1, 2, 0, -9, 1, 3, -6, -8, 3,
    -- layer=1 filter=95 channel=62
    0, -8, 7, -7, -1, 4, 3, 1, -10,
    -- layer=1 filter=95 channel=63
    -3, -2, -1, -5, -11, 2, -2, 8, -10,
    -- layer=1 filter=95 channel=64
    8, -3, -6, 5, -8, 5, -4, -3, 5,
    -- layer=1 filter=95 channel=65
    -2, -11, 1, 8, 6, -2, 1, 7, 3,
    -- layer=1 filter=95 channel=66
    -10, -9, -12, 6, 8, -3, -11, 8, 0,
    -- layer=1 filter=95 channel=67
    -3, 3, -2, 1, 8, 3, 2, 2, -6,
    -- layer=1 filter=95 channel=68
    3, -6, 8, 0, -8, -1, -6, -2, -2,
    -- layer=1 filter=95 channel=69
    6, -9, -8, 5, 10, 4, -2, 5, 5,
    -- layer=1 filter=95 channel=70
    -3, -3, -5, -8, -10, -8, 5, 4, 8,
    -- layer=1 filter=95 channel=71
    4, 3, 5, 4, -3, 2, -5, -9, -9,
    -- layer=1 filter=95 channel=72
    7, 7, -2, 7, 6, 7, -1, 0, 7,
    -- layer=1 filter=95 channel=73
    -9, 3, -7, -3, -4, -10, -6, -10, -5,
    -- layer=1 filter=95 channel=74
    -11, -7, -7, -11, -4, -4, 2, 5, -3,
    -- layer=1 filter=95 channel=75
    -8, 7, -8, -9, 1, 3, -2, 9, -6,
    -- layer=1 filter=95 channel=76
    0, -1, -11, 4, -5, 0, -10, 7, -11,
    -- layer=1 filter=95 channel=77
    -10, -7, -7, -1, 2, 3, -9, 5, 6,
    -- layer=1 filter=95 channel=78
    0, 8, 6, 4, -8, -6, 7, -5, 0,
    -- layer=1 filter=95 channel=79
    9, 5, -3, -3, -11, 2, 4, 5, -10,
    -- layer=1 filter=95 channel=80
    3, -2, 6, 10, -8, 0, 0, -5, -9,
    -- layer=1 filter=95 channel=81
    -2, -4, 0, 3, 4, 2, -2, -8, -1,
    -- layer=1 filter=95 channel=82
    5, -9, -11, -9, -7, 3, 7, 6, 6,
    -- layer=1 filter=95 channel=83
    -11, 5, -7, 1, 0, -5, -1, -10, 8,
    -- layer=1 filter=95 channel=84
    7, -7, 1, -10, -10, 3, -6, -6, -2,
    -- layer=1 filter=95 channel=85
    -10, 7, 0, -1, -2, 4, 2, -8, -1,
    -- layer=1 filter=95 channel=86
    5, 5, 0, -13, -9, -10, -11, -6, -10,
    -- layer=1 filter=95 channel=87
    -5, -8, -9, -10, 3, 6, -6, -6, -11,
    -- layer=1 filter=95 channel=88
    4, 3, 9, 1, 0, -3, -2, 7, -11,
    -- layer=1 filter=95 channel=89
    1, 4, 8, -9, -8, -1, -5, -3, -1,
    -- layer=1 filter=95 channel=90
    -10, -6, -11, -4, -8, -9, -10, 0, -3,
    -- layer=1 filter=95 channel=91
    -11, -9, 4, 6, -6, 4, 0, -12, -5,
    -- layer=1 filter=95 channel=92
    3, -2, 2, 0, -6, -6, 7, 0, 3,
    -- layer=1 filter=95 channel=93
    -8, -1, -2, 4, -3, 6, 8, 0, 3,
    -- layer=1 filter=95 channel=94
    -5, -3, 0, -4, -2, -8, 1, 8, -1,
    -- layer=1 filter=95 channel=95
    12, -1, 2, -1, -6, 6, 5, -10, -9,
    -- layer=1 filter=95 channel=96
    -11, -5, 7, -10, -2, 4, -5, 1, 0,
    -- layer=1 filter=95 channel=97
    0, 5, 2, -11, 0, -3, 0, 5, -10,
    -- layer=1 filter=95 channel=98
    0, 0, 8, -12, 2, -13, 6, -9, -3,
    -- layer=1 filter=95 channel=99
    -5, 4, 1, 1, 9, -6, 0, -10, -1,
    -- layer=1 filter=95 channel=100
    -1, -8, 2, -3, -4, -3, -2, 1, 2,
    -- layer=1 filter=95 channel=101
    -5, 7, -9, -6, -5, 8, -7, 8, 8,
    -- layer=1 filter=95 channel=102
    6, 3, 8, -8, 4, 4, -5, -5, -1,
    -- layer=1 filter=95 channel=103
    -6, -4, 0, -12, -8, -1, -4, -5, 6,
    -- layer=1 filter=95 channel=104
    -8, 0, 3, 1, -2, -3, -4, 8, 0,
    -- layer=1 filter=95 channel=105
    -2, -2, 1, 1, -2, 3, 2, -8, -5,
    -- layer=1 filter=95 channel=106
    -7, -8, -8, 4, 7, 6, -6, -3, 3,
    -- layer=1 filter=95 channel=107
    11, 4, 10, -3, 4, 9, -5, -6, 0,
    -- layer=1 filter=95 channel=108
    3, -1, 0, 9, 0, -5, -7, -2, -9,
    -- layer=1 filter=95 channel=109
    1, 1, 3, -6, 4, 9, 5, 3, -2,
    -- layer=1 filter=95 channel=110
    -9, -1, 4, 6, 3, 4, 0, 8, 0,
    -- layer=1 filter=95 channel=111
    6, 1, -9, -2, -9, -6, -9, -7, -1,
    -- layer=1 filter=95 channel=112
    0, 5, -5, -1, -4, 2, -2, -6, 1,
    -- layer=1 filter=95 channel=113
    9, 1, -6, 0, -2, -5, 0, 4, 9,
    -- layer=1 filter=95 channel=114
    -8, 3, -1, -9, 3, 9, -7, -3, 8,
    -- layer=1 filter=95 channel=115
    -3, -2, -6, -5, -1, 5, -7, -4, -9,
    -- layer=1 filter=95 channel=116
    -7, 0, -4, -7, -1, 8, 8, -10, 0,
    -- layer=1 filter=95 channel=117
    2, 0, 4, 10, -2, -7, 4, 5, 2,
    -- layer=1 filter=95 channel=118
    -8, 7, -7, -9, 0, 5, 4, -12, 3,
    -- layer=1 filter=95 channel=119
    1, 0, 8, 1, 8, 0, 1, 8, -9,
    -- layer=1 filter=95 channel=120
    -4, -3, -4, -6, 1, 1, 6, 7, -5,
    -- layer=1 filter=95 channel=121
    -1, -11, -6, 2, -4, -6, 3, 1, 8,
    -- layer=1 filter=95 channel=122
    6, 8, -4, 3, 10, -6, 4, -4, 0,
    -- layer=1 filter=95 channel=123
    8, -7, 4, -10, 7, 1, 6, 5, -10,
    -- layer=1 filter=95 channel=124
    8, 1, -5, -9, 0, -4, -8, -8, -3,
    -- layer=1 filter=95 channel=125
    6, 0, -7, 3, -1, 9, 0, 2, 4,
    -- layer=1 filter=95 channel=126
    -4, 5, 0, -7, 3, -6, -6, -9, 1,
    -- layer=1 filter=95 channel=127
    -7, 3, -4, 1, -11, -5, 2, 6, 0,
    -- layer=1 filter=96 channel=0
    15, -6, -7, 0, 0, -3, -7, 0, -6,
    -- layer=1 filter=96 channel=1
    23, 19, -2, -2, 30, 27, -34, -29, -21,
    -- layer=1 filter=96 channel=2
    12, 24, 3, -16, -43, -39, 3, -68, -35,
    -- layer=1 filter=96 channel=3
    9, -16, -1, 5, 2, -5, 10, -1, -5,
    -- layer=1 filter=96 channel=4
    -3, -2, 0, -1, -9, -2, 10, -4, 7,
    -- layer=1 filter=96 channel=5
    9, 26, -17, 19, 38, 36, -60, -39, 5,
    -- layer=1 filter=96 channel=6
    55, 43, 24, 19, 9, -21, -23, -30, -35,
    -- layer=1 filter=96 channel=7
    -6, -36, -30, 5, -9, -38, 17, -20, -12,
    -- layer=1 filter=96 channel=8
    4, 0, -19, 8, 23, 9, -25, -40, -1,
    -- layer=1 filter=96 channel=9
    0, -13, 6, 34, -39, -3, -39, -19, -15,
    -- layer=1 filter=96 channel=10
    2, -42, -29, 2, 26, -30, 29, -2, 0,
    -- layer=1 filter=96 channel=11
    6, -3, -1, 17, -10, 5, 25, 38, 27,
    -- layer=1 filter=96 channel=12
    -87, -45, 0, 34, -41, -44, -51, -72, -50,
    -- layer=1 filter=96 channel=13
    56, 53, 32, 1, 8, 3, -24, -39, -44,
    -- layer=1 filter=96 channel=14
    -23, -37, -14, -12, 0, -48, 6, -7, -3,
    -- layer=1 filter=96 channel=15
    10, 34, 1, -60, -35, 6, -27, -39, -5,
    -- layer=1 filter=96 channel=16
    20, -17, -44, 7, 12, -8, -41, -55, -6,
    -- layer=1 filter=96 channel=17
    28, 15, -5, 8, 12, 6, -18, -8, -12,
    -- layer=1 filter=96 channel=18
    12, 3, 25, 26, 7, -12, 36, 32, 18,
    -- layer=1 filter=96 channel=19
    17, 14, -15, 26, 7, -37, 9, 25, 50,
    -- layer=1 filter=96 channel=20
    60, 63, 25, 5, 13, -10, -30, -35, -57,
    -- layer=1 filter=96 channel=21
    28, 33, 39, 0, 0, -7, -47, -48, -59,
    -- layer=1 filter=96 channel=22
    36, 58, 39, 5, -3, 0, -46, -41, -69,
    -- layer=1 filter=96 channel=23
    -47, -24, -53, -57, -56, -41, 11, -14, -27,
    -- layer=1 filter=96 channel=24
    5, -10, -5, -22, -13, -5, -43, -28, -19,
    -- layer=1 filter=96 channel=25
    8, -15, -47, 21, -14, -28, 16, -49, -37,
    -- layer=1 filter=96 channel=26
    14, 10, 20, 2, 10, -5, -11, -13, -19,
    -- layer=1 filter=96 channel=27
    -12, -7, 11, 1, 7, 15, 19, 18, 23,
    -- layer=1 filter=96 channel=28
    -14, -14, -25, -4, -10, -39, -8, -12, -23,
    -- layer=1 filter=96 channel=29
    8, -4, 21, 19, 25, 29, 6, -3, -3,
    -- layer=1 filter=96 channel=30
    15, 5, 9, 38, 38, -12, 43, 14, 21,
    -- layer=1 filter=96 channel=31
    -14, 14, 31, 27, 30, -4, 4, -7, 6,
    -- layer=1 filter=96 channel=32
    3, 13, 19, 45, 7, -4, 39, 8, 8,
    -- layer=1 filter=96 channel=33
    24, 6, -3, 2, 5, 3, 10, -4, -3,
    -- layer=1 filter=96 channel=34
    29, 29, -3, 15, -5, 0, 17, -4, -5,
    -- layer=1 filter=96 channel=35
    -5, 5, 4, -3, -5, 8, 6, -3, 8,
    -- layer=1 filter=96 channel=36
    -2, -12, -1, 10, -4, -3, 21, 39, 21,
    -- layer=1 filter=96 channel=37
    24, 5, -18, 18, 54, 35, -56, -30, 15,
    -- layer=1 filter=96 channel=38
    43, 64, 30, 9, 7, -2, -35, -41, -47,
    -- layer=1 filter=96 channel=39
    -5, -7, 0, 10, 2, 4, -9, 17, 16,
    -- layer=1 filter=96 channel=40
    39, 46, 31, 7, 6, -27, -2, -5, -33,
    -- layer=1 filter=96 channel=41
    -5, -14, 7, 72, -27, -10, 61, 5, 9,
    -- layer=1 filter=96 channel=42
    26, 3, -5, -34, -60, -44, -7, -56, -74,
    -- layer=1 filter=96 channel=43
    13, -17, -34, 4, 2, -19, -21, -26, -15,
    -- layer=1 filter=96 channel=44
    17, 22, 16, 20, 22, 7, 6, 5, -13,
    -- layer=1 filter=96 channel=45
    34, 14, 15, -2, 16, 0, -43, -42, -28,
    -- layer=1 filter=96 channel=46
    9, 6, -26, 5, 18, -33, -53, -25, 32,
    -- layer=1 filter=96 channel=47
    -59, -7, 10, 15, -26, 26, 39, -16, -13,
    -- layer=1 filter=96 channel=48
    34, 39, 20, 7, -9, 8, -15, -43, -46,
    -- layer=1 filter=96 channel=49
    10, 19, 0, 25, 0, -7, -16, -37, -40,
    -- layer=1 filter=96 channel=50
    0, 4, 10, -1, -8, -12, -2, -22, -25,
    -- layer=1 filter=96 channel=51
    21, 26, 13, -1, 4, -9, -16, -51, -44,
    -- layer=1 filter=96 channel=52
    -10, -23, -8, -14, -21, -17, 4, 2, 17,
    -- layer=1 filter=96 channel=53
    14, 7, 22, 18, 7, 5, 3, 7, 2,
    -- layer=1 filter=96 channel=54
    33, -19, -63, 22, 15, -23, 17, -44, -13,
    -- layer=1 filter=96 channel=55
    -27, -46, -28, 1, 10, 19, 30, 19, 36,
    -- layer=1 filter=96 channel=56
    -7, -9, 3, 4, 5, -1, 10, -1, 3,
    -- layer=1 filter=96 channel=57
    21, 0, -1, 5, 27, -3, 20, -16, 0,
    -- layer=1 filter=96 channel=58
    -46, -23, -61, -6, -45, -56, 58, -49, 5,
    -- layer=1 filter=96 channel=59
    -1, 1, -5, 3, -9, -8, 8, 10, 7,
    -- layer=1 filter=96 channel=60
    -12, -16, -12, -11, -7, -3, -5, -17, 10,
    -- layer=1 filter=96 channel=61
    6, 4, -9, 12, 8, 6, -1, 2, 3,
    -- layer=1 filter=96 channel=62
    22, 0, -35, -2, 38, 5, -47, -52, -7,
    -- layer=1 filter=96 channel=63
    1, -4, 8, 22, -8, -7, 33, 29, 11,
    -- layer=1 filter=96 channel=64
    26, 41, 11, 4, 1, 15, -15, -14, -21,
    -- layer=1 filter=96 channel=65
    31, 30, 34, -4, -4, -13, -31, -58, -44,
    -- layer=1 filter=96 channel=66
    3, -7, -15, 11, 0, 9, 3, 8, 2,
    -- layer=1 filter=96 channel=67
    12, 24, -1, 14, 16, 20, -12, -30, -31,
    -- layer=1 filter=96 channel=68
    13, -1, 18, 36, 20, 4, -4, 5, -16,
    -- layer=1 filter=96 channel=69
    1, -10, -28, -46, 2, -1, -73, -28, -5,
    -- layer=1 filter=96 channel=70
    -7, 4, -13, 5, 18, 20, -15, -38, -24,
    -- layer=1 filter=96 channel=71
    11, -9, -11, -15, -14, -12, -30, -32, 0,
    -- layer=1 filter=96 channel=72
    -12, 14, 20, 34, -17, -40, 14, 5, 54,
    -- layer=1 filter=96 channel=73
    -5, -2, -16, 5, -5, -4, -10, -17, -11,
    -- layer=1 filter=96 channel=74
    30, 3, 20, 42, 14, -19, -30, -7, -34,
    -- layer=1 filter=96 channel=75
    -13, -9, 18, 0, -42, -51, -23, -28, 15,
    -- layer=1 filter=96 channel=76
    19, 6, 16, 21, 1, -11, 14, -6, -21,
    -- layer=1 filter=96 channel=77
    21, 25, 35, -11, -4, 5, -20, -32, -40,
    -- layer=1 filter=96 channel=78
    -3, 0, -3, -1, 4, -19, -7, -5, -2,
    -- layer=1 filter=96 channel=79
    25, 16, -13, -21, 0, -11, -41, -50, 0,
    -- layer=1 filter=96 channel=80
    1, -1, 4, 5, -6, -6, -3, 4, -6,
    -- layer=1 filter=96 channel=81
    -11, -4, -17, -16, -42, -18, -17, -26, -14,
    -- layer=1 filter=96 channel=82
    39, 33, 45, 7, 6, 0, -30, -45, -61,
    -- layer=1 filter=96 channel=83
    6, -6, 0, -3, 22, 10, -42, -32, -22,
    -- layer=1 filter=96 channel=84
    39, 12, 39, 51, 0, -1, 28, 10, -25,
    -- layer=1 filter=96 channel=85
    -36, -22, -14, 22, -22, -34, 32, 2, -1,
    -- layer=1 filter=96 channel=86
    -3, -2, -21, 16, 14, 2, 15, 22, 17,
    -- layer=1 filter=96 channel=87
    -25, 18, -12, 30, 0, -5, -7, 10, 28,
    -- layer=1 filter=96 channel=88
    20, 26, 18, -3, 11, 0, -19, -32, -39,
    -- layer=1 filter=96 channel=89
    23, 29, 40, -7, -21, -11, -45, -42, -71,
    -- layer=1 filter=96 channel=90
    6, -5, 14, -1, 18, 6, -27, -14, -16,
    -- layer=1 filter=96 channel=91
    42, 60, 43, 17, 18, 3, -2, -26, -51,
    -- layer=1 filter=96 channel=92
    13, -15, -9, -21, -16, -16, -12, -8, -5,
    -- layer=1 filter=96 channel=93
    19, 1, -6, 0, -2, -9, -41, -39, -25,
    -- layer=1 filter=96 channel=94
    3, 3, -2, 19, -8, -4, 3, 2, 0,
    -- layer=1 filter=96 channel=95
    42, 31, 39, 69, 26, -8, 12, 17, 0,
    -- layer=1 filter=96 channel=96
    1, 13, 13, 16, 8, 0, 2, 7, -6,
    -- layer=1 filter=96 channel=97
    11, 7, -7, 4, 1, 3, -21, -14, -6,
    -- layer=1 filter=96 channel=98
    18, -1, -20, -2, -7, -4, -54, -54, -36,
    -- layer=1 filter=96 channel=99
    -2, -53, -16, -32, -2, -47, -35, -18, -23,
    -- layer=1 filter=96 channel=100
    -2, 2, 6, 14, 12, 10, 26, 35, 23,
    -- layer=1 filter=96 channel=101
    47, 46, 35, 23, 9, -5, -39, -41, -65,
    -- layer=1 filter=96 channel=102
    34, 30, 11, 23, 5, 4, -23, -16, -7,
    -- layer=1 filter=96 channel=103
    -6, 5, 12, 19, 8, 6, 33, 16, 23,
    -- layer=1 filter=96 channel=104
    -56, -23, -27, -9, -28, -29, 26, -27, -6,
    -- layer=1 filter=96 channel=105
    1, 0, -10, 0, -8, -1, -10, 8, -2,
    -- layer=1 filter=96 channel=106
    48, 47, 29, 35, 17, 0, -23, -38, -61,
    -- layer=1 filter=96 channel=107
    3, 13, -4, -3, -3, 6, -9, -7, -4,
    -- layer=1 filter=96 channel=108
    11, -14, -21, 8, 4, -20, -3, 1, -19,
    -- layer=1 filter=96 channel=109
    9, 5, 6, 10, 3, -3, -3, 1, 6,
    -- layer=1 filter=96 channel=110
    0, -2, 1, 1, 0, 4, -1, 0, -8,
    -- layer=1 filter=96 channel=111
    32, 6, 22, 36, 21, -17, 4, -3, -17,
    -- layer=1 filter=96 channel=112
    31, 0, 10, 18, -7, 4, -12, -9, -27,
    -- layer=1 filter=96 channel=113
    49, 39, 10, 10, -3, -29, -14, -43, -63,
    -- layer=1 filter=96 channel=114
    -31, -24, -36, -5, 13, 26, -29, -35, -8,
    -- layer=1 filter=96 channel=115
    3, -28, -15, -2, -9, -16, 13, -5, 14,
    -- layer=1 filter=96 channel=116
    2, -8, -6, -3, 2, 1, 8, 5, -1,
    -- layer=1 filter=96 channel=117
    18, -15, 23, -7, -11, 25, -32, -14, -51,
    -- layer=1 filter=96 channel=118
    22, 1, 31, 43, 22, -10, 7, 2, -15,
    -- layer=1 filter=96 channel=119
    3, -1, 8, 38, 31, -2, 23, 4, 7,
    -- layer=1 filter=96 channel=120
    8, 29, 16, -8, 2, -2, -11, -52, -56,
    -- layer=1 filter=96 channel=121
    -15, -24, -11, 0, 4, -4, -3, 10, 36,
    -- layer=1 filter=96 channel=122
    -1, -8, 4, -9, 5, -10, -9, 0, -6,
    -- layer=1 filter=96 channel=123
    -21, -35, -5, 1, 7, -7, 22, 7, 37,
    -- layer=1 filter=96 channel=124
    -3, -13, 1, -3, -17, -2, -10, -13, -13,
    -- layer=1 filter=96 channel=125
    25, 32, 0, 23, 40, 15, -12, -42, -70,
    -- layer=1 filter=96 channel=126
    -13, -5, 25, -9, 30, 51, -56, -52, -2,
    -- layer=1 filter=96 channel=127
    12, 7, 33, 43, 40, 8, 22, 38, 23,
    -- layer=1 filter=97 channel=0
    -9, -12, -1, 6, -6, -15, -8, 10, -10,
    -- layer=1 filter=97 channel=1
    -18, -33, -23, -35, -30, -21, 5, -19, -14,
    -- layer=1 filter=97 channel=2
    33, 29, 32, 31, 34, 29, 52, 54, 65,
    -- layer=1 filter=97 channel=3
    -8, 7, 13, 6, 6, -6, 7, 2, 12,
    -- layer=1 filter=97 channel=4
    9, 0, 8, -5, 8, 6, -8, -3, 5,
    -- layer=1 filter=97 channel=5
    -72, -103, -68, -92, -87, -75, -40, -24, -55,
    -- layer=1 filter=97 channel=6
    39, 16, 0, 5, 13, -2, 20, 0, -1,
    -- layer=1 filter=97 channel=7
    -38, -51, -47, -49, -60, -71, -41, 20, -53,
    -- layer=1 filter=97 channel=8
    -42, -80, -43, -146, -142, -102, -67, -70, -52,
    -- layer=1 filter=97 channel=9
    -6, 10, -18, 4, 21, -15, 40, 26, 41,
    -- layer=1 filter=97 channel=10
    -38, -46, -42, -39, -32, -34, -30, 24, -24,
    -- layer=1 filter=97 channel=11
    -3, 11, 7, 12, 9, 18, 12, 11, 5,
    -- layer=1 filter=97 channel=12
    7, -7, -3, 15, 17, 32, 61, 60, 58,
    -- layer=1 filter=97 channel=13
    21, 21, 16, 13, 9, 20, 3, -9, 10,
    -- layer=1 filter=97 channel=14
    -54, -10, 3, 11, -15, -10, 2, 73, -20,
    -- layer=1 filter=97 channel=15
    -22, -33, 25, -27, -24, -18, 6, 0, -42,
    -- layer=1 filter=97 channel=16
    -51, -102, -44, -133, -125, -92, -29, -73, -78,
    -- layer=1 filter=97 channel=17
    18, 11, 10, -5, -1, 6, 13, 0, -11,
    -- layer=1 filter=97 channel=18
    -19, -23, -12, 14, -1, -15, 12, 41, 27,
    -- layer=1 filter=97 channel=19
    -69, -64, -72, -104, -127, -104, -48, -94, -71,
    -- layer=1 filter=97 channel=20
    41, 21, 29, 9, 4, 12, 12, 9, -5,
    -- layer=1 filter=97 channel=21
    -9, -9, -11, -8, -3, -1, -7, -1, -9,
    -- layer=1 filter=97 channel=22
    36, 37, 23, 10, 3, 4, 20, 4, 1,
    -- layer=1 filter=97 channel=23
    -11, -32, -8, -3, -24, -17, 25, -4, -34,
    -- layer=1 filter=97 channel=24
    -26, 2, 10, -8, -15, 8, -6, -10, 33,
    -- layer=1 filter=97 channel=25
    -19, -58, -64, -58, -68, -83, -43, -39, -59,
    -- layer=1 filter=97 channel=26
    7, 22, 41, 3, 5, 44, 22, 8, 29,
    -- layer=1 filter=97 channel=27
    -28, -11, -19, -2, 4, 6, 8, 21, -4,
    -- layer=1 filter=97 channel=28
    -34, -18, -25, -23, -30, -22, -33, 7, -8,
    -- layer=1 filter=97 channel=29
    -25, -3, 0, -7, -3, -4, -13, -6, -3,
    -- layer=1 filter=97 channel=30
    -73, -116, -76, -46, -72, -84, -21, 10, -7,
    -- layer=1 filter=97 channel=31
    6, -22, -32, -7, 12, 8, 49, 62, 50,
    -- layer=1 filter=97 channel=32
    -27, -29, 18, -12, -44, 21, 18, -10, 44,
    -- layer=1 filter=97 channel=33
    16, 12, 8, 0, -7, 11, 10, 5, 8,
    -- layer=1 filter=97 channel=34
    2, -3, -11, 10, -7, -8, -4, 14, -1,
    -- layer=1 filter=97 channel=35
    -11, -2, -10, -13, -12, -7, -9, -14, 2,
    -- layer=1 filter=97 channel=36
    5, 14, 17, 16, 24, 16, 12, 19, 6,
    -- layer=1 filter=97 channel=37
    -73, -74, -57, -77, -89, -83, -47, -74, -62,
    -- layer=1 filter=97 channel=38
    14, 9, 6, 9, 15, 1, 9, -6, 9,
    -- layer=1 filter=97 channel=39
    -3, -11, -15, -28, -3, -18, -6, -4, -7,
    -- layer=1 filter=97 channel=40
    6, -7, 0, 11, 4, -6, 45, 54, 19,
    -- layer=1 filter=97 channel=41
    5, -18, 13, -7, -25, -6, 18, 14, 48,
    -- layer=1 filter=97 channel=42
    25, 6, 29, 15, 38, 19, 57, 45, 27,
    -- layer=1 filter=97 channel=43
    -49, -71, -47, -118, -121, -106, -58, -55, -51,
    -- layer=1 filter=97 channel=44
    -19, -34, 41, -11, -42, 32, 13, -27, 53,
    -- layer=1 filter=97 channel=45
    -10, 0, 21, -17, 0, -1, 2, -23, -9,
    -- layer=1 filter=97 channel=46
    -93, -58, -28, -91, -101, -53, -31, -74, -48,
    -- layer=1 filter=97 channel=47
    22, -20, -26, 20, -6, -27, 41, 10, -21,
    -- layer=1 filter=97 channel=48
    7, -18, -8, 8, -5, 7, -17, 0, -4,
    -- layer=1 filter=97 channel=49
    -5, -3, -17, -6, -12, -10, 6, -2, -6,
    -- layer=1 filter=97 channel=50
    10, 12, 17, 5, 17, 16, 29, 20, 31,
    -- layer=1 filter=97 channel=51
    -7, -5, 7, -8, 8, 0, -7, 9, 2,
    -- layer=1 filter=97 channel=52
    9, 16, 12, 20, 16, -1, 17, 2, 4,
    -- layer=1 filter=97 channel=53
    -3, -11, -6, -17, -19, -8, -15, -17, -8,
    -- layer=1 filter=97 channel=54
    -49, -29, -58, -74, -38, -50, -30, -43, -29,
    -- layer=1 filter=97 channel=55
    10, 23, 23, 15, 35, 18, 24, 37, 12,
    -- layer=1 filter=97 channel=56
    3, -4, 7, -1, 0, -10, -10, -10, 2,
    -- layer=1 filter=97 channel=57
    7, 3, -12, -6, -13, 0, 4, 45, -2,
    -- layer=1 filter=97 channel=58
    -41, -97, -67, -27, -95, -57, 2, 36, -70,
    -- layer=1 filter=97 channel=59
    -6, -8, -1, 3, -3, -3, -9, -10, 7,
    -- layer=1 filter=97 channel=60
    8, 11, 13, 14, 20, 18, 15, 10, 15,
    -- layer=1 filter=97 channel=61
    0, -14, -9, -7, 3, -14, -2, -7, 0,
    -- layer=1 filter=97 channel=62
    -88, -104, -31, -128, -158, -113, -72, -112, -79,
    -- layer=1 filter=97 channel=63
    4, 15, 5, 4, 19, 10, 7, 10, 16,
    -- layer=1 filter=97 channel=64
    17, 11, 0, 5, -10, -8, -7, 1, -6,
    -- layer=1 filter=97 channel=65
    0, -12, 2, -5, 7, -12, -11, -18, -1,
    -- layer=1 filter=97 channel=66
    5, -7, 0, -3, -2, -6, 0, 2, -4,
    -- layer=1 filter=97 channel=67
    2, -35, -47, -24, -4, -20, -39, -27, -17,
    -- layer=1 filter=97 channel=68
    -50, -18, 37, -49, -53, 27, 4, -31, 57,
    -- layer=1 filter=97 channel=69
    -18, -34, 23, -28, -40, 19, -12, 12, -19,
    -- layer=1 filter=97 channel=70
    6, -11, -40, 5, -19, -16, 10, 22, -15,
    -- layer=1 filter=97 channel=71
    -10, -24, -16, -31, 0, 6, -5, -3, 14,
    -- layer=1 filter=97 channel=72
    -29, -37, -23, -75, -33, -41, -13, -22, 10,
    -- layer=1 filter=97 channel=73
    -6, -2, -5, -7, 7, -9, -5, 10, -2,
    -- layer=1 filter=97 channel=74
    -17, -42, 15, -14, -29, 32, 43, 19, 76,
    -- layer=1 filter=97 channel=75
    -33, -14, 21, -19, -23, -30, 53, 49, 28,
    -- layer=1 filter=97 channel=76
    -14, 2, 12, -9, -15, -2, 10, -7, 29,
    -- layer=1 filter=97 channel=77
    -2, -18, -13, -12, 1, -4, -18, 1, 6,
    -- layer=1 filter=97 channel=78
    2, 11, 2, 7, 12, -3, -5, 10, -4,
    -- layer=1 filter=97 channel=79
    -28, -66, -19, -94, -105, -77, -12, -46, -58,
    -- layer=1 filter=97 channel=80
    5, -2, -7, 0, 8, -5, 6, 7, 6,
    -- layer=1 filter=97 channel=81
    -16, -26, -17, -14, -17, -5, 6, -2, 17,
    -- layer=1 filter=97 channel=82
    -7, -23, -12, -2, -13, 7, -18, -1, -9,
    -- layer=1 filter=97 channel=83
    -19, -19, 8, -16, -24, 13, -9, -41, 9,
    -- layer=1 filter=97 channel=84
    -101, -104, -41, -24, -59, -29, 3, 4, 55,
    -- layer=1 filter=97 channel=85
    0, -1, -25, 6, -35, -27, 19, -14, -44,
    -- layer=1 filter=97 channel=86
    14, 20, 7, 11, 20, 11, 0, 8, -5,
    -- layer=1 filter=97 channel=87
    -43, -23, -65, -68, -42, -57, -3, -25, -11,
    -- layer=1 filter=97 channel=88
    -1, -23, -24, -3, -11, -8, -9, -9, 0,
    -- layer=1 filter=97 channel=89
    -17, -8, 0, -16, -21, -5, 9, -16, 7,
    -- layer=1 filter=97 channel=90
    -29, -8, 31, -24, -62, 35, 7, -29, 26,
    -- layer=1 filter=97 channel=91
    27, 27, 1, 15, 7, -1, 22, 6, 3,
    -- layer=1 filter=97 channel=92
    -13, 14, 20, 6, 9, 27, 7, 95, 19,
    -- layer=1 filter=97 channel=93
    -4, 11, 4, 6, 5, -2, 3, -2, 8,
    -- layer=1 filter=97 channel=94
    -9, 2, 0, 3, -4, -5, -12, 5, -3,
    -- layer=1 filter=97 channel=95
    -93, -118, -48, -38, -72, -47, -17, 0, 23,
    -- layer=1 filter=97 channel=96
    -3, 5, 6, 12, 4, 0, 5, 1, 17,
    -- layer=1 filter=97 channel=97
    11, -2, -8, 13, 9, 2, -4, -1, 6,
    -- layer=1 filter=97 channel=98
    -11, -9, -2, -56, -72, -36, -51, -37, -24,
    -- layer=1 filter=97 channel=99
    -69, -47, -37, -23, -6, -9, -32, 17, 14,
    -- layer=1 filter=97 channel=100
    3, 7, 18, -5, 19, 11, -8, 6, -4,
    -- layer=1 filter=97 channel=101
    28, 10, 2, 21, 7, 17, 13, 3, 20,
    -- layer=1 filter=97 channel=102
    9, -6, -4, 9, 3, -6, -13, 1, -13,
    -- layer=1 filter=97 channel=103
    -5, 5, 12, 6, 13, -7, 12, 13, 4,
    -- layer=1 filter=97 channel=104
    15, -3, -22, -3, -3, -16, 18, 14, -13,
    -- layer=1 filter=97 channel=105
    5, 1, 6, 1, 2, -8, -9, 0, 4,
    -- layer=1 filter=97 channel=106
    37, 25, 24, 32, 13, 31, 33, 0, 28,
    -- layer=1 filter=97 channel=107
    14, 11, -5, 3, 0, 15, -1, 0, 18,
    -- layer=1 filter=97 channel=108
    -67, -59, 11, -59, -82, 2, -9, -50, 7,
    -- layer=1 filter=97 channel=109
    4, 5, 9, 0, -6, -7, -8, -6, 3,
    -- layer=1 filter=97 channel=110
    -8, -4, 0, 9, 10, -4, -11, 2, -10,
    -- layer=1 filter=97 channel=111
    -65, -103, -34, 12, -16, -61, 13, 42, 25,
    -- layer=1 filter=97 channel=112
    -41, -33, -14, 14, -12, -19, 39, 42, 51,
    -- layer=1 filter=97 channel=113
    10, -13, -8, -2, -4, -10, 15, -7, 5,
    -- layer=1 filter=97 channel=114
    -49, -54, -47, -32, -15, -31, -19, 11, -30,
    -- layer=1 filter=97 channel=115
    8, 8, 6, 6, 16, 0, 10, 12, 3,
    -- layer=1 filter=97 channel=116
    -10, 3, 9, 6, 8, 0, -2, -6, -10,
    -- layer=1 filter=97 channel=117
    -122, -96, -24, 3, -59, -52, 9, 78, 29,
    -- layer=1 filter=97 channel=118
    -39, -74, -28, -21, -41, -18, 7, 8, 49,
    -- layer=1 filter=97 channel=119
    -39, -24, -4, -47, -76, 4, -15, -58, 15,
    -- layer=1 filter=97 channel=120
    8, -13, -18, -4, 4, -2, -2, 0, -19,
    -- layer=1 filter=97 channel=121
    1, 17, 30, -7, 0, -2, 8, 11, -9,
    -- layer=1 filter=97 channel=122
    -6, -3, 7, 4, 0, -5, -1, 8, -3,
    -- layer=1 filter=97 channel=123
    19, 11, 29, 4, 28, 25, 7, 30, 9,
    -- layer=1 filter=97 channel=124
    3, 2, -3, -1, -9, -13, -3, 2, -1,
    -- layer=1 filter=97 channel=125
    32, -3, -1, 4, -15, 3, 1, 17, 4,
    -- layer=1 filter=97 channel=126
    -49, -60, -22, -94, -89, -59, -78, -73, -28,
    -- layer=1 filter=97 channel=127
    -73, -114, -48, -28, -51, -47, 0, 3, 27,
    -- layer=1 filter=98 channel=0
    -1, -8, -26, -9, -5, -9, 11, 5, 3,
    -- layer=1 filter=98 channel=1
    -52, -42, -19, 16, 24, -7, -33, -13, -16,
    -- layer=1 filter=98 channel=2
    19, 5, -7, 24, -20, -13, 37, 6, -19,
    -- layer=1 filter=98 channel=3
    0, 1, 13, 6, 12, 3, 9, 14, 15,
    -- layer=1 filter=98 channel=4
    -1, -9, -6, -17, -7, 2, -6, -16, 7,
    -- layer=1 filter=98 channel=5
    -27, -36, -8, 40, 41, 5, -19, 7, 17,
    -- layer=1 filter=98 channel=6
    -20, 14, -7, -16, 23, 38, -30, 2, 0,
    -- layer=1 filter=98 channel=7
    -21, -2, -21, 10, 20, -19, 52, 28, 19,
    -- layer=1 filter=98 channel=8
    -20, -4, 3, 40, 26, -7, -26, -23, -16,
    -- layer=1 filter=98 channel=9
    -5, -14, -44, 0, -30, -9, -23, -92, -66,
    -- layer=1 filter=98 channel=10
    9, 16, -26, 28, 43, -22, 53, 48, 30,
    -- layer=1 filter=98 channel=11
    41, 8, 0, 36, 4, 8, 61, 32, 3,
    -- layer=1 filter=98 channel=12
    -17, -28, -24, 50, 28, 36, -22, -48, -45,
    -- layer=1 filter=98 channel=13
    1, 15, 29, -8, 10, 30, -45, -17, 0,
    -- layer=1 filter=98 channel=14
    0, -39, -45, -41, 24, -9, 35, 3, -18,
    -- layer=1 filter=98 channel=15
    -33, -14, 33, 24, 0, 15, -5, 18, -35,
    -- layer=1 filter=98 channel=16
    -28, -5, 9, 43, 16, -4, -29, -24, -8,
    -- layer=1 filter=98 channel=17
    -10, -1, 18, 13, 4, 6, -2, -1, -17,
    -- layer=1 filter=98 channel=18
    31, 25, 1, -22, -3, -36, 12, -28, -15,
    -- layer=1 filter=98 channel=19
    11, 2, -3, 33, -13, 0, -35, -40, -32,
    -- layer=1 filter=98 channel=20
    5, 32, 43, 5, 28, 40, -46, -16, -7,
    -- layer=1 filter=98 channel=21
    -22, 11, 42, -11, 37, 33, -30, 0, 25,
    -- layer=1 filter=98 channel=22
    1, 31, 28, 9, 26, 38, -23, -24, -14,
    -- layer=1 filter=98 channel=23
    -16, -48, -55, 29, -27, -20, 58, 21, 29,
    -- layer=1 filter=98 channel=24
    -27, -11, -12, -24, -9, -11, -6, 8, 14,
    -- layer=1 filter=98 channel=25
    -29, -9, 1, 22, 15, -3, 12, 12, 11,
    -- layer=1 filter=98 channel=26
    -15, -9, 5, 7, -16, -11, 4, -3, -16,
    -- layer=1 filter=98 channel=27
    57, 44, 21, 38, 32, 21, 56, 45, 34,
    -- layer=1 filter=98 channel=28
    -49, 11, -20, -9, 28, -7, 9, 9, -14,
    -- layer=1 filter=98 channel=29
    5, -18, -14, 17, 6, -15, 14, 4, -18,
    -- layer=1 filter=98 channel=30
    16, -17, -25, -31, -14, -32, -19, -34, -42,
    -- layer=1 filter=98 channel=31
    60, 40, 3, 25, 19, 7, 9, -12, 6,
    -- layer=1 filter=98 channel=32
    -38, -79, -63, -4, -11, -49, 18, 31, -11,
    -- layer=1 filter=98 channel=33
    -1, -21, -19, -26, -26, -18, -24, -7, -25,
    -- layer=1 filter=98 channel=34
    -49, -60, -56, -27, -27, -24, -11, -10, -12,
    -- layer=1 filter=98 channel=35
    -16, -7, -19, 16, 6, -11, 1, -10, -13,
    -- layer=1 filter=98 channel=36
    40, 9, 0, 22, -2, -4, 63, 24, 19,
    -- layer=1 filter=98 channel=37
    -23, -11, 22, 60, 23, 11, 3, 14, 36,
    -- layer=1 filter=98 channel=38
    -2, 23, 35, -19, 39, 32, -33, -3, 12,
    -- layer=1 filter=98 channel=39
    31, 28, 23, 37, 4, -1, 3, 18, 9,
    -- layer=1 filter=98 channel=40
    41, 44, 26, -4, 43, 31, -4, 13, 11,
    -- layer=1 filter=98 channel=41
    -45, -74, -97, 3, -66, -71, -15, -4, -72,
    -- layer=1 filter=98 channel=42
    40, 1, -2, 22, -3, -18, 13, -2, -39,
    -- layer=1 filter=98 channel=43
    -42, 0, -18, 40, 7, -5, -10, -8, -18,
    -- layer=1 filter=98 channel=44
    -36, -51, -29, 0, -13, -36, 13, 25, 3,
    -- layer=1 filter=98 channel=45
    -43, 5, 18, -8, 4, 26, -16, 19, 18,
    -- layer=1 filter=98 channel=46
    31, 2, 30, 44, 44, 14, 2, -11, -29,
    -- layer=1 filter=98 channel=47
    -16, -46, -31, 18, 20, 22, 50, 22, 29,
    -- layer=1 filter=98 channel=48
    -20, 22, 16, -13, 3, 18, -47, -6, 16,
    -- layer=1 filter=98 channel=49
    0, 12, 13, 19, 27, 16, 1, 8, 14,
    -- layer=1 filter=98 channel=50
    25, 8, 0, 1, -13, -18, -23, -8, -31,
    -- layer=1 filter=98 channel=51
    -15, 21, 16, -7, 33, 17, -3, 11, 11,
    -- layer=1 filter=98 channel=52
    21, 11, 19, 24, -3, 11, -15, -9, -2,
    -- layer=1 filter=98 channel=53
    35, 15, 10, 19, 8, 7, -2, 17, 5,
    -- layer=1 filter=98 channel=54
    -41, -23, -4, 43, -4, -15, 12, 9, 13,
    -- layer=1 filter=98 channel=55
    8, -20, -28, 33, 0, -4, 49, 40, 13,
    -- layer=1 filter=98 channel=56
    -9, -8, 9, 2, 7, 8, 8, -10, -6,
    -- layer=1 filter=98 channel=57
    22, 27, 14, 38, 66, 18, 40, 29, 35,
    -- layer=1 filter=98 channel=58
    -2, -49, -24, 30, -13, -40, 58, 7, 40,
    -- layer=1 filter=98 channel=59
    -6, -5, 5, 10, 5, -5, -22, -3, -14,
    -- layer=1 filter=98 channel=60
    3, -22, -18, -20, -2, -22, 8, -34, -8,
    -- layer=1 filter=98 channel=61
    7, 4, -1, 9, -11, -4, 6, -8, -11,
    -- layer=1 filter=98 channel=62
    -16, 0, 6, 46, 2, -10, -22, -1, -13,
    -- layer=1 filter=98 channel=63
    24, 6, -22, -5, -16, -40, 45, 4, 12,
    -- layer=1 filter=98 channel=64
    -27, -9, -2, -20, 10, 22, -31, -18, 5,
    -- layer=1 filter=98 channel=65
    -22, 33, 8, -26, 28, 26, -55, -10, -13,
    -- layer=1 filter=98 channel=66
    -1, -11, -22, 11, -1, -20, 44, 22, 5,
    -- layer=1 filter=98 channel=67
    -9, 33, 42, -6, 80, 71, -13, 29, 42,
    -- layer=1 filter=98 channel=68
    -64, -43, -25, 3, -48, -17, 25, 10, 12,
    -- layer=1 filter=98 channel=69
    -25, -18, 28, 28, 17, -7, -14, 4, -2,
    -- layer=1 filter=98 channel=70
    23, -21, -6, 9, 34, 10, -3, 36, 32,
    -- layer=1 filter=98 channel=71
    -33, 2, -27, -1, -25, -28, -14, 13, -1,
    -- layer=1 filter=98 channel=72
    26, -19, -20, 12, -23, 8, -23, -59, -66,
    -- layer=1 filter=98 channel=73
    -13, -21, -7, 3, -5, 0, -6, -7, 0,
    -- layer=1 filter=98 channel=74
    -11, 12, 0, -38, -23, 6, -3, -19, 19,
    -- layer=1 filter=98 channel=75
    6, -39, -35, -18, -40, -38, -42, -62, -77,
    -- layer=1 filter=98 channel=76
    -28, -24, -23, 11, -38, -17, 5, 4, -2,
    -- layer=1 filter=98 channel=77
    -41, -9, 24, -63, -1, 40, -51, -5, 14,
    -- layer=1 filter=98 channel=78
    -5, 11, -33, -6, 24, -6, 25, 34, 0,
    -- layer=1 filter=98 channel=79
    -8, 3, 37, 31, 19, -7, -34, -19, -12,
    -- layer=1 filter=98 channel=80
    7, -15, 1, 8, 7, 18, -2, -7, -24,
    -- layer=1 filter=98 channel=81
    -46, -26, -4, -19, -57, -13, -27, -20, 16,
    -- layer=1 filter=98 channel=82
    -23, 26, 22, -36, 33, 27, -29, 15, 13,
    -- layer=1 filter=98 channel=83
    -46, -28, 0, -8, -19, 2, -36, 8, -2,
    -- layer=1 filter=98 channel=84
    6, 10, -10, -19, -61, -39, -29, -47, -30,
    -- layer=1 filter=98 channel=85
    -27, -34, -52, 30, -19, -24, 45, 31, 44,
    -- layer=1 filter=98 channel=86
    42, 21, 7, 42, 34, 9, 32, 17, 12,
    -- layer=1 filter=98 channel=87
    41, 21, 19, 29, 19, -13, -17, -31, -30,
    -- layer=1 filter=98 channel=88
    5, 22, 18, 0, 42, 16, -4, 19, 14,
    -- layer=1 filter=98 channel=89
    -30, 26, 15, -28, 14, 39, -50, -17, 13,
    -- layer=1 filter=98 channel=90
    -51, -73, -6, -12, -49, -38, 24, 7, 10,
    -- layer=1 filter=98 channel=91
    -2, 17, 34, -4, 21, 36, -28, -13, 16,
    -- layer=1 filter=98 channel=92
    -46, -68, -3, -12, -39, -20, 3, 4, -24,
    -- layer=1 filter=98 channel=93
    -33, -11, -8, -34, -6, -1, -34, -10, 0,
    -- layer=1 filter=98 channel=94
    -11, -2, -15, -18, -10, -18, 5, -3, -16,
    -- layer=1 filter=98 channel=95
    17, -9, -30, -43, -56, -42, -10, -58, -36,
    -- layer=1 filter=98 channel=96
    -6, 2, -27, 0, -13, -28, 17, 0, 16,
    -- layer=1 filter=98 channel=97
    -20, -22, -9, -32, -33, -10, -17, -8, 1,
    -- layer=1 filter=98 channel=98
    -13, 17, 25, 36, 18, 2, -19, -6, 2,
    -- layer=1 filter=98 channel=99
    -29, 8, -17, -15, 33, -8, 30, 50, -7,
    -- layer=1 filter=98 channel=100
    21, 9, -1, 14, 10, 0, 37, 27, 33,
    -- layer=1 filter=98 channel=101
    0, 24, 15, -19, 29, 33, -29, -9, 6,
    -- layer=1 filter=98 channel=102
    -32, -14, -17, -55, -14, -4, -47, -26, -14,
    -- layer=1 filter=98 channel=103
    27, 18, 12, 24, 20, 1, 30, 23, 2,
    -- layer=1 filter=98 channel=104
    3, -26, -42, -3, -8, -44, 1, 40, -25,
    -- layer=1 filter=98 channel=105
    -13, -18, -23, -10, -20, -21, 21, -4, -13,
    -- layer=1 filter=98 channel=106
    -6, 3, 8, -20, 5, 28, -16, -16, -9,
    -- layer=1 filter=98 channel=107
    -9, -11, -9, -11, 5, -4, -4, -5, -11,
    -- layer=1 filter=98 channel=108
    -30, -61, -36, 0, 13, -50, 12, 41, -7,
    -- layer=1 filter=98 channel=109
    0, 8, -6, -7, 4, -1, 8, 7, -8,
    -- layer=1 filter=98 channel=110
    0, 1, -7, -7, 16, -7, -3, 13, -2,
    -- layer=1 filter=98 channel=111
    22, 4, -5, -33, 0, -36, 5, -19, -2,
    -- layer=1 filter=98 channel=112
    8, -20, -20, -38, -56, -61, -12, -25, 0,
    -- layer=1 filter=98 channel=113
    25, 17, 27, 46, 27, 9, 6, 30, -4,
    -- layer=1 filter=98 channel=114
    27, 9, 35, 46, 9, 0, -28, -11, -31,
    -- layer=1 filter=98 channel=115
    21, 21, -13, 42, 33, 6, 21, 30, 10,
    -- layer=1 filter=98 channel=116
    5, -8, -6, 8, -4, -10, -12, 2, -12,
    -- layer=1 filter=98 channel=117
    34, -2, -28, -31, 0, -26, -12, -2, -14,
    -- layer=1 filter=98 channel=118
    24, 13, 11, -23, -31, -9, -8, -34, 0,
    -- layer=1 filter=98 channel=119
    -61, -104, -59, -29, -54, -50, 17, 29, -19,
    -- layer=1 filter=98 channel=120
    -34, -7, 24, -6, 22, 37, -30, -12, 38,
    -- layer=1 filter=98 channel=121
    46, -3, -8, 10, 37, -23, 27, -16, -29,
    -- layer=1 filter=98 channel=122
    4, 9, 9, 6, -10, 8, 0, 6, 1,
    -- layer=1 filter=98 channel=123
    29, -24, -28, 1, -16, -34, 37, 11, -4,
    -- layer=1 filter=98 channel=124
    -2, -2, 10, 24, -3, -6, 11, -2, 13,
    -- layer=1 filter=98 channel=125
    17, 11, -6, -20, 49, 5, 19, 48, 44,
    -- layer=1 filter=98 channel=126
    -36, -37, 3, 17, 9, 17, 13, 23, 20,
    -- layer=1 filter=98 channel=127
    20, 8, -9, -32, -33, -32, -11, -30, -15,
    -- layer=1 filter=99 channel=0
    6, -20, -8, -4, -7, -1, -16, 0, 1,
    -- layer=1 filter=99 channel=1
    10, 0, 3, 10, 38, -12, 1, -7, -14,
    -- layer=1 filter=99 channel=2
    -8, 16, 14, -1, 1, -12, 0, -15, -21,
    -- layer=1 filter=99 channel=3
    -7, 2, -12, -8, -11, -11, -7, -1, 0,
    -- layer=1 filter=99 channel=4
    -5, 1, -4, 1, -2, 7, 0, 12, -1,
    -- layer=1 filter=99 channel=5
    8, -1, 10, 28, 38, -14, 9, 3, -14,
    -- layer=1 filter=99 channel=6
    9, 9, -9, -16, -22, 3, -18, 9, -36,
    -- layer=1 filter=99 channel=7
    -16, 28, -2, -5, 42, 9, 17, -5, 8,
    -- layer=1 filter=99 channel=8
    42, 22, 27, 22, 47, -21, 35, 3, 2,
    -- layer=1 filter=99 channel=9
    5, -4, 17, 13, 9, 0, -36, 17, -6,
    -- layer=1 filter=99 channel=10
    -8, 24, 16, 0, 29, 10, 10, -15, 4,
    -- layer=1 filter=99 channel=11
    -8, -9, -9, -5, 2, 4, 26, 28, 18,
    -- layer=1 filter=99 channel=12
    3, 7, -21, -28, -25, -21, 4, 41, -42,
    -- layer=1 filter=99 channel=13
    -10, 1, -6, -10, 5, -6, -8, 10, 15,
    -- layer=1 filter=99 channel=14
    -37, 12, -23, -15, -11, -7, -31, -36, -24,
    -- layer=1 filter=99 channel=15
    10, 16, 12, 24, 42, -5, 38, 25, 9,
    -- layer=1 filter=99 channel=16
    33, 14, 19, 27, 45, 2, 23, 7, 1,
    -- layer=1 filter=99 channel=17
    -7, 0, 0, -16, 3, -15, 7, 13, 3,
    -- layer=1 filter=99 channel=18
    1, -4, -4, 18, 11, -19, -6, 5, 4,
    -- layer=1 filter=99 channel=19
    16, 52, 41, 78, 53, 36, 46, 67, 34,
    -- layer=1 filter=99 channel=20
    -4, -5, 5, -4, -2, -7, -3, 1, -1,
    -- layer=1 filter=99 channel=21
    -18, -17, -4, -24, 0, 11, -3, -1, -5,
    -- layer=1 filter=99 channel=22
    -13, -9, 3, -8, 26, 14, 15, 31, -6,
    -- layer=1 filter=99 channel=23
    8, 69, -8, 2, 27, 7, 14, 2, 0,
    -- layer=1 filter=99 channel=24
    5, -13, 11, 7, -7, -20, -3, -21, 2,
    -- layer=1 filter=99 channel=25
    7, 28, 18, 22, 58, 11, 42, -9, -1,
    -- layer=1 filter=99 channel=26
    -2, 3, 5, 6, 22, -11, -8, -18, -7,
    -- layer=1 filter=99 channel=27
    4, -10, -13, 0, -20, -31, 2, -3, 0,
    -- layer=1 filter=99 channel=28
    -12, -2, 10, -3, 28, 11, 20, -21, -9,
    -- layer=1 filter=99 channel=29
    0, 12, 13, -7, -7, 2, -2, 2, 16,
    -- layer=1 filter=99 channel=30
    -9, -10, -8, 36, -1, 1, -10, 11, 1,
    -- layer=1 filter=99 channel=31
    17, 6, -5, 16, -8, -3, -13, 2, -25,
    -- layer=1 filter=99 channel=32
    6, 17, 8, 0, 13, 12, 6, -10, 23,
    -- layer=1 filter=99 channel=33
    1, -12, 4, 15, 9, -2, 8, 0, -10,
    -- layer=1 filter=99 channel=34
    8, -2, 3, 0, 9, -9, 2, -6, -1,
    -- layer=1 filter=99 channel=35
    -8, 3, 3, 4, 4, -1, 18, 10, 0,
    -- layer=1 filter=99 channel=36
    -4, -19, -12, -8, -2, 3, 19, -4, -1,
    -- layer=1 filter=99 channel=37
    18, 5, 24, 39, 35, -18, 11, -4, 2,
    -- layer=1 filter=99 channel=38
    -7, -17, 7, -4, -8, 1, -5, 12, 13,
    -- layer=1 filter=99 channel=39
    3, 1, 5, -7, -2, -11, 5, -5, -8,
    -- layer=1 filter=99 channel=40
    -8, 6, 3, 3, -8, -3, -2, -8, -8,
    -- layer=1 filter=99 channel=41
    0, 34, -6, 19, 37, 20, 4, 24, 43,
    -- layer=1 filter=99 channel=42
    -24, 23, -1, 3, -3, -1, -10, -25, -10,
    -- layer=1 filter=99 channel=43
    24, 6, 17, 0, 39, -25, 27, 6, -21,
    -- layer=1 filter=99 channel=44
    -10, 7, -3, -8, 13, 6, -3, -40, 7,
    -- layer=1 filter=99 channel=45
    2, -10, 12, -7, 5, -4, -3, -3, 1,
    -- layer=1 filter=99 channel=46
    -25, 1, -17, 25, 25, -8, 30, 27, 3,
    -- layer=1 filter=99 channel=47
    17, 59, -6, 28, 27, -4, -18, 3, 8,
    -- layer=1 filter=99 channel=48
    -14, -21, -24, -3, -17, -17, -5, 3, -4,
    -- layer=1 filter=99 channel=49
    12, -1, -2, 6, -6, 7, -16, 18, -16,
    -- layer=1 filter=99 channel=50
    4, -10, 16, -7, -11, -27, -4, 4, -1,
    -- layer=1 filter=99 channel=51
    -22, -4, -7, -22, -7, 16, 9, -4, 1,
    -- layer=1 filter=99 channel=52
    11, -14, 12, -7, 10, -8, 0, -6, -5,
    -- layer=1 filter=99 channel=53
    0, 7, 3, 8, 11, 6, 19, 5, 22,
    -- layer=1 filter=99 channel=54
    9, 30, 6, 34, 55, 3, 49, -6, 8,
    -- layer=1 filter=99 channel=55
    18, 1, 5, 14, -6, 0, 7, 8, -5,
    -- layer=1 filter=99 channel=56
    12, -3, 4, -4, 10, 3, 2, 6, 4,
    -- layer=1 filter=99 channel=57
    -7, 8, 29, 8, 31, 13, 22, -17, 9,
    -- layer=1 filter=99 channel=58
    18, 70, 1, 35, 43, 23, 11, -5, 0,
    -- layer=1 filter=99 channel=59
    0, 0, 8, 2, 16, 11, 0, 15, 15,
    -- layer=1 filter=99 channel=60
    2, 20, 19, 5, 8, 9, 7, 19, 18,
    -- layer=1 filter=99 channel=61
    1, 7, -13, 7, -5, -4, 10, -1, 1,
    -- layer=1 filter=99 channel=62
    28, 37, 41, 32, 53, -9, 40, 1, 5,
    -- layer=1 filter=99 channel=63
    -12, -22, -19, -16, -21, -8, -12, -10, 11,
    -- layer=1 filter=99 channel=64
    -11, -7, 5, 0, 8, 2, -4, 13, -3,
    -- layer=1 filter=99 channel=65
    -17, -31, -15, -14, -10, 1, -4, 13, 9,
    -- layer=1 filter=99 channel=66
    -13, -17, -12, -19, -12, 0, 3, -10, -22,
    -- layer=1 filter=99 channel=67
    8, -13, -11, -13, -2, -25, 3, 21, 16,
    -- layer=1 filter=99 channel=68
    12, 15, 13, 0, 4, 28, 7, -19, 7,
    -- layer=1 filter=99 channel=69
    3, -1, 5, 4, 20, -42, 16, -11, -17,
    -- layer=1 filter=99 channel=70
    7, -12, -9, -2, -3, -23, -22, -3, -43,
    -- layer=1 filter=99 channel=71
    -11, -1, -9, -10, 0, -18, -4, -5, 4,
    -- layer=1 filter=99 channel=72
    -12, 1, -16, 40, 24, 11, 17, 40, -3,
    -- layer=1 filter=99 channel=73
    -2, -6, 7, -4, 4, 2, -13, -12, -8,
    -- layer=1 filter=99 channel=74
    10, 9, 7, 15, 13, 4, -3, -7, 18,
    -- layer=1 filter=99 channel=75
    -44, -16, -50, -2, -32, -28, -33, -1, -39,
    -- layer=1 filter=99 channel=76
    -16, 3, -31, -13, -9, -9, 2, 0, 13,
    -- layer=1 filter=99 channel=77
    -8, -24, -5, -16, -19, -17, -1, 4, 15,
    -- layer=1 filter=99 channel=78
    -5, -13, 3, -8, 10, -1, 0, -6, 7,
    -- layer=1 filter=99 channel=79
    21, 7, 4, 16, 38, -14, 6, 0, -9,
    -- layer=1 filter=99 channel=80
    5, 5, -1, 6, 11, 18, 20, 12, 9,
    -- layer=1 filter=99 channel=81
    -5, 0, -6, -9, -8, -22, -4, -6, -18,
    -- layer=1 filter=99 channel=82
    -25, -21, -9, -35, -8, -12, -18, 4, -2,
    -- layer=1 filter=99 channel=83
    -21, 0, 18, -18, -15, -25, 8, 6, 4,
    -- layer=1 filter=99 channel=84
    24, 36, -9, 21, 35, -15, 10, 9, 7,
    -- layer=1 filter=99 channel=85
    18, 73, -1, 28, 40, -1, 3, 6, -9,
    -- layer=1 filter=99 channel=86
    -11, -9, -9, -1, -3, 3, 22, 18, 9,
    -- layer=1 filter=99 channel=87
    8, 18, 16, 65, 25, 12, 20, 56, 19,
    -- layer=1 filter=99 channel=88
    -6, -3, -7, 10, 5, 6, 21, 17, -1,
    -- layer=1 filter=99 channel=89
    -2, -4, -16, -32, -14, 1, -16, 3, -2,
    -- layer=1 filter=99 channel=90
    -10, 10, 12, -18, 2, 2, -8, -25, -1,
    -- layer=1 filter=99 channel=91
    -14, -18, -12, -19, -5, 9, 0, 19, 1,
    -- layer=1 filter=99 channel=92
    -17, -9, 4, -6, 7, 13, 10, -4, 42,
    -- layer=1 filter=99 channel=93
    -16, -26, -18, -22, -9, -15, -3, -11, 0,
    -- layer=1 filter=99 channel=94
    5, -19, -4, -5, -6, 15, -6, 3, 1,
    -- layer=1 filter=99 channel=95
    21, 8, -14, 10, 0, -6, -1, -11, 11,
    -- layer=1 filter=99 channel=96
    -1, -14, -5, 3, 16, 8, 9, -8, -15,
    -- layer=1 filter=99 channel=97
    -6, -24, 0, -23, -15, 3, -9, -9, 0,
    -- layer=1 filter=99 channel=98
    7, -2, 10, 4, 36, -7, 23, -3, -15,
    -- layer=1 filter=99 channel=99
    5, -5, 41, -6, -14, -3, 2, -31, 0,
    -- layer=1 filter=99 channel=100
    3, 1, -21, -1, -1, 8, 25, 27, 33,
    -- layer=1 filter=99 channel=101
    0, -5, -14, -19, 0, -1, 1, 13, 1,
    -- layer=1 filter=99 channel=102
    -21, -26, 1, -22, -16, -12, -20, 0, -3,
    -- layer=1 filter=99 channel=103
    -2, -18, -20, 4, 10, 4, 12, 15, 15,
    -- layer=1 filter=99 channel=104
    -2, 26, 0, 9, 21, -6, -8, 4, 14,
    -- layer=1 filter=99 channel=105
    2, -15, -1, -13, -20, -4, 0, -1, -15,
    -- layer=1 filter=99 channel=106
    3, 12, -19, -1, -7, 0, -4, -2, 8,
    -- layer=1 filter=99 channel=107
    -12, 0, -24, -22, -4, -3, -1, 0, -1,
    -- layer=1 filter=99 channel=108
    -7, 16, -13, -24, 17, -3, 3, -10, -1,
    -- layer=1 filter=99 channel=109
    11, 0, -5, -12, 3, 3, 6, -1, 0,
    -- layer=1 filter=99 channel=110
    -8, -1, -7, -10, 4, -3, 0, -9, 8,
    -- layer=1 filter=99 channel=111
    3, 12, -3, 25, 16, -31, -10, 8, 2,
    -- layer=1 filter=99 channel=112
    40, 31, -33, 27, 14, -14, 30, 20, 26,
    -- layer=1 filter=99 channel=113
    -15, 20, -15, -23, -3, -6, -26, -14, -32,
    -- layer=1 filter=99 channel=114
    23, 11, 4, 21, 16, -23, 30, 21, -2,
    -- layer=1 filter=99 channel=115
    -15, 5, 8, 5, 21, 13, 24, 1, 18,
    -- layer=1 filter=99 channel=116
    -6, 3, -2, -10, -8, -10, -7, -4, -5,
    -- layer=1 filter=99 channel=117
    19, 27, -18, 40, 5, -9, 40, 14, 23,
    -- layer=1 filter=99 channel=118
    10, 11, -13, 25, 1, -30, -17, -11, 3,
    -- layer=1 filter=99 channel=119
    -1, 17, 4, 7, 22, 6, -1, 0, 7,
    -- layer=1 filter=99 channel=120
    -8, -7, -1, -15, 13, -9, -1, 0, 8,
    -- layer=1 filter=99 channel=121
    -18, -9, -14, 5, -2, -4, -2, 17, 7,
    -- layer=1 filter=99 channel=122
    -4, 1, -1, 10, 3, -6, 0, -3, -9,
    -- layer=1 filter=99 channel=123
    -16, 3, -15, 6, -6, -13, -3, 15, 3,
    -- layer=1 filter=99 channel=124
    6, 10, 13, 16, 7, 6, 27, 13, 21,
    -- layer=1 filter=99 channel=125
    2, -19, -25, 15, -1, -2, -22, 0, -9,
    -- layer=1 filter=99 channel=126
    22, 14, 6, 2, 23, -21, 7, 2, -24,
    -- layer=1 filter=99 channel=127
    0, 3, -27, 11, 4, -12, 9, -8, 0,
    -- layer=1 filter=100 channel=0
    9, 3, 11, 5, 3, -12, 5, 8, -4,
    -- layer=1 filter=100 channel=1
    -19, 0, -18, 6, 7, -6, -14, -13, 22,
    -- layer=1 filter=100 channel=2
    -18, 3, 43, 0, 2, 13, 7, 16, 25,
    -- layer=1 filter=100 channel=3
    -11, -3, 0, -1, 7, 5, 1, 4, 5,
    -- layer=1 filter=100 channel=4
    -8, 9, 7, -7, -8, 5, 5, -4, -4,
    -- layer=1 filter=100 channel=5
    -13, -2, -10, 5, 24, 22, -27, -10, 15,
    -- layer=1 filter=100 channel=6
    4, -4, -24, -10, -12, -1, -26, -7, 41,
    -- layer=1 filter=100 channel=7
    -49, -60, 12, -92, -50, -70, -68, -39, -101,
    -- layer=1 filter=100 channel=8
    -31, -11, -27, 36, 33, -5, -30, 1, 24,
    -- layer=1 filter=100 channel=9
    -38, -32, 32, 10, 8, 44, -21, -6, 11,
    -- layer=1 filter=100 channel=10
    -56, -50, 10, -91, -60, -101, -68, -68, -86,
    -- layer=1 filter=100 channel=11
    13, 12, 4, 14, 9, -6, 7, 8, -11,
    -- layer=1 filter=100 channel=12
    -5, -8, 17, -4, -29, 19, -18, 3, 2,
    -- layer=1 filter=100 channel=13
    -13, -19, -33, -27, 0, -31, -15, 21, 7,
    -- layer=1 filter=100 channel=14
    -70, -46, 35, -106, -29, -18, -71, -23, -56,
    -- layer=1 filter=100 channel=15
    17, 12, -37, -11, 14, -1, -8, 5, 47,
    -- layer=1 filter=100 channel=16
    -12, -8, -22, 29, 32, 0, -13, 1, 29,
    -- layer=1 filter=100 channel=17
    26, 1, -2, 20, -2, -17, 16, 2, 1,
    -- layer=1 filter=100 channel=18
    -24, -19, 14, 9, 16, 12, 3, -16, 10,
    -- layer=1 filter=100 channel=19
    -37, -22, -7, -1, 46, 28, -17, -1, 41,
    -- layer=1 filter=100 channel=20
    -22, -4, -27, -21, -20, -18, -4, -1, -18,
    -- layer=1 filter=100 channel=21
    -37, -41, -54, -20, -22, -12, -21, -40, -27,
    -- layer=1 filter=100 channel=22
    -37, -36, -40, -16, 2, -22, -20, -17, 6,
    -- layer=1 filter=100 channel=23
    -9, -4, -22, -21, -17, -42, 19, -3, 5,
    -- layer=1 filter=100 channel=24
    -8, -44, -10, -17, 21, 1, 3, 13, 25,
    -- layer=1 filter=100 channel=25
    -52, -35, -30, 0, -49, -45, -95, -63, -66,
    -- layer=1 filter=100 channel=26
    2, -17, -3, -1, 42, -26, 20, 34, 46,
    -- layer=1 filter=100 channel=27
    -33, -20, -19, -35, -22, -25, -49, -39, -24,
    -- layer=1 filter=100 channel=28
    -42, -53, 16, -47, -57, -75, -66, -35, -65,
    -- layer=1 filter=100 channel=29
    -31, -13, -6, -33, -30, 5, -26, -31, -7,
    -- layer=1 filter=100 channel=30
    -5, -17, 28, 3, 28, 19, -21, 0, 10,
    -- layer=1 filter=100 channel=31
    -39, -37, -1, -30, -19, -13, -24, -12, -5,
    -- layer=1 filter=100 channel=32
    5, 9, 0, 9, 25, -25, -7, 33, 35,
    -- layer=1 filter=100 channel=33
    8, -8, 3, -6, 4, -10, 0, 5, 2,
    -- layer=1 filter=100 channel=34
    7, 12, 27, 3, 8, 15, -10, 2, -11,
    -- layer=1 filter=100 channel=35
    -4, 2, -16, 0, -7, -15, 2, 4, -6,
    -- layer=1 filter=100 channel=36
    29, 20, 15, 31, 23, 14, 28, 11, 0,
    -- layer=1 filter=100 channel=37
    0, -2, -10, 29, 16, 7, -16, -7, 27,
    -- layer=1 filter=100 channel=38
    -34, -34, -23, -46, -28, -36, -39, -16, -12,
    -- layer=1 filter=100 channel=39
    9, 2, -1, 27, 3, -2, 6, 0, 1,
    -- layer=1 filter=100 channel=40
    -64, -57, -27, -50, -57, -39, -30, -3, 4,
    -- layer=1 filter=100 channel=41
    5, 0, 6, 15, 38, 15, 14, 27, 22,
    -- layer=1 filter=100 channel=42
    -22, -3, 38, -31, -17, 21, 25, -22, 20,
    -- layer=1 filter=100 channel=43
    -14, -25, -35, 28, 35, -12, -36, -14, 1,
    -- layer=1 filter=100 channel=44
    -9, 19, -12, 7, 42, -13, 14, 44, 42,
    -- layer=1 filter=100 channel=45
    -27, -24, -20, -30, 7, -34, -42, 5, 5,
    -- layer=1 filter=100 channel=46
    -46, -8, -1, -8, 34, 28, -34, -21, 19,
    -- layer=1 filter=100 channel=47
    -28, -15, -53, -35, -23, -23, -9, -13, 10,
    -- layer=1 filter=100 channel=48
    -7, -19, -11, -10, -24, -9, -6, -23, -21,
    -- layer=1 filter=100 channel=49
    -24, -17, 0, -19, -33, 3, -25, -9, -11,
    -- layer=1 filter=100 channel=50
    -21, -19, 9, -17, -32, -8, -3, -7, 2,
    -- layer=1 filter=100 channel=51
    -28, -33, -16, -49, -20, -33, -23, -46, -26,
    -- layer=1 filter=100 channel=52
    15, -3, -12, -8, -6, 9, 9, 18, 6,
    -- layer=1 filter=100 channel=53
    -16, -4, 10, 0, -6, -3, -18, -17, -10,
    -- layer=1 filter=100 channel=54
    -42, -4, -23, -4, -27, -43, -53, -52, -6,
    -- layer=1 filter=100 channel=55
    20, 5, -6, 31, 19, 1, 0, 0, 4,
    -- layer=1 filter=100 channel=56
    -1, 5, -8, 8, -11, -2, 3, -12, -3,
    -- layer=1 filter=100 channel=57
    -84, -52, 1, -97, -55, -96, -74, -50, -74,
    -- layer=1 filter=100 channel=58
    -93, -52, -35, -54, -92, -107, -7, -62, -49,
    -- layer=1 filter=100 channel=59
    5, -3, 2, -12, -12, 1, -4, -5, -11,
    -- layer=1 filter=100 channel=60
    -6, 9, 3, -5, 1, 14, -8, -10, 4,
    -- layer=1 filter=100 channel=61
    -7, 9, -5, 10, -8, -9, 5, 1, -7,
    -- layer=1 filter=100 channel=62
    -16, -17, -19, 32, 30, 11, -12, -5, 15,
    -- layer=1 filter=100 channel=63
    8, 17, 13, 33, 8, 11, 25, 0, -3,
    -- layer=1 filter=100 channel=64
    -10, 8, 9, 7, 6, -7, 0, -8, 7,
    -- layer=1 filter=100 channel=65
    -1, 0, 0, -2, -5, -12, -10, -23, -10,
    -- layer=1 filter=100 channel=66
    19, 14, -1, 22, 11, 5, 12, -8, 1,
    -- layer=1 filter=100 channel=67
    -34, -48, -63, 8, -27, -18, -11, -16, 0,
    -- layer=1 filter=100 channel=68
    -3, 4, 3, 13, 39, -22, 27, 25, 19,
    -- layer=1 filter=100 channel=69
    16, -11, -14, 20, 36, -15, 3, 31, 38,
    -- layer=1 filter=100 channel=70
    26, 39, -7, -21, -15, 5, -18, -14, 3,
    -- layer=1 filter=100 channel=71
    -29, -10, -17, 9, 16, 15, -17, 0, 12,
    -- layer=1 filter=100 channel=72
    -12, -16, -2, 24, 37, 29, -9, 3, 42,
    -- layer=1 filter=100 channel=73
    1, -6, 0, -6, 1, 0, -7, -2, 4,
    -- layer=1 filter=100 channel=74
    -38, 31, -1, -4, 16, -6, -3, -1, 16,
    -- layer=1 filter=100 channel=75
    -39, -25, -11, -30, -2, 19, -29, 6, 18,
    -- layer=1 filter=100 channel=76
    0, 0, -4, 20, 9, 0, 17, 9, 7,
    -- layer=1 filter=100 channel=77
    -19, -21, -28, -15, -14, -8, -15, -3, 0,
    -- layer=1 filter=100 channel=78
    9, -5, 14, -3, -12, -10, -4, -4, -9,
    -- layer=1 filter=100 channel=79
    -27, -3, -11, 38, 26, 5, -9, 5, 30,
    -- layer=1 filter=100 channel=80
    -5, 7, 8, -10, 6, 9, 3, -1, -7,
    -- layer=1 filter=100 channel=81
    -42, -47, -30, 18, 10, 3, -13, -2, 9,
    -- layer=1 filter=100 channel=82
    -35, -44, -50, -41, -48, -34, -21, -28, -3,
    -- layer=1 filter=100 channel=83
    1, -31, -25, -16, 22, -28, -11, 30, 33,
    -- layer=1 filter=100 channel=84
    -11, 12, 34, 15, 8, 21, 5, 10, 28,
    -- layer=1 filter=100 channel=85
    -37, -8, -30, -45, -20, -62, -10, -38, -3,
    -- layer=1 filter=100 channel=86
    28, 20, 1, 18, 2, 4, 1, -1, -10,
    -- layer=1 filter=100 channel=87
    -50, -25, 24, -10, 32, 39, -45, -14, 59,
    -- layer=1 filter=100 channel=88
    -24, -19, -3, -23, -8, -12, -9, -15, -14,
    -- layer=1 filter=100 channel=89
    -51, -10, -27, -25, -9, -19, -25, 1, -3,
    -- layer=1 filter=100 channel=90
    0, -26, -32, -2, 42, -41, 9, 34, 32,
    -- layer=1 filter=100 channel=91
    -16, -2, -12, -34, -30, -36, -40, -31, -26,
    -- layer=1 filter=100 channel=92
    -4, 25, -34, -64, 16, -38, -16, 53, 14,
    -- layer=1 filter=100 channel=93
    1, 1, -2, -7, 4, -13, -5, -4, 3,
    -- layer=1 filter=100 channel=94
    18, 0, 11, 5, 8, 3, 16, 6, -11,
    -- layer=1 filter=100 channel=95
    -5, 17, 29, 21, 32, 24, 1, 19, 17,
    -- layer=1 filter=100 channel=96
    -3, 0, 0, 0, 0, 2, 5, 8, 10,
    -- layer=1 filter=100 channel=97
    12, 15, 7, 15, 1, 0, 5, 11, -9,
    -- layer=1 filter=100 channel=98
    -13, -32, -23, 26, 13, -33, -25, -2, 20,
    -- layer=1 filter=100 channel=99
    -67, -77, -15, -101, -80, -86, -41, 0, -64,
    -- layer=1 filter=100 channel=100
    11, 17, -3, 23, 10, 16, 7, -10, -15,
    -- layer=1 filter=100 channel=101
    -18, -11, -8, -30, -41, -24, -20, -31, -11,
    -- layer=1 filter=100 channel=102
    13, 19, 12, 8, -18, -5, 10, -5, -15,
    -- layer=1 filter=100 channel=103
    -22, 0, -10, -10, -12, -2, -8, -32, -19,
    -- layer=1 filter=100 channel=104
    -49, -17, -12, -13, 8, -21, 10, -17, 26,
    -- layer=1 filter=100 channel=105
    5, 14, 8, 14, 9, -7, -1, 10, -10,
    -- layer=1 filter=100 channel=106
    -31, -2, -28, -31, 0, -27, -24, 0, -9,
    -- layer=1 filter=100 channel=107
    17, 6, 9, 4, -6, 5, -6, -1, -1,
    -- layer=1 filter=100 channel=108
    9, -17, -37, -14, 41, -28, -2, 26, 21,
    -- layer=1 filter=100 channel=109
    -2, -10, 7, -2, 3, -7, -7, -1, -3,
    -- layer=1 filter=100 channel=110
    -9, 5, 0, 0, 6, -5, -12, -12, 6,
    -- layer=1 filter=100 channel=111
    0, 10, 47, -3, 18, 19, 12, -4, 4,
    -- layer=1 filter=100 channel=112
    -9, 8, 7, 11, 5, 0, 18, -3, 7,
    -- layer=1 filter=100 channel=113
    -6, 5, 5, -10, -29, 24, -5, -33, 4,
    -- layer=1 filter=100 channel=114
    1, 0, -16, 33, 38, 7, -16, -16, 17,
    -- layer=1 filter=100 channel=115
    8, 14, 20, 3, -3, -16, -12, -22, -34,
    -- layer=1 filter=100 channel=116
    -8, -10, 1, -5, 10, 1, -8, -1, -9,
    -- layer=1 filter=100 channel=117
    -6, -8, 32, -11, -30, -19, 13, -19, -26,
    -- layer=1 filter=100 channel=118
    -13, 5, 12, 8, 36, 22, -11, 3, 23,
    -- layer=1 filter=100 channel=119
    23, -4, -10, -3, 45, -19, 18, 31, 35,
    -- layer=1 filter=100 channel=120
    -20, -35, -31, -11, -45, -37, -39, -56, -44,
    -- layer=1 filter=100 channel=121
    -22, -22, -1, -21, 15, 22, -45, -19, 0,
    -- layer=1 filter=100 channel=122
    -2, -4, 6, 6, -3, 0, 7, -9, 10,
    -- layer=1 filter=100 channel=123
    -8, 3, -12, -10, 7, 28, -19, -4, -8,
    -- layer=1 filter=100 channel=124
    -11, -12, 4, -6, -8, -12, 0, 0, 3,
    -- layer=1 filter=100 channel=125
    13, 10, -2, 7, -4, -14, -20, -47, 13,
    -- layer=1 filter=100 channel=126
    -24, -28, -7, -4, 2, -31, -14, 28, 15,
    -- layer=1 filter=100 channel=127
    5, 7, 35, 8, 31, 15, -1, 13, 17,
    -- layer=1 filter=101 channel=0
    -31, -21, -8, -9, -37, -20, -20, -11, -14,
    -- layer=1 filter=101 channel=1
    4, -8, -24, -26, -16, -11, -52, -2, 29,
    -- layer=1 filter=101 channel=2
    -33, -11, 20, -2, 17, 6, 10, -24, -31,
    -- layer=1 filter=101 channel=3
    0, -8, 3, 2, -1, 8, 0, 4, 2,
    -- layer=1 filter=101 channel=4
    -2, -1, 4, -4, 7, 0, -12, 1, 0,
    -- layer=1 filter=101 channel=5
    -8, 12, -32, -28, -4, 16, -65, -24, 46,
    -- layer=1 filter=101 channel=6
    -11, -18, -1, -9, -4, 12, 8, -17, -25,
    -- layer=1 filter=101 channel=7
    -33, -24, -1, -9, -25, -19, 31, 14, -17,
    -- layer=1 filter=101 channel=8
    9, -6, -26, -29, -10, -17, -54, -17, 36,
    -- layer=1 filter=101 channel=9
    -31, -4, -14, 15, -7, -24, 0, -21, -29,
    -- layer=1 filter=101 channel=10
    -18, -18, 7, -1, -18, -2, 35, 19, -3,
    -- layer=1 filter=101 channel=11
    -39, -16, -22, -28, -35, -11, -15, -32, -24,
    -- layer=1 filter=101 channel=12
    20, -51, -12, -3, -14, 21, 9, 13, -16,
    -- layer=1 filter=101 channel=13
    8, 39, -3, 6, 38, 4, 8, 17, 27,
    -- layer=1 filter=101 channel=14
    -23, -31, 11, 12, -7, -1, 21, 28, -17,
    -- layer=1 filter=101 channel=15
    -3, 41, -21, -28, -4, 26, -45, -20, 71,
    -- layer=1 filter=101 channel=16
    -24, -20, -37, -34, -7, -4, -79, -19, 40,
    -- layer=1 filter=101 channel=17
    2, -11, -29, -23, 7, -36, -18, -2, 5,
    -- layer=1 filter=101 channel=18
    -21, -22, -45, 10, -26, 16, -13, -23, -31,
    -- layer=1 filter=101 channel=19
    -29, -32, -1, 0, 22, 0, 9, -18, -5,
    -- layer=1 filter=101 channel=20
    -9, 9, -13, -6, -6, -17, -8, 11, 10,
    -- layer=1 filter=101 channel=21
    3, -18, 21, 10, 0, -2, 10, -5, -4,
    -- layer=1 filter=101 channel=22
    13, 10, 9, -1, 12, -8, -30, 17, 42,
    -- layer=1 filter=101 channel=23
    36, 8, -4, -28, -55, 19, 12, -28, 11,
    -- layer=1 filter=101 channel=24
    6, 28, -6, -17, 35, -3, -34, -7, 24,
    -- layer=1 filter=101 channel=25
    -31, -21, -3, -7, -21, -24, 11, 0, -23,
    -- layer=1 filter=101 channel=26
    -35, 15, -27, -26, 29, -8, -36, -30, 24,
    -- layer=1 filter=101 channel=27
    -15, -23, 21, 0, -19, -10, -12, -21, -59,
    -- layer=1 filter=101 channel=28
    -30, -28, 11, 0, -12, 1, 22, 20, -10,
    -- layer=1 filter=101 channel=29
    -11, -4, -3, -11, -17, 11, -23, -17, -4,
    -- layer=1 filter=101 channel=30
    -37, -41, -19, 28, 10, 0, 3, -16, -50,
    -- layer=1 filter=101 channel=31
    -15, -60, -6, 2, -31, 32, 0, -9, -7,
    -- layer=1 filter=101 channel=32
    -12, 42, -4, -11, 28, 31, -28, -44, 34,
    -- layer=1 filter=101 channel=33
    18, -11, 8, -1, -1, 0, 5, -2, 14,
    -- layer=1 filter=101 channel=34
    4, 0, -2, 23, -9, 5, -3, -14, -12,
    -- layer=1 filter=101 channel=35
    -7, -7, 4, -10, -4, 0, -2, 7, 1,
    -- layer=1 filter=101 channel=36
    -46, -34, -21, -19, -22, -9, -30, -26, -31,
    -- layer=1 filter=101 channel=37
    -27, -9, -19, -31, 5, -6, -51, -13, 46,
    -- layer=1 filter=101 channel=38
    3, 1, -7, 19, 6, 0, 7, 18, -1,
    -- layer=1 filter=101 channel=39
    3, -19, -8, -2, 7, -19, -10, 4, 28,
    -- layer=1 filter=101 channel=40
    -39, -46, -27, 6, -30, -5, 22, -24, -44,
    -- layer=1 filter=101 channel=41
    -9, 17, -28, 2, 6, 4, 3, -33, 9,
    -- layer=1 filter=101 channel=42
    -27, -15, 36, -36, -8, -1, 5, -3, -39,
    -- layer=1 filter=101 channel=43
    -9, -23, -9, -25, -19, -33, -46, -15, 36,
    -- layer=1 filter=101 channel=44
    -19, 38, -34, -3, 14, 16, -30, -41, 16,
    -- layer=1 filter=101 channel=45
    10, 45, -39, -20, 35, -4, -28, -7, 62,
    -- layer=1 filter=101 channel=46
    -28, -68, -26, -33, -47, 11, -33, -48, -31,
    -- layer=1 filter=101 channel=47
    15, 2, -21, -23, -48, 47, 1, -40, 5,
    -- layer=1 filter=101 channel=48
    -5, -7, 5, 2, -20, -22, 1, -1, -20,
    -- layer=1 filter=101 channel=49
    -12, 16, 2, -12, -25, 34, 12, -28, -10,
    -- layer=1 filter=101 channel=50
    6, -8, -2, 7, -1, 1, -5, -10, 8,
    -- layer=1 filter=101 channel=51
    -17, -16, 17, 9, -26, 10, 21, 3, -26,
    -- layer=1 filter=101 channel=52
    -3, 7, -22, -10, 13, 5, 4, 2, -2,
    -- layer=1 filter=101 channel=53
    5, -8, -10, -10, 6, -3, 1, -1, 5,
    -- layer=1 filter=101 channel=54
    -42, -26, -4, -20, -20, -30, 40, -24, -33,
    -- layer=1 filter=101 channel=55
    -53, -24, -6, -59, -18, 17, -57, -54, 0,
    -- layer=1 filter=101 channel=56
    10, -3, 3, 3, 6, -8, -6, -2, -10,
    -- layer=1 filter=101 channel=57
    -28, -27, 12, 9, -10, -4, 35, 2, -29,
    -- layer=1 filter=101 channel=58
    -3, -1, -21, -23, -49, 11, 34, -17, -18,
    -- layer=1 filter=101 channel=59
    -8, -3, -7, 2, 6, -8, 2, 4, -8,
    -- layer=1 filter=101 channel=60
    -15, 18, 12, 17, -11, 2, -10, 7, -18,
    -- layer=1 filter=101 channel=61
    -5, 10, -6, -9, 4, -2, 0, -1, -4,
    -- layer=1 filter=101 channel=62
    -3, -21, -32, -21, 3, -26, -61, -23, 58,
    -- layer=1 filter=101 channel=63
    -28, -20, -25, -2, -58, 2, -26, -47, -39,
    -- layer=1 filter=101 channel=64
    -4, -26, -11, 3, -29, -11, 8, -13, -3,
    -- layer=1 filter=101 channel=65
    -5, -6, -6, 1, -7, -8, -8, 6, -31,
    -- layer=1 filter=101 channel=66
    -14, -35, -16, -21, -31, 3, -36, -5, -24,
    -- layer=1 filter=101 channel=67
    10, -2, 39, 24, -18, 18, 23, 7, -9,
    -- layer=1 filter=101 channel=68
    -31, 45, -28, -16, 14, 11, -27, -21, 25,
    -- layer=1 filter=101 channel=69
    -2, 31, -19, -32, 19, 21, -60, -29, 79,
    -- layer=1 filter=101 channel=70
    -18, 0, 13, -5, -6, 49, -7, -19, -17,
    -- layer=1 filter=101 channel=71
    7, -28, 22, 4, 14, 7, -11, 4, 5,
    -- layer=1 filter=101 channel=72
    -2, -20, -30, -10, 3, -6, -13, -47, -33,
    -- layer=1 filter=101 channel=73
    7, -12, 6, -11, -4, 3, -9, 4, 1,
    -- layer=1 filter=101 channel=74
    -58, -5, -48, 6, -3, -16, -7, -24, -42,
    -- layer=1 filter=101 channel=75
    -8, -60, 4, 5, -35, -9, 0, -8, -25,
    -- layer=1 filter=101 channel=76
    -44, 16, -29, 9, 10, -21, 0, -8, -6,
    -- layer=1 filter=101 channel=77
    24, 12, 2, 11, 31, -2, 8, 37, 4,
    -- layer=1 filter=101 channel=78
    -6, 0, 0, -8, -5, 5, -10, -2, -3,
    -- layer=1 filter=101 channel=79
    -7, -13, -34, -28, -6, -4, -57, -20, 53,
    -- layer=1 filter=101 channel=80
    0, -1, -9, -7, -3, 6, 5, 8, -1,
    -- layer=1 filter=101 channel=81
    2, 6, -1, 1, 2, -17, 9, 14, 28,
    -- layer=1 filter=101 channel=82
    7, 9, 0, 2, -3, -21, 12, 8, 0,
    -- layer=1 filter=101 channel=83
    11, 17, -46, -12, 22, -17, -9, 7, 54,
    -- layer=1 filter=101 channel=84
    -46, 10, -24, -1, -20, -23, -10, -56, -49,
    -- layer=1 filter=101 channel=85
    17, -5, 0, 5, -24, 7, 35, -21, 33,
    -- layer=1 filter=101 channel=86
    -22, -25, -12, -21, -20, -5, -28, 0, -14,
    -- layer=1 filter=101 channel=87
    -38, -42, -8, -9, 0, 10, -2, -29, -53,
    -- layer=1 filter=101 channel=88
    -22, 8, 44, -24, 10, 6, 10, 12, -9,
    -- layer=1 filter=101 channel=89
    6, 11, -23, 4, -12, 0, -7, -14, -5,
    -- layer=1 filter=101 channel=90
    -8, 25, -32, -17, 37, 8, -18, -21, 24,
    -- layer=1 filter=101 channel=91
    5, -11, 0, -3, -20, -15, 21, -3, -24,
    -- layer=1 filter=101 channel=92
    -35, 51, -14, 0, 26, 20, 1, -32, 32,
    -- layer=1 filter=101 channel=93
    11, -2, -12, 3, -9, -20, -7, -5, 13,
    -- layer=1 filter=101 channel=94
    -15, -21, -9, -17, -28, 5, -24, 6, -29,
    -- layer=1 filter=101 channel=95
    -36, -15, -36, 6, -32, -17, -3, -66, -40,
    -- layer=1 filter=101 channel=96
    -17, -3, 12, -8, -15, 0, -2, -11, -19,
    -- layer=1 filter=101 channel=97
    -1, -10, -8, -15, -8, -41, -23, -3, -6,
    -- layer=1 filter=101 channel=98
    14, -6, -38, -26, -5, -42, -50, -17, 48,
    -- layer=1 filter=101 channel=99
    -25, -4, -9, -2, 5, -4, 0, 16, -1,
    -- layer=1 filter=101 channel=100
    -39, 8, -28, -1, -25, 12, -16, -35, -33,
    -- layer=1 filter=101 channel=101
    -9, 6, -6, 4, -7, 1, 5, -19, -19,
    -- layer=1 filter=101 channel=102
    -24, -38, -34, -7, -26, -14, -15, -12, -49,
    -- layer=1 filter=101 channel=103
    -28, 15, -22, -17, 2, -8, -21, -36, -30,
    -- layer=1 filter=101 channel=104
    15, -12, -3, 2, -32, 20, 11, -35, 27,
    -- layer=1 filter=101 channel=105
    -3, -27, 0, -7, -32, -25, -9, 6, -26,
    -- layer=1 filter=101 channel=106
    -1, 33, -24, -1, 2, 10, -7, -25, 9,
    -- layer=1 filter=101 channel=107
    5, 7, 8, -9, -5, -4, -3, 1, -1,
    -- layer=1 filter=101 channel=108
    -13, 54, -28, -28, 34, 25, -33, -27, 48,
    -- layer=1 filter=101 channel=109
    -8, 0, -9, -9, 7, 2, 7, -7, -1,
    -- layer=1 filter=101 channel=110
    0, -8, -2, 0, -5, -6, 1, 0, -11,
    -- layer=1 filter=101 channel=111
    -24, -21, -43, 10, -37, 0, 5, -23, -40,
    -- layer=1 filter=101 channel=112
    4, 5, -28, 0, -50, 5, 5, -24, -17,
    -- layer=1 filter=101 channel=113
    -21, -13, 33, 12, -24, 26, 6, -15, 4,
    -- layer=1 filter=101 channel=114
    -28, 4, -20, -53, -21, 18, -68, -28, 36,
    -- layer=1 filter=101 channel=115
    -11, -13, -9, -14, -19, -16, 5, 1, -11,
    -- layer=1 filter=101 channel=116
    -9, 2, 1, 7, -7, 9, 2, -5, 0,
    -- layer=1 filter=101 channel=117
    -24, -17, -2, 12, -29, -24, 23, -18, -33,
    -- layer=1 filter=101 channel=118
    -52, 4, -30, 14, -12, -19, -9, -50, -51,
    -- layer=1 filter=101 channel=119
    -20, 32, -15, -17, 37, 6, -16, -31, 36,
    -- layer=1 filter=101 channel=120
    -12, -5, 12, 16, -27, -13, 10, -4, -17,
    -- layer=1 filter=101 channel=121
    -47, -76, 17, 18, 13, 12, -11, -6, -48,
    -- layer=1 filter=101 channel=122
    -4, 9, -9, 10, 6, -8, 10, 4, -6,
    -- layer=1 filter=101 channel=123
    -27, -36, 3, -17, -5, 16, -12, -10, -38,
    -- layer=1 filter=101 channel=124
    -11, -5, 11, -3, -1, 2, -9, 1, -5,
    -- layer=1 filter=101 channel=125
    -39, -26, 23, 5, -32, 37, 37, -30, -25,
    -- layer=1 filter=101 channel=126
    20, 2, -31, -14, 3, -54, -58, -12, 58,
    -- layer=1 filter=101 channel=127
    -31, -10, -14, 15, -35, 1, -3, -31, -39,
    -- layer=1 filter=102 channel=0
    -3, 10, -1, -12, 0, 3, 10, 12, 16,
    -- layer=1 filter=102 channel=1
    -7, -17, -8, -5, -5, -8, -8, 8, 18,
    -- layer=1 filter=102 channel=2
    2, 3, 3, 2, -14, -4, 1, -1, -23,
    -- layer=1 filter=102 channel=3
    4, -2, -9, 9, -6, 8, -4, -11, -3,
    -- layer=1 filter=102 channel=4
    -8, 0, 3, 6, 0, 0, -8, 1, -6,
    -- layer=1 filter=102 channel=5
    -16, -17, -20, -29, -33, -32, -11, -3, 15,
    -- layer=1 filter=102 channel=6
    -41, -41, -30, -46, -45, -36, -15, -25, -44,
    -- layer=1 filter=102 channel=7
    -24, -45, -23, -33, -60, -27, -14, 8, -43,
    -- layer=1 filter=102 channel=8
    -25, -29, 0, -14, -50, -39, -9, 8, 21,
    -- layer=1 filter=102 channel=9
    -7, -5, -7, -17, -16, -5, -33, -17, -14,
    -- layer=1 filter=102 channel=10
    1, -31, -10, -25, -52, -23, 17, 24, -15,
    -- layer=1 filter=102 channel=11
    -11, 2, 0, -12, 5, -2, 1, -9, 1,
    -- layer=1 filter=102 channel=12
    21, 17, -17, -21, -6, -16, -1, -11, -14,
    -- layer=1 filter=102 channel=13
    -2, 12, 20, 7, 8, -2, 11, 3, 6,
    -- layer=1 filter=102 channel=14
    -56, -31, -4, -26, -39, -39, -8, -32, -52,
    -- layer=1 filter=102 channel=15
    -39, -66, -26, -63, -43, -41, -28, -48, -11,
    -- layer=1 filter=102 channel=16
    -37, -50, -34, -9, -40, -37, -5, 10, 19,
    -- layer=1 filter=102 channel=17
    1, 0, 1, -7, 0, 9, -5, 5, 13,
    -- layer=1 filter=102 channel=18
    -16, -31, -16, -49, -28, -24, 6, -19, -52,
    -- layer=1 filter=102 channel=19
    -30, -39, -46, -50, -30, -41, -12, -43, -26,
    -- layer=1 filter=102 channel=20
    25, 15, 12, 13, 18, 20, 21, 9, 10,
    -- layer=1 filter=102 channel=21
    -10, -8, 0, -13, -7, 0, -14, -8, -24,
    -- layer=1 filter=102 channel=22
    0, 10, 12, 0, -13, -1, 4, 0, 20,
    -- layer=1 filter=102 channel=23
    -11, -5, -13, -2, -1, 0, 14, -10, 1,
    -- layer=1 filter=102 channel=24
    7, 0, 0, -12, 5, 9, 0, 1, 0,
    -- layer=1 filter=102 channel=25
    -4, -31, -9, -25, -36, -19, -18, 0, -5,
    -- layer=1 filter=102 channel=26
    -3, -16, 12, -2, -8, 11, 12, -14, 13,
    -- layer=1 filter=102 channel=27
    -27, -31, -30, -33, -26, -37, -28, -16, -37,
    -- layer=1 filter=102 channel=28
    -19, -18, -14, 7, -13, 1, -1, 13, -16,
    -- layer=1 filter=102 channel=29
    -27, -26, -31, -18, -9, -14, -24, -20, -28,
    -- layer=1 filter=102 channel=30
    -63, -62, -80, -58, -71, -49, -16, -56, -118,
    -- layer=1 filter=102 channel=31
    -22, -25, -31, -26, -36, -49, -3, -36, -41,
    -- layer=1 filter=102 channel=32
    -40, -78, -15, -37, -57, -30, -20, -51, -25,
    -- layer=1 filter=102 channel=33
    -3, -11, 4, -3, 2, -1, -6, -1, -1,
    -- layer=1 filter=102 channel=34
    -6, -34, -24, -14, -24, -32, -4, -18, -38,
    -- layer=1 filter=102 channel=35
    -13, -14, -2, -17, -5, -19, -15, -7, -8,
    -- layer=1 filter=102 channel=36
    4, 16, 21, 10, 9, 18, 20, 21, 17,
    -- layer=1 filter=102 channel=37
    -9, -28, -20, -7, -31, -28, 3, -3, 30,
    -- layer=1 filter=102 channel=38
    12, 13, 7, 4, 14, 4, 1, 5, 5,
    -- layer=1 filter=102 channel=39
    -5, -3, -3, 0, -10, -9, 1, 4, -7,
    -- layer=1 filter=102 channel=40
    -54, -36, -20, -19, -51, -30, 18, -15, -31,
    -- layer=1 filter=102 channel=41
    0, -7, -4, -6, -47, -2, -21, -35, -43,
    -- layer=1 filter=102 channel=42
    -2, -14, -27, -5, 0, -8, 5, -27, -22,
    -- layer=1 filter=102 channel=43
    -5, -20, 3, -25, -21, -27, -8, 5, 24,
    -- layer=1 filter=102 channel=44
    -16, -77, -16, -29, -48, -42, -1, -59, -27,
    -- layer=1 filter=102 channel=45
    -16, -27, -11, -15, -14, 0, -7, -18, -5,
    -- layer=1 filter=102 channel=46
    -27, -15, 11, -42, -26, -47, -23, -39, -26,
    -- layer=1 filter=102 channel=47
    -20, 5, -14, -3, -17, 12, -2, 13, -12,
    -- layer=1 filter=102 channel=48
    -5, -6, -13, -14, -5, 1, 1, 3, -14,
    -- layer=1 filter=102 channel=49
    0, -10, 2, -21, -12, -13, -9, -15, -28,
    -- layer=1 filter=102 channel=50
    0, 2, -5, 1, -9, 8, -5, 4, 0,
    -- layer=1 filter=102 channel=51
    -14, -8, -9, -16, -10, -12, 5, -7, -18,
    -- layer=1 filter=102 channel=52
    -6, -3, 6, -3, -4, 7, 3, 4, -3,
    -- layer=1 filter=102 channel=53
    1, -7, -12, -5, 0, -13, -12, -14, -8,
    -- layer=1 filter=102 channel=54
    14, -26, -8, -38, -36, -8, 9, -6, 4,
    -- layer=1 filter=102 channel=55
    3, 6, 0, 12, 0, 0, 16, 0, 1,
    -- layer=1 filter=102 channel=56
    -11, -3, -10, -4, -8, 8, 9, -6, 5,
    -- layer=1 filter=102 channel=57
    -5, -35, 2, -13, -40, 9, 20, 16, 0,
    -- layer=1 filter=102 channel=58
    -36, -48, -54, -32, -72, -48, 5, 26, -35,
    -- layer=1 filter=102 channel=59
    0, -5, -5, 2, -9, -12, 4, -7, 6,
    -- layer=1 filter=102 channel=60
    -12, -9, 4, -3, -8, -16, 0, -10, -6,
    -- layer=1 filter=102 channel=61
    -2, -11, -4, 10, 6, 7, -10, -2, 6,
    -- layer=1 filter=102 channel=62
    -46, -63, -23, -44, -60, -31, -6, -10, 12,
    -- layer=1 filter=102 channel=63
    0, -14, -1, -3, -3, -10, -15, -4, -11,
    -- layer=1 filter=102 channel=64
    2, 8, 4, 9, -3, 2, 2, 9, 5,
    -- layer=1 filter=102 channel=65
    -10, -5, -3, -2, -20, -1, -14, -6, -25,
    -- layer=1 filter=102 channel=66
    0, 1, 4, -7, 10, 2, 0, 5, 16,
    -- layer=1 filter=102 channel=67
    23, -4, 0, -15, -3, -8, -4, -18, -23,
    -- layer=1 filter=102 channel=68
    -32, -90, -33, -20, -90, -67, -34, -79, -29,
    -- layer=1 filter=102 channel=69
    -17, -21, -1, -24, -26, -35, -9, 0, 11,
    -- layer=1 filter=102 channel=70
    12, -10, 11, -31, -55, -49, -8, -15, -43,
    -- layer=1 filter=102 channel=71
    -6, -1, -2, 16, -3, -4, -4, 2, 10,
    -- layer=1 filter=102 channel=72
    -14, 4, -8, -6, -6, -5, -23, -27, -36,
    -- layer=1 filter=102 channel=73
    -9, 10, 9, 9, -3, 2, 0, 11, 7,
    -- layer=1 filter=102 channel=74
    -8, -15, -9, -12, -40, -33, -8, -28, -19,
    -- layer=1 filter=102 channel=75
    -77, -31, -7, -34, -24, -19, 12, -35, -46,
    -- layer=1 filter=102 channel=76
    -12, -23, -12, -1, -5, -2, -10, -12, -28,
    -- layer=1 filter=102 channel=77
    -15, -12, -8, -3, -5, -11, -7, -8, -5,
    -- layer=1 filter=102 channel=78
    -1, 4, 0, -4, 1, -2, 12, 8, 0,
    -- layer=1 filter=102 channel=79
    -10, -30, -1, -18, -25, -19, 22, 3, 29,
    -- layer=1 filter=102 channel=80
    1, 0, 6, 7, -7, -6, -5, 0, -2,
    -- layer=1 filter=102 channel=81
    -9, -19, -14, -10, -7, -7, -12, 12, 7,
    -- layer=1 filter=102 channel=82
    4, 1, 0, 2, -12, -3, -3, -20, -16,
    -- layer=1 filter=102 channel=83
    -21, -14, -10, -10, -14, -13, -1, -11, 20,
    -- layer=1 filter=102 channel=84
    -63, -76, -42, -60, -64, -52, -30, -52, -58,
    -- layer=1 filter=102 channel=85
    -7, -2, -21, -25, -40, 8, 16, -11, -3,
    -- layer=1 filter=102 channel=86
    4, 14, 3, 17, 19, 5, 11, 10, 14,
    -- layer=1 filter=102 channel=87
    -16, -58, -33, -39, -38, -22, -51, -85, -55,
    -- layer=1 filter=102 channel=88
    -8, -4, 0, -13, -2, -3, -4, -24, -28,
    -- layer=1 filter=102 channel=89
    -14, -21, -6, -16, -11, -6, -18, -33, -19,
    -- layer=1 filter=102 channel=90
    -23, -83, -31, -19, -64, -30, 4, -42, -20,
    -- layer=1 filter=102 channel=91
    10, 23, 22, 19, 17, 15, 16, 10, 12,
    -- layer=1 filter=102 channel=92
    -25, -25, 9, -21, -8, -1, 0, -18, 14,
    -- layer=1 filter=102 channel=93
    9, 13, 20, 6, 0, 7, 2, 1, 22,
    -- layer=1 filter=102 channel=94
    -1, 9, -4, 4, 0, -1, -4, 12, 0,
    -- layer=1 filter=102 channel=95
    -66, -78, -44, -48, -59, -52, -50, -84, -76,
    -- layer=1 filter=102 channel=96
    -2, -10, 4, 3, -4, -9, 6, 7, 6,
    -- layer=1 filter=102 channel=97
    5, 17, 19, 11, 4, 20, 15, 19, 23,
    -- layer=1 filter=102 channel=98
    13, -1, 33, 4, -10, -2, 0, 4, 30,
    -- layer=1 filter=102 channel=99
    -34, -50, -44, -36, -42, -30, 0, 12, -49,
    -- layer=1 filter=102 channel=100
    -7, -16, -14, -14, -12, -3, -11, -5, -2,
    -- layer=1 filter=102 channel=101
    16, 14, 2, 0, 1, 16, 14, 6, 0,
    -- layer=1 filter=102 channel=102
    2, -7, 2, -4, 6, 4, -1, 0, -5,
    -- layer=1 filter=102 channel=103
    -6, -12, -6, -8, -21, -15, -1, -25, -6,
    -- layer=1 filter=102 channel=104
    -2, 9, 2, 12, 0, 13, 2, 12, -5,
    -- layer=1 filter=102 channel=105
    -1, 11, 14, 9, 14, 8, 5, 13, 22,
    -- layer=1 filter=102 channel=106
    0, -2, 18, -3, 7, 4, 9, -15, 0,
    -- layer=1 filter=102 channel=107
    3, 13, 5, -2, 16, 16, -1, 0, 1,
    -- layer=1 filter=102 channel=108
    -47, -103, -22, -44, -61, -37, -19, -76, -45,
    -- layer=1 filter=102 channel=109
    6, 8, -8, 5, -6, -7, 5, -2, -8,
    -- layer=1 filter=102 channel=110
    -3, 11, -1, 1, 10, -8, -2, 2, 6,
    -- layer=1 filter=102 channel=111
    -42, -55, -20, -33, -50, -27, 3, -16, -65,
    -- layer=1 filter=102 channel=112
    -11, -12, -3, -9, -6, -7, 22, -10, -19,
    -- layer=1 filter=102 channel=113
    -25, -50, -32, -20, -31, -36, -15, -45, -28,
    -- layer=1 filter=102 channel=114
    -40, -49, -63, -12, -41, -39, -21, 4, 4,
    -- layer=1 filter=102 channel=115
    2, 15, 11, 4, 21, 23, 23, 24, 33,
    -- layer=1 filter=102 channel=116
    7, 0, 1, 0, 0, -1, 0, 0, 9,
    -- layer=1 filter=102 channel=117
    -68, -84, 0, -60, -53, -80, 23, -18, -64,
    -- layer=1 filter=102 channel=118
    -16, -85, -44, -43, -35, -36, 0, -43, -48,
    -- layer=1 filter=102 channel=119
    -54, -94, -37, -50, -78, -44, -31, -75, -48,
    -- layer=1 filter=102 channel=120
    2, 4, -5, -6, -12, -5, -5, 12, -11,
    -- layer=1 filter=102 channel=121
    -16, -18, -5, 1, -13, -12, -20, -18, -27,
    -- layer=1 filter=102 channel=122
    0, -8, -8, -1, 8, -1, -2, 5, -10,
    -- layer=1 filter=102 channel=123
    -15, -11, -5, -16, -1, -4, -8, -11, -20,
    -- layer=1 filter=102 channel=124
    -5, -1, 3, -2, -4, -9, -1, -4, -6,
    -- layer=1 filter=102 channel=125
    11, -6, -1, -37, -55, -41, 5, -24, -34,
    -- layer=1 filter=102 channel=126
    -28, -13, 8, -33, -54, -58, -45, -18, -7,
    -- layer=1 filter=102 channel=127
    -69, -81, -37, -64, -59, -66, -11, -68, -81,
    -- layer=1 filter=103 channel=0
    -11, -3, -6, 9, 4, 3, -11, -7, -3,
    -- layer=1 filter=103 channel=1
    -5, -10, -11, 8, -1, 0, 2, -7, 0,
    -- layer=1 filter=103 channel=2
    7, -5, 3, -11, -12, -13, -7, -9, 10,
    -- layer=1 filter=103 channel=3
    -7, 7, -10, 1, -1, -4, 7, 11, 2,
    -- layer=1 filter=103 channel=4
    -11, 6, -10, -2, 0, -8, -11, -8, 6,
    -- layer=1 filter=103 channel=5
    7, -9, 0, -1, -5, 8, -6, -3, -8,
    -- layer=1 filter=103 channel=6
    -8, -11, 0, 4, -18, -10, 4, 1, -4,
    -- layer=1 filter=103 channel=7
    -15, 7, 2, 12, 1, -10, 4, -3, -27,
    -- layer=1 filter=103 channel=8
    -8, -9, -6, -9, 0, -1, 0, 1, -10,
    -- layer=1 filter=103 channel=9
    3, -8, 3, 3, 6, -12, 1, 5, 19,
    -- layer=1 filter=103 channel=10
    -2, 3, -10, 7, -1, -6, 0, 10, -17,
    -- layer=1 filter=103 channel=11
    0, -21, -8, -5, -1, 0, -2, 2, 2,
    -- layer=1 filter=103 channel=12
    -5, -2, -2, -2, 6, -1, 14, -1, -3,
    -- layer=1 filter=103 channel=13
    -10, 0, -12, 0, -1, -2, -5, -3, -15,
    -- layer=1 filter=103 channel=14
    -10, -6, 8, 7, -5, -3, 5, -11, 5,
    -- layer=1 filter=103 channel=15
    6, -8, 6, -11, 3, -9, -9, -7, -8,
    -- layer=1 filter=103 channel=16
    -1, 4, -3, -6, -2, -8, -2, -4, -5,
    -- layer=1 filter=103 channel=17
    4, 6, -12, -5, -9, -11, 0, -2, 2,
    -- layer=1 filter=103 channel=18
    -5, -2, -13, -6, -7, 2, 11, 5, -1,
    -- layer=1 filter=103 channel=19
    4, -8, 8, 0, 4, 6, 0, -4, 2,
    -- layer=1 filter=103 channel=20
    -12, -12, -9, 1, -9, -17, 0, -3, -12,
    -- layer=1 filter=103 channel=21
    -4, -2, -4, 6, -9, 3, -2, -10, -7,
    -- layer=1 filter=103 channel=22
    -11, -13, 0, -1, 0, -7, -13, -15, -11,
    -- layer=1 filter=103 channel=23
    -2, 0, -13, 8, -11, -10, -1, 7, 7,
    -- layer=1 filter=103 channel=24
    2, 6, 3, -14, 3, -20, -15, -14, -13,
    -- layer=1 filter=103 channel=25
    -12, -1, 6, 3, 3, 2, -4, 5, -12,
    -- layer=1 filter=103 channel=26
    -1, -3, 5, -5, -18, 1, -11, 2, -7,
    -- layer=1 filter=103 channel=27
    -8, -7, 7, -5, -9, -3, -2, -8, 9,
    -- layer=1 filter=103 channel=28
    -4, 6, 2, 7, -2, 5, 9, -12, 0,
    -- layer=1 filter=103 channel=29
    -8, 9, -5, 5, -9, 2, -1, -9, 1,
    -- layer=1 filter=103 channel=30
    5, 8, 0, -2, -6, -5, -1, -8, 0,
    -- layer=1 filter=103 channel=31
    8, 4, -4, -9, 2, -1, 2, -6, 1,
    -- layer=1 filter=103 channel=32
    1, -5, -10, -6, 2, -9, -9, 6, 0,
    -- layer=1 filter=103 channel=33
    -8, -9, 0, 2, 3, -7, 9, 5, -7,
    -- layer=1 filter=103 channel=34
    4, -5, 8, 6, -1, 5, 2, -9, -8,
    -- layer=1 filter=103 channel=35
    -5, -7, 4, 1, -6, 7, -7, -7, -6,
    -- layer=1 filter=103 channel=36
    -13, 1, -14, -10, 2, 7, 7, -3, 0,
    -- layer=1 filter=103 channel=37
    12, 3, -5, -8, -12, 7, -1, -6, -14,
    -- layer=1 filter=103 channel=38
    9, 1, -13, -1, -16, 0, -7, -5, -4,
    -- layer=1 filter=103 channel=39
    3, -2, 1, -4, -7, -12, -9, 4, -2,
    -- layer=1 filter=103 channel=40
    -4, -9, -12, 9, -14, -20, 3, 0, -16,
    -- layer=1 filter=103 channel=41
    -8, -6, -7, -9, -10, 1, -6, 1, 0,
    -- layer=1 filter=103 channel=42
    9, 1, -7, -1, -1, -11, 8, -6, 1,
    -- layer=1 filter=103 channel=43
    -6, 6, -2, 0, 2, 8, -9, -5, 2,
    -- layer=1 filter=103 channel=44
    3, 3, -12, -1, -1, 7, 8, -5, 2,
    -- layer=1 filter=103 channel=45
    3, -7, -8, 7, 4, -3, 5, -3, 1,
    -- layer=1 filter=103 channel=46
    4, 0, 8, -14, -7, -14, -5, 1, 0,
    -- layer=1 filter=103 channel=47
    -4, -8, 0, -2, -1, 0, -8, -8, 0,
    -- layer=1 filter=103 channel=48
    5, 3, -6, 8, -4, -11, 0, 5, -3,
    -- layer=1 filter=103 channel=49
    8, -8, 7, -9, -2, 7, 2, 4, -4,
    -- layer=1 filter=103 channel=50
    -9, 4, 0, 2, -1, 6, 5, -9, -7,
    -- layer=1 filter=103 channel=51
    6, -13, 7, -8, -10, 4, 0, -3, -5,
    -- layer=1 filter=103 channel=52
    2, 8, 1, -3, -2, 10, 10, -5, -9,
    -- layer=1 filter=103 channel=53
    0, 0, -10, 9, -7, 0, -6, -11, 8,
    -- layer=1 filter=103 channel=54
    -8, 4, 5, -15, -7, 5, -1, 6, -3,
    -- layer=1 filter=103 channel=55
    -12, -5, -8, -7, -13, -5, -14, -13, -12,
    -- layer=1 filter=103 channel=56
    0, -2, 0, 5, 4, -6, -6, -8, -9,
    -- layer=1 filter=103 channel=57
    1, -4, 0, 3, -8, 4, 5, -12, -9,
    -- layer=1 filter=103 channel=58
    -12, 1, 5, 3, 11, -11, -13, 15, -2,
    -- layer=1 filter=103 channel=59
    7, -8, -8, 0, 7, -2, -10, 5, 3,
    -- layer=1 filter=103 channel=60
    -7, 0, -6, -5, -7, -3, 10, 6, -6,
    -- layer=1 filter=103 channel=61
    -9, 9, 5, 8, -4, 1, 4, 7, -8,
    -- layer=1 filter=103 channel=62
    -6, 6, 4, 4, -6, -3, -2, -12, -4,
    -- layer=1 filter=103 channel=63
    -15, 3, 0, -12, -10, -5, -12, -3, -5,
    -- layer=1 filter=103 channel=64
    0, -8, -10, -7, -11, -11, -2, -4, -10,
    -- layer=1 filter=103 channel=65
    6, 7, 4, 2, 4, -6, -5, -1, -11,
    -- layer=1 filter=103 channel=66
    1, -7, -6, -11, 0, -12, 7, -6, 6,
    -- layer=1 filter=103 channel=67
    8, 3, 5, 8, 12, -10, 0, 5, -2,
    -- layer=1 filter=103 channel=68
    -9, 3, -10, -12, 3, 5, -11, -9, -6,
    -- layer=1 filter=103 channel=69
    -7, 5, -16, 9, 1, -1, -9, -10, -10,
    -- layer=1 filter=103 channel=70
    -10, 3, 13, 1, 0, 6, 1, 5, -11,
    -- layer=1 filter=103 channel=71
    8, -9, -13, -9, -16, -4, -4, -13, 0,
    -- layer=1 filter=103 channel=72
    7, 0, 5, -7, -5, 3, -4, 2, -3,
    -- layer=1 filter=103 channel=73
    -8, -4, -10, 2, 0, 1, -3, -10, 8,
    -- layer=1 filter=103 channel=74
    3, 7, -7, 7, -6, 5, -1, -6, -11,
    -- layer=1 filter=103 channel=75
    9, 2, 11, -5, 0, 0, 12, 7, 14,
    -- layer=1 filter=103 channel=76
    -2, 7, -4, 6, -8, -4, -4, -7, -10,
    -- layer=1 filter=103 channel=77
    6, 2, -7, 4, 3, -7, 6, -1, -3,
    -- layer=1 filter=103 channel=78
    -11, 8, -7, -5, 3, 2, -6, -4, 0,
    -- layer=1 filter=103 channel=79
    2, 7, -12, -1, 2, -3, -15, -11, -14,
    -- layer=1 filter=103 channel=80
    3, 0, 0, -12, -7, 4, -11, 7, -9,
    -- layer=1 filter=103 channel=81
    -11, -5, -8, 2, -12, -14, -10, -13, 0,
    -- layer=1 filter=103 channel=82
    -4, -5, -5, -6, 2, -11, 4, -9, -13,
    -- layer=1 filter=103 channel=83
    2, -2, 0, -6, -2, -1, 5, -2, 7,
    -- layer=1 filter=103 channel=84
    -16, -16, 2, 5, -10, 9, -7, -8, -4,
    -- layer=1 filter=103 channel=85
    -1, 4, -7, 8, 7, -5, -6, 3, -7,
    -- layer=1 filter=103 channel=86
    -9, -13, -13, -8, 3, -11, -8, 0, -5,
    -- layer=1 filter=103 channel=87
    7, -6, 0, 6, -1, 4, 4, -8, -8,
    -- layer=1 filter=103 channel=88
    3, 1, 5, 4, 7, 2, -9, -5, 7,
    -- layer=1 filter=103 channel=89
    2, 2, 4, -10, -6, 4, -2, -6, -6,
    -- layer=1 filter=103 channel=90
    4, -4, -3, -9, -10, -3, -6, -11, -12,
    -- layer=1 filter=103 channel=91
    -1, -1, -15, -9, 3, -7, 5, -2, 1,
    -- layer=1 filter=103 channel=92
    3, -7, -7, 8, 8, 6, 9, 8, 0,
    -- layer=1 filter=103 channel=93
    1, 7, 1, -6, -12, -9, -11, -10, -2,
    -- layer=1 filter=103 channel=94
    5, 0, 5, -3, 3, 3, 6, 1, 0,
    -- layer=1 filter=103 channel=95
    -9, -6, -7, -12, -4, 3, 4, -5, -10,
    -- layer=1 filter=103 channel=96
    -2, -2, -11, -8, -6, -4, 9, 7, -10,
    -- layer=1 filter=103 channel=97
    -1, -2, -12, -3, -6, 1, 6, -5, -10,
    -- layer=1 filter=103 channel=98
    -6, -8, -12, -6, -11, 6, -10, 1, 1,
    -- layer=1 filter=103 channel=99
    -11, -1, -5, 9, -2, 2, -3, -10, 4,
    -- layer=1 filter=103 channel=100
    -10, 1, -4, -3, -2, 2, 1, -5, -1,
    -- layer=1 filter=103 channel=101
    -8, 3, -13, 2, -4, 5, -9, -1, 4,
    -- layer=1 filter=103 channel=102
    -7, 8, -6, 0, -4, -6, -10, -5, -1,
    -- layer=1 filter=103 channel=103
    0, -20, -6, 1, 3, -2, 8, -4, -2,
    -- layer=1 filter=103 channel=104
    2, 7, 6, 8, -11, -8, 8, 0, 8,
    -- layer=1 filter=103 channel=105
    -8, 0, 0, 6, -4, 4, 4, -10, -5,
    -- layer=1 filter=103 channel=106
    0, -16, -12, -16, -2, -4, 5, -10, 2,
    -- layer=1 filter=103 channel=107
    5, 5, 6, -7, 8, 1, -8, -7, -3,
    -- layer=1 filter=103 channel=108
    -21, -10, 3, -9, -7, -9, -21, -2, 8,
    -- layer=1 filter=103 channel=109
    0, 5, 7, 7, -4, 4, 1, 1, -8,
    -- layer=1 filter=103 channel=110
    -4, -6, 6, 5, -5, 0, -9, -8, 0,
    -- layer=1 filter=103 channel=111
    -4, 3, 8, -1, -2, -3, -2, 0, -3,
    -- layer=1 filter=103 channel=112
    4, -9, -6, -5, 8, -7, -5, -4, 0,
    -- layer=1 filter=103 channel=113
    5, -6, -4, 0, -10, -6, -4, -2, -6,
    -- layer=1 filter=103 channel=114
    7, -7, 9, -1, 7, 10, 0, -9, 0,
    -- layer=1 filter=103 channel=115
    -6, 5, 4, 0, -6, -10, -5, -4, -11,
    -- layer=1 filter=103 channel=116
    11, -3, -9, -5, 10, 4, -8, -2, 0,
    -- layer=1 filter=103 channel=117
    -19, 0, -1, -4, -11, -1, 11, -3, -13,
    -- layer=1 filter=103 channel=118
    -2, -3, -8, 0, -9, 7, 8, 7, 0,
    -- layer=1 filter=103 channel=119
    -20, -3, -13, -10, 5, 2, -19, 0, -3,
    -- layer=1 filter=103 channel=120
    1, -10, -4, -1, -4, -9, -10, -5, -2,
    -- layer=1 filter=103 channel=121
    5, -6, 8, -22, -6, -11, 0, -9, 8,
    -- layer=1 filter=103 channel=122
    0, -7, -1, 9, 0, -9, -5, 5, 2,
    -- layer=1 filter=103 channel=123
    -2, -3, -6, -13, 0, 5, 7, -2, 7,
    -- layer=1 filter=103 channel=124
    7, -4, 1, 1, 7, -4, -10, -4, 0,
    -- layer=1 filter=103 channel=125
    -9, -11, 4, -3, -4, 13, 8, 7, -25,
    -- layer=1 filter=103 channel=126
    -11, -3, -2, -1, -9, -10, 7, 7, 4,
    -- layer=1 filter=103 channel=127
    -6, 4, -2, -11, 3, 0, 16, 10, 3,
    -- layer=1 filter=104 channel=0
    -4, -1, 1, -1, 0, -3, -10, 3, -6,
    -- layer=1 filter=104 channel=1
    0, -5, 2, 2, -5, -7, 2, 8, 8,
    -- layer=1 filter=104 channel=2
    1, 9, 0, -9, -4, -9, -11, -6, 2,
    -- layer=1 filter=104 channel=3
    -5, -5, 1, 1, 7, -3, -2, 2, -9,
    -- layer=1 filter=104 channel=4
    2, 2, -10, -10, -6, 0, 4, 4, 7,
    -- layer=1 filter=104 channel=5
    -1, 5, 0, 3, 2, -5, -7, -4, -3,
    -- layer=1 filter=104 channel=6
    -10, 0, 7, -10, -8, 1, -7, -11, -9,
    -- layer=1 filter=104 channel=7
    1, 1, -7, 4, 5, -3, 3, -3, -12,
    -- layer=1 filter=104 channel=8
    9, -9, -5, -7, -9, -4, -8, -1, -8,
    -- layer=1 filter=104 channel=9
    -2, 3, -6, 4, 5, -1, 6, 8, 6,
    -- layer=1 filter=104 channel=10
    -12, -14, -1, -12, -9, -7, -5, -14, -1,
    -- layer=1 filter=104 channel=11
    -4, -13, -3, 1, -6, -7, 0, -7, -1,
    -- layer=1 filter=104 channel=12
    4, -6, 7, 5, 0, -9, -8, -6, 6,
    -- layer=1 filter=104 channel=13
    -12, -10, -8, -11, -1, 5, -3, 1, -10,
    -- layer=1 filter=104 channel=14
    -3, -2, 9, -7, 7, -3, 0, -9, 0,
    -- layer=1 filter=104 channel=15
    -3, 1, -4, 0, -7, 5, -7, -3, 0,
    -- layer=1 filter=104 channel=16
    -9, 4, -5, 7, -7, -9, 4, 6, -4,
    -- layer=1 filter=104 channel=17
    -7, -7, -8, -7, -6, 5, 0, 3, 4,
    -- layer=1 filter=104 channel=18
    1, -10, -10, -10, 9, -3, 1, 11, -6,
    -- layer=1 filter=104 channel=19
    1, -2, 8, 2, 0, 3, 7, -5, 6,
    -- layer=1 filter=104 channel=20
    -7, -3, -10, -11, -6, -4, -1, 7, -7,
    -- layer=1 filter=104 channel=21
    -10, 7, -3, -1, 2, -10, -3, -2, 1,
    -- layer=1 filter=104 channel=22
    7, 0, 5, -10, -5, -2, -4, -6, 1,
    -- layer=1 filter=104 channel=23
    -1, 9, -4, -6, 6, 8, 0, -3, 4,
    -- layer=1 filter=104 channel=24
    -11, 7, 0, -11, 0, 3, 5, 1, 1,
    -- layer=1 filter=104 channel=25
    -1, -6, -3, -9, 9, -5, -6, 6, -9,
    -- layer=1 filter=104 channel=26
    5, -1, -6, 2, 0, -8, -1, -8, 2,
    -- layer=1 filter=104 channel=27
    -12, -10, -2, 0, -2, -2, 3, -7, -9,
    -- layer=1 filter=104 channel=28
    5, -6, 6, 0, 3, 4, -9, 5, 9,
    -- layer=1 filter=104 channel=29
    5, -6, 2, -12, 0, 5, -12, -10, -8,
    -- layer=1 filter=104 channel=30
    -1, 1, -2, 0, 8, -8, -11, 2, 10,
    -- layer=1 filter=104 channel=31
    5, 1, -11, -2, 2, -13, -4, 3, -5,
    -- layer=1 filter=104 channel=32
    -2, -9, -3, -5, 3, 0, -6, 2, -1,
    -- layer=1 filter=104 channel=33
    1, -5, 8, -6, -10, -9, -4, -5, 6,
    -- layer=1 filter=104 channel=34
    -9, 9, 8, 1, 5, 5, 1, -6, 8,
    -- layer=1 filter=104 channel=35
    -4, 1, 8, 11, 4, 4, 7, -5, 0,
    -- layer=1 filter=104 channel=36
    -2, 8, -10, -7, -8, 1, 6, -1, -9,
    -- layer=1 filter=104 channel=37
    3, 6, 7, -5, 5, -4, 2, -9, -4,
    -- layer=1 filter=104 channel=38
    -11, -5, -11, 4, -11, -3, 5, 7, 4,
    -- layer=1 filter=104 channel=39
    0, -5, -1, -4, -7, -4, 4, 3, 8,
    -- layer=1 filter=104 channel=40
    -10, 5, -1, 4, 4, 0, -5, 0, 0,
    -- layer=1 filter=104 channel=41
    -1, -10, -9, -6, 4, -7, -1, -8, 7,
    -- layer=1 filter=104 channel=42
    -6, 13, 3, -12, 3, -4, -5, -1, 4,
    -- layer=1 filter=104 channel=43
    -4, -10, 1, 5, 7, -1, -11, 2, 6,
    -- layer=1 filter=104 channel=44
    -5, -4, 6, 6, -9, 0, 3, -4, 5,
    -- layer=1 filter=104 channel=45
    -6, 7, 1, 4, -9, 0, 6, 4, -4,
    -- layer=1 filter=104 channel=46
    6, 4, 15, 1, -6, -5, 2, -2, -5,
    -- layer=1 filter=104 channel=47
    5, 8, 0, -6, 0, -4, -4, 3, 5,
    -- layer=1 filter=104 channel=48
    -1, 5, 7, 5, -2, -3, 8, -10, -11,
    -- layer=1 filter=104 channel=49
    8, -11, -4, -4, -5, -2, -3, -6, -7,
    -- layer=1 filter=104 channel=50
    5, 1, 7, 6, 3, 1, 5, 5, -5,
    -- layer=1 filter=104 channel=51
    -3, -8, -9, 8, -1, -8, -8, 0, 3,
    -- layer=1 filter=104 channel=52
    4, -7, 0, 2, -5, -3, -1, -7, 1,
    -- layer=1 filter=104 channel=53
    2, 9, -3, -4, -7, -10, 9, 8, 7,
    -- layer=1 filter=104 channel=54
    -10, 1, 2, 2, -4, -6, 4, -1, -3,
    -- layer=1 filter=104 channel=55
    7, -1, 0, -8, -10, 9, -1, -11, -12,
    -- layer=1 filter=104 channel=56
    8, -2, -5, 4, -2, 6, 9, -8, 0,
    -- layer=1 filter=104 channel=57
    -12, 0, 3, -10, 5, -3, 0, 1, 1,
    -- layer=1 filter=104 channel=58
    -12, -8, 9, 3, -5, -6, 3, 3, -8,
    -- layer=1 filter=104 channel=59
    3, -8, 3, -3, 5, 8, -4, -1, 4,
    -- layer=1 filter=104 channel=60
    -5, -6, -10, -3, 6, 6, -8, -3, -2,
    -- layer=1 filter=104 channel=61
    0, 5, 3, 3, -5, 9, 0, 4, -7,
    -- layer=1 filter=104 channel=62
    -4, 5, -2, -1, 8, -12, -2, 0, -6,
    -- layer=1 filter=104 channel=63
    -2, -10, -7, -13, 3, 0, 0, -5, 3,
    -- layer=1 filter=104 channel=64
    0, 8, -9, -11, -9, 8, -5, -8, -6,
    -- layer=1 filter=104 channel=65
    -8, -9, 2, -11, -1, -4, -4, -7, 5,
    -- layer=1 filter=104 channel=66
    3, 0, -11, 2, -5, -3, 3, -3, 0,
    -- layer=1 filter=104 channel=67
    3, 3, -8, 9, -2, 7, 0, 4, -10,
    -- layer=1 filter=104 channel=68
    9, -5, 0, 8, -3, -9, 7, 6, -10,
    -- layer=1 filter=104 channel=69
    1, -8, 4, 4, -13, -7, -14, 2, 3,
    -- layer=1 filter=104 channel=70
    1, 0, 2, 10, -4, 1, 8, 3, 3,
    -- layer=1 filter=104 channel=71
    6, 2, -7, 0, -13, 5, -8, -1, -9,
    -- layer=1 filter=104 channel=72
    -12, 1, -1, 2, -3, -4, -11, -5, -2,
    -- layer=1 filter=104 channel=73
    -9, -7, -4, -9, -11, -6, 8, 8, 1,
    -- layer=1 filter=104 channel=74
    -8, 0, 9, 8, -4, 5, 0, -7, 1,
    -- layer=1 filter=104 channel=75
    -10, -12, 1, -10, -5, 3, -11, 4, 8,
    -- layer=1 filter=104 channel=76
    -7, -5, 6, 4, 3, -8, -11, -12, 8,
    -- layer=1 filter=104 channel=77
    -2, 1, 5, -2, 4, -8, -6, -2, 2,
    -- layer=1 filter=104 channel=78
    6, -6, -9, 3, 9, 8, -10, -5, 1,
    -- layer=1 filter=104 channel=79
    4, -4, 4, 2, 1, 6, 10, -7, 1,
    -- layer=1 filter=104 channel=80
    9, -2, -2, 0, 4, 6, 8, -4, 8,
    -- layer=1 filter=104 channel=81
    -4, -2, -2, -3, -5, 3, -12, -9, 0,
    -- layer=1 filter=104 channel=82
    0, -4, 6, 4, 4, -9, -8, -8, 8,
    -- layer=1 filter=104 channel=83
    -3, -7, 6, 7, -10, -9, -11, -12, -1,
    -- layer=1 filter=104 channel=84
    -4, 0, 0, -8, 0, -3, -12, -3, -4,
    -- layer=1 filter=104 channel=85
    8, 9, 3, -7, 3, 2, 2, -5, -5,
    -- layer=1 filter=104 channel=86
    -4, -10, -8, -8, -2, -3, -7, 4, 0,
    -- layer=1 filter=104 channel=87
    3, 2, 8, -8, -10, -8, 0, 7, -6,
    -- layer=1 filter=104 channel=88
    -7, 1, -11, -8, 8, -11, -1, -4, 0,
    -- layer=1 filter=104 channel=89
    -11, -10, 1, -4, -3, -11, 1, 7, -6,
    -- layer=1 filter=104 channel=90
    0, 3, -6, -5, 7, 2, -10, -6, 0,
    -- layer=1 filter=104 channel=91
    2, -8, 3, -1, -10, -4, -10, -8, 6,
    -- layer=1 filter=104 channel=92
    -6, -9, -7, -10, 1, -8, -10, -4, 6,
    -- layer=1 filter=104 channel=93
    -1, 0, 7, -9, 0, 0, 1, 0, -7,
    -- layer=1 filter=104 channel=94
    -8, -5, 2, 0, -5, 1, -4, -5, -9,
    -- layer=1 filter=104 channel=95
    7, -10, 5, -9, -8, -7, -13, 6, 0,
    -- layer=1 filter=104 channel=96
    -10, 0, -10, -5, -1, 3, 6, 0, 3,
    -- layer=1 filter=104 channel=97
    3, -5, -4, 3, 0, 6, 3, -2, 6,
    -- layer=1 filter=104 channel=98
    0, -3, -3, -7, 5, 0, -7, -6, 7,
    -- layer=1 filter=104 channel=99
    -6, 7, -9, -8, -1, 7, -9, -1, -1,
    -- layer=1 filter=104 channel=100
    -4, -1, -6, -12, -8, -5, -7, -4, 5,
    -- layer=1 filter=104 channel=101
    3, -6, 3, 1, -11, 8, 2, 1, 3,
    -- layer=1 filter=104 channel=102
    -11, -10, 1, -6, -5, 3, -5, -4, -10,
    -- layer=1 filter=104 channel=103
    1, 6, -1, -6, -8, -5, -2, -7, 1,
    -- layer=1 filter=104 channel=104
    2, -4, 8, -1, -7, 0, -7, 3, -8,
    -- layer=1 filter=104 channel=105
    3, 1, -8, -1, 2, 2, 6, 2, -5,
    -- layer=1 filter=104 channel=106
    -6, -5, -14, -11, -7, 5, 4, -9, -1,
    -- layer=1 filter=104 channel=107
    -7, 0, 7, -7, -6, -2, -1, -11, -11,
    -- layer=1 filter=104 channel=108
    -2, 1, -4, 6, -6, -6, -8, 7, -11,
    -- layer=1 filter=104 channel=109
    7, 0, -7, 2, -6, 8, -5, 10, 4,
    -- layer=1 filter=104 channel=110
    5, -5, -3, -2, 2, -3, -7, 6, -1,
    -- layer=1 filter=104 channel=111
    -8, 7, 2, -10, -1, -4, -3, -5, -11,
    -- layer=1 filter=104 channel=112
    -4, -9, -11, 0, -9, 3, 0, -11, 7,
    -- layer=1 filter=104 channel=113
    0, -5, 2, -5, -2, 3, -2, 4, -6,
    -- layer=1 filter=104 channel=114
    11, 11, -4, 8, 0, -7, 4, -5, 3,
    -- layer=1 filter=104 channel=115
    0, -5, -4, -3, 2, -9, -9, -9, -3,
    -- layer=1 filter=104 channel=116
    3, -1, -6, 1, 0, 4, 7, 3, -1,
    -- layer=1 filter=104 channel=117
    -1, -10, -3, -2, -4, -3, -4, -4, -14,
    -- layer=1 filter=104 channel=118
    -4, -7, -3, -10, -1, 9, 6, -5, -4,
    -- layer=1 filter=104 channel=119
    -12, -5, 2, 3, 0, -9, -13, -9, 2,
    -- layer=1 filter=104 channel=120
    -12, -10, 0, -2, 4, -7, -1, -5, 8,
    -- layer=1 filter=104 channel=121
    0, 5, 9, -17, -16, -8, -13, -5, 6,
    -- layer=1 filter=104 channel=122
    3, -4, 1, -9, 2, 0, -7, 8, 0,
    -- layer=1 filter=104 channel=123
    -12, 4, -2, 2, -11, -8, -4, 5, -2,
    -- layer=1 filter=104 channel=124
    3, 1, -3, -8, -3, 6, 5, -8, 1,
    -- layer=1 filter=104 channel=125
    -8, -8, 1, -3, -5, -5, 2, 0, 1,
    -- layer=1 filter=104 channel=126
    7, 8, -3, 8, 9, -2, 1, -11, 0,
    -- layer=1 filter=104 channel=127
    1, -5, -6, -6, -1, 6, -8, 5, 8,
    -- layer=1 filter=105 channel=0
    -7, 0, 7, 4, -9, -7, -12, -11, 4,
    -- layer=1 filter=105 channel=1
    0, 4, -7, -4, -4, 6, -11, 5, -1,
    -- layer=1 filter=105 channel=2
    5, -8, -4, -2, -4, 8, 1, 9, 0,
    -- layer=1 filter=105 channel=3
    0, -9, -1, 3, 4, -4, 1, -2, 8,
    -- layer=1 filter=105 channel=4
    -10, 5, -1, 1, -6, -5, -5, -7, -4,
    -- layer=1 filter=105 channel=5
    1, -6, 1, -1, 1, -6, -14, -14, -8,
    -- layer=1 filter=105 channel=6
    -3, -5, -8, 9, -2, -5, 2, 6, 9,
    -- layer=1 filter=105 channel=7
    -9, 0, 3, 0, 0, 2, 4, -15, -4,
    -- layer=1 filter=105 channel=8
    3, -3, 8, -10, -10, -3, 2, -3, -8,
    -- layer=1 filter=105 channel=9
    1, -3, -7, -11, 0, -5, -1, -10, -12,
    -- layer=1 filter=105 channel=10
    2, -4, -10, 5, -8, -7, -6, 9, 4,
    -- layer=1 filter=105 channel=11
    0, -2, -11, 4, -12, -9, 0, -10, 3,
    -- layer=1 filter=105 channel=12
    -9, -7, 4, 5, 5, 9, 11, 5, -7,
    -- layer=1 filter=105 channel=13
    6, -7, 6, 9, 8, -4, 5, 3, -10,
    -- layer=1 filter=105 channel=14
    7, 2, 0, 1, -8, -15, -8, 7, -7,
    -- layer=1 filter=105 channel=15
    3, -12, -9, -7, -4, -4, -8, 2, -6,
    -- layer=1 filter=105 channel=16
    -8, -4, -13, -6, 0, 6, -6, 2, -3,
    -- layer=1 filter=105 channel=17
    -9, -7, 3, -7, -10, 3, 0, 0, -2,
    -- layer=1 filter=105 channel=18
    -10, -10, 0, -4, 0, 6, -10, -7, -4,
    -- layer=1 filter=105 channel=19
    4, -11, -5, -3, 3, 3, 6, -9, 0,
    -- layer=1 filter=105 channel=20
    1, -1, -4, -11, -8, 3, -6, -2, -6,
    -- layer=1 filter=105 channel=21
    -3, -1, 5, -8, 6, -3, -7, 4, -6,
    -- layer=1 filter=105 channel=22
    -2, -1, -6, -5, 1, -8, 4, -6, -14,
    -- layer=1 filter=105 channel=23
    -8, 7, 9, -12, 9, -7, -9, 7, -2,
    -- layer=1 filter=105 channel=24
    4, 4, -2, 6, 4, 3, -1, -15, -6,
    -- layer=1 filter=105 channel=25
    -3, -7, -1, -17, -7, -5, -10, -6, -14,
    -- layer=1 filter=105 channel=26
    0, 3, -7, -10, -13, 0, 2, -5, -7,
    -- layer=1 filter=105 channel=27
    -3, -3, 0, -4, 7, -9, -10, -3, 0,
    -- layer=1 filter=105 channel=28
    4, -2, -2, -6, 0, -10, -6, -7, 4,
    -- layer=1 filter=105 channel=29
    6, -11, -12, -6, 5, -2, -3, -4, -6,
    -- layer=1 filter=105 channel=30
    -1, 6, -1, -2, 7, -5, 5, -5, 5,
    -- layer=1 filter=105 channel=31
    0, -9, 1, 0, 8, 13, -3, 2, -4,
    -- layer=1 filter=105 channel=32
    -7, 0, -4, 5, 2, 2, 0, -1, 4,
    -- layer=1 filter=105 channel=33
    12, 7, -8, 3, 4, 7, 3, 9, 0,
    -- layer=1 filter=105 channel=34
    -9, -1, 2, 7, 7, -1, -2, -7, 0,
    -- layer=1 filter=105 channel=35
    -10, -7, 2, -5, -7, -2, -12, 5, -11,
    -- layer=1 filter=105 channel=36
    0, -4, -6, -4, -9, 4, 1, -8, 6,
    -- layer=1 filter=105 channel=37
    2, -1, 3, -10, -5, -10, -10, 0, 0,
    -- layer=1 filter=105 channel=38
    -1, -1, -1, -9, 1, 10, -9, 0, -11,
    -- layer=1 filter=105 channel=39
    -7, 0, -5, 7, -4, 5, -5, -2, -2,
    -- layer=1 filter=105 channel=40
    -5, 0, -1, 7, -10, -4, 8, 6, 9,
    -- layer=1 filter=105 channel=41
    2, 6, -1, -8, -3, -2, -4, -2, -1,
    -- layer=1 filter=105 channel=42
    -4, -8, -9, -9, -2, -9, 6, 3, 1,
    -- layer=1 filter=105 channel=43
    2, -8, 0, 8, -7, -2, -8, 3, -6,
    -- layer=1 filter=105 channel=44
    0, -7, -9, -5, -14, -1, 6, 4, 7,
    -- layer=1 filter=105 channel=45
    -4, -2, 0, 2, 5, 5, 0, 0, 6,
    -- layer=1 filter=105 channel=46
    -2, 5, -6, 9, -6, 0, 10, 6, -3,
    -- layer=1 filter=105 channel=47
    -6, -8, 5, -6, 8, -3, 3, 4, 1,
    -- layer=1 filter=105 channel=48
    0, -8, -8, 5, -12, -6, 6, -8, -5,
    -- layer=1 filter=105 channel=49
    2, -13, 4, -7, -5, -8, -7, -15, -13,
    -- layer=1 filter=105 channel=50
    1, 0, -2, 3, 7, -6, 4, -10, 6,
    -- layer=1 filter=105 channel=51
    -8, 3, -8, -8, -9, -5, 3, 7, -11,
    -- layer=1 filter=105 channel=52
    9, 9, -1, 1, 3, 5, -10, 1, -7,
    -- layer=1 filter=105 channel=53
    5, 2, 0, -2, -1, -5, 0, 6, -9,
    -- layer=1 filter=105 channel=54
    0, 1, -1, -12, -4, 4, -1, 6, 6,
    -- layer=1 filter=105 channel=55
    -1, -11, -2, 1, 4, -7, 4, -10, -5,
    -- layer=1 filter=105 channel=56
    2, -9, 9, 9, 2, -10, 6, 0, 1,
    -- layer=1 filter=105 channel=57
    3, -13, -11, -4, 0, 5, -11, 0, -3,
    -- layer=1 filter=105 channel=58
    0, 0, -2, 0, -9, 4, 0, -2, 2,
    -- layer=1 filter=105 channel=59
    7, -9, -6, 4, -1, 4, -4, -9, 6,
    -- layer=1 filter=105 channel=60
    -1, 2, -6, -5, -8, -5, -10, -7, -9,
    -- layer=1 filter=105 channel=61
    8, 1, -5, -7, -11, 2, 6, -2, 8,
    -- layer=1 filter=105 channel=62
    2, 3, -3, -8, 3, -13, 3, 2, -8,
    -- layer=1 filter=105 channel=63
    -11, -13, -7, -9, -4, 7, 5, -6, 3,
    -- layer=1 filter=105 channel=64
    -9, 5, 5, 5, 3, -11, 3, -12, -2,
    -- layer=1 filter=105 channel=65
    0, -7, 6, -7, 3, -10, 6, -13, 3,
    -- layer=1 filter=105 channel=66
    -8, -9, 7, -4, -4, -2, -6, -9, 0,
    -- layer=1 filter=105 channel=67
    8, -9, -2, 1, -6, -3, -5, 4, 9,
    -- layer=1 filter=105 channel=68
    -7, -9, 0, 8, -2, -10, 0, -11, 0,
    -- layer=1 filter=105 channel=69
    -1, -14, 0, 0, -10, 0, -3, -7, -6,
    -- layer=1 filter=105 channel=70
    -7, -5, 0, 8, -6, -3, 11, 10, 8,
    -- layer=1 filter=105 channel=71
    -1, 0, -2, 0, 3, -12, -13, -3, -7,
    -- layer=1 filter=105 channel=72
    -10, 1, -4, -7, 5, 2, -6, -1, 6,
    -- layer=1 filter=105 channel=73
    -3, 0, 3, -11, 7, 6, 5, -2, 3,
    -- layer=1 filter=105 channel=74
    -5, 0, 2, -7, 6, -3, 7, 6, 0,
    -- layer=1 filter=105 channel=75
    5, -3, -2, -11, -8, 2, -1, -7, -8,
    -- layer=1 filter=105 channel=76
    -7, 2, -2, -3, 2, 3, -10, 3, 5,
    -- layer=1 filter=105 channel=77
    8, 5, 0, -9, 6, -8, 0, 2, -2,
    -- layer=1 filter=105 channel=78
    -7, 6, -7, 7, -3, 4, -4, 9, -10,
    -- layer=1 filter=105 channel=79
    -2, -12, -7, -17, -7, -3, -6, -9, 1,
    -- layer=1 filter=105 channel=80
    -5, 5, 2, -10, -4, -9, -6, -9, 0,
    -- layer=1 filter=105 channel=81
    7, 5, 2, -6, 6, 3, -7, 6, 3,
    -- layer=1 filter=105 channel=82
    2, 8, 6, -13, -9, 7, -2, -8, -9,
    -- layer=1 filter=105 channel=83
    0, 5, -5, -9, 4, 0, -10, -7, 1,
    -- layer=1 filter=105 channel=84
    -3, -2, -3, 0, -17, -3, -11, -3, -7,
    -- layer=1 filter=105 channel=85
    -8, 2, 5, -5, -10, -2, 1, -5, 0,
    -- layer=1 filter=105 channel=86
    -9, -3, -9, -2, 0, -5, -8, 3, 2,
    -- layer=1 filter=105 channel=87
    -8, -6, -3, -7, -9, 0, 5, 5, 0,
    -- layer=1 filter=105 channel=88
    -10, -9, 0, 6, 0, 0, 2, 2, -6,
    -- layer=1 filter=105 channel=89
    3, -2, 7, -9, 6, 6, -8, 0, 0,
    -- layer=1 filter=105 channel=90
    -11, -12, -6, -10, 5, -8, -7, -13, 2,
    -- layer=1 filter=105 channel=91
    -1, 3, 6, 5, 0, 12, 1, 1, -6,
    -- layer=1 filter=105 channel=92
    -6, 0, -10, -9, -1, 3, -11, -4, -9,
    -- layer=1 filter=105 channel=93
    -1, 5, -11, -12, -3, -2, -7, -3, -6,
    -- layer=1 filter=105 channel=94
    -10, 6, 1, 1, 5, -11, 0, 2, -4,
    -- layer=1 filter=105 channel=95
    -11, 4, 2, -12, 0, -3, 3, -12, 7,
    -- layer=1 filter=105 channel=96
    -1, -2, -6, -1, 0, -10, 0, -10, -5,
    -- layer=1 filter=105 channel=97
    0, -3, 1, 0, 2, -10, -9, 3, -8,
    -- layer=1 filter=105 channel=98
    3, 6, -9, -12, 0, -2, 1, -6, -4,
    -- layer=1 filter=105 channel=99
    -9, 10, -10, -9, 0, -8, 0, -5, 9,
    -- layer=1 filter=105 channel=100
    8, -1, -6, 7, 7, 0, 2, 7, 5,
    -- layer=1 filter=105 channel=101
    -9, 6, 7, 5, -5, 5, -11, -11, -10,
    -- layer=1 filter=105 channel=102
    -3, 0, 0, 0, 4, -9, -9, -5, -4,
    -- layer=1 filter=105 channel=103
    7, -4, 4, -5, -6, 4, -5, -10, -8,
    -- layer=1 filter=105 channel=104
    4, 2, 0, -1, -9, 4, -3, 1, 8,
    -- layer=1 filter=105 channel=105
    6, 2, 0, -3, 4, -10, -1, 3, -6,
    -- layer=1 filter=105 channel=106
    -4, -12, 3, -3, -6, 0, -1, -4, -3,
    -- layer=1 filter=105 channel=107
    -2, -1, 1, -2, -9, 2, 0, -4, 7,
    -- layer=1 filter=105 channel=108
    -2, 3, -8, 5, -2, -14, -15, -2, 2,
    -- layer=1 filter=105 channel=109
    -3, -4, 10, -3, 0, -1, 2, 0, 3,
    -- layer=1 filter=105 channel=110
    0, -7, -7, 8, -10, -1, 7, -4, -9,
    -- layer=1 filter=105 channel=111
    0, 5, -12, -2, 5, 3, 3, -3, -8,
    -- layer=1 filter=105 channel=112
    6, -9, -7, 9, -8, -6, -5, 2, -4,
    -- layer=1 filter=105 channel=113
    -8, -6, -5, -9, 0, 1, -11, -8, 0,
    -- layer=1 filter=105 channel=114
    -5, 1, -12, -9, 4, -11, 2, 4, -5,
    -- layer=1 filter=105 channel=115
    6, -4, -8, 6, -7, 1, -5, 9, 0,
    -- layer=1 filter=105 channel=116
    -3, -2, -5, 6, -10, 5, 5, 8, 7,
    -- layer=1 filter=105 channel=117
    9, -9, -13, 0, -7, -9, -1, 7, -3,
    -- layer=1 filter=105 channel=118
    -5, -8, -5, -7, -11, 3, -6, 1, 3,
    -- layer=1 filter=105 channel=119
    -4, -11, -9, -7, -2, -3, -1, -12, 7,
    -- layer=1 filter=105 channel=120
    3, -2, -3, -5, 2, 1, -14, -9, -14,
    -- layer=1 filter=105 channel=121
    6, -12, 0, 0, 3, -2, -10, 5, -7,
    -- layer=1 filter=105 channel=122
    -9, 1, 8, -10, -6, -2, 6, -3, 6,
    -- layer=1 filter=105 channel=123
    -3, -7, 4, 6, -6, 6, -1, 6, -11,
    -- layer=1 filter=105 channel=124
    -9, -8, -1, -1, -2, 5, -3, -1, 7,
    -- layer=1 filter=105 channel=125
    -2, 6, 6, -6, 11, -1, 1, 3, -6,
    -- layer=1 filter=105 channel=126
    5, -5, -2, -11, -6, -9, 2, -3, 5,
    -- layer=1 filter=105 channel=127
    -3, 3, 3, -12, -14, -8, 0, -3, 0,
    -- layer=1 filter=106 channel=0
    3, -6, -3, 20, 10, -7, -4, -5, 10,
    -- layer=1 filter=106 channel=1
    -13, 30, 8, -10, 6, 33, 4, 8, 5,
    -- layer=1 filter=106 channel=2
    -3, 50, 32, -10, -13, -14, -5, -15, 4,
    -- layer=1 filter=106 channel=3
    2, -3, 3, 0, 6, -2, 9, 5, 1,
    -- layer=1 filter=106 channel=4
    -2, 13, -3, 7, -10, -4, -11, -10, 6,
    -- layer=1 filter=106 channel=5
    5, 48, 6, -28, 15, 17, 14, 13, 28,
    -- layer=1 filter=106 channel=6
    -7, 47, 56, -53, 1, 35, -80, -41, -33,
    -- layer=1 filter=106 channel=7
    -58, -16, 56, -73, -55, -12, -47, -81, -35,
    -- layer=1 filter=106 channel=8
    12, 27, 0, 7, 11, 4, 2, 16, 29,
    -- layer=1 filter=106 channel=9
    -2, 4, 1, 56, 0, 10, -59, -6, 43,
    -- layer=1 filter=106 channel=10
    -39, -5, 47, -58, -51, -8, -53, -84, -4,
    -- layer=1 filter=106 channel=11
    11, -23, -18, 22, 4, 0, 19, 18, 13,
    -- layer=1 filter=106 channel=12
    1, -8, 39, -7, -10, -30, 8, 25, 55,
    -- layer=1 filter=106 channel=13
    38, 50, 33, -13, 0, -15, -26, -24, -24,
    -- layer=1 filter=106 channel=14
    -42, -24, 49, -4, 19, -21, -48, -86, -3,
    -- layer=1 filter=106 channel=15
    35, 32, 8, -36, 5, 0, 18, -16, 25,
    -- layer=1 filter=106 channel=16
    -14, 13, -11, -30, -3, -19, 5, 14, 26,
    -- layer=1 filter=106 channel=17
    37, 2, -17, 10, 21, -8, -1, -3, 10,
    -- layer=1 filter=106 channel=18
    -4, -5, -2, 19, 12, -20, 14, 16, 10,
    -- layer=1 filter=106 channel=19
    31, 43, 45, 64, 30, 21, 15, 36, 66,
    -- layer=1 filter=106 channel=20
    26, 45, 29, -37, -11, -17, -25, -20, -30,
    -- layer=1 filter=106 channel=21
    -41, 23, 24, -30, -29, -24, -32, -45, -50,
    -- layer=1 filter=106 channel=22
    -16, 13, 6, -36, -15, 0, -18, -28, -8,
    -- layer=1 filter=106 channel=23
    -16, 16, 38, -55, -29, -4, -31, -14, -25,
    -- layer=1 filter=106 channel=24
    13, 18, 11, -21, -22, -6, -22, -25, 0,
    -- layer=1 filter=106 channel=25
    -62, -3, 27, -51, -59, -14, -27, -49, -1,
    -- layer=1 filter=106 channel=26
    55, 33, 1, -16, -2, -10, -31, -13, -21,
    -- layer=1 filter=106 channel=27
    -48, -56, -62, -34, -38, -20, 14, -2, 4,
    -- layer=1 filter=106 channel=28
    -46, -23, 52, -56, -55, -20, -37, -64, -8,
    -- layer=1 filter=106 channel=29
    -36, -30, -30, -27, -37, -4, -22, -2, -13,
    -- layer=1 filter=106 channel=30
    2, 3, 27, 66, 29, -1, -1, 3, 21,
    -- layer=1 filter=106 channel=31
    -27, 3, 13, -9, 0, -45, -11, -31, -7,
    -- layer=1 filter=106 channel=32
    49, 22, 12, 3, -12, -4, -32, -21, -22,
    -- layer=1 filter=106 channel=33
    0, -10, 0, 9, -1, 14, -1, -7, 8,
    -- layer=1 filter=106 channel=34
    -13, 6, 21, -7, -1, 32, -2, -22, 10,
    -- layer=1 filter=106 channel=35
    -3, 7, -4, -8, -13, 3, -4, -17, 0,
    -- layer=1 filter=106 channel=36
    24, -10, -19, 40, 13, 15, 38, 42, 20,
    -- layer=1 filter=106 channel=37
    7, 35, 21, 1, 19, 5, 14, 3, 36,
    -- layer=1 filter=106 channel=38
    19, 58, 26, -30, -19, -23, -56, -49, -41,
    -- layer=1 filter=106 channel=39
    -8, -22, -23, -7, 11, -9, 11, 0, 20,
    -- layer=1 filter=106 channel=40
    -44, -3, 0, -22, -24, -44, -47, -39, -52,
    -- layer=1 filter=106 channel=41
    57, 10, 0, 58, -7, -8, -29, 27, 21,
    -- layer=1 filter=106 channel=42
    2, 60, 49, -33, 12, -8, -16, -19, 4,
    -- layer=1 filter=106 channel=43
    -19, -2, -10, -19, 3, -6, 1, -1, 26,
    -- layer=1 filter=106 channel=44
    57, 16, 13, -10, -10, 11, -24, -37, -16,
    -- layer=1 filter=106 channel=45
    23, 10, 10, -34, -6, -21, -32, -23, -19,
    -- layer=1 filter=106 channel=46
    71, 90, 71, 36, 43, 39, 23, 25, 31,
    -- layer=1 filter=106 channel=47
    -15, -11, 34, -27, -48, -6, -35, -23, -33,
    -- layer=1 filter=106 channel=48
    -8, 16, 19, -14, -1, -9, -24, -35, -41,
    -- layer=1 filter=106 channel=49
    -5, 21, 11, -15, -8, 19, -48, -38, -18,
    -- layer=1 filter=106 channel=50
    -21, 0, 15, 13, 0, -10, -2, -30, 7,
    -- layer=1 filter=106 channel=51
    -4, 18, 40, -47, -40, -8, -71, -74, -36,
    -- layer=1 filter=106 channel=52
    -2, -1, 2, 9, 12, 11, 5, 6, 24,
    -- layer=1 filter=106 channel=53
    16, 0, -1, -12, 10, 7, 1, 6, 3,
    -- layer=1 filter=106 channel=54
    -27, -3, 12, -31, -43, -17, -17, -22, 19,
    -- layer=1 filter=106 channel=55
    -8, -18, -25, 14, 15, 14, 27, 30, 23,
    -- layer=1 filter=106 channel=56
    -10, -9, -11, 1, -7, -11, -11, -5, 6,
    -- layer=1 filter=106 channel=57
    -64, -1, 37, -65, -77, -37, -65, -105, -44,
    -- layer=1 filter=106 channel=58
    -74, 0, 27, -109, -96, -54, -65, -85, -50,
    -- layer=1 filter=106 channel=59
    -4, -10, -15, -3, -12, -8, -12, -7, -18,
    -- layer=1 filter=106 channel=60
    11, 6, 0, 23, 13, 20, 24, 4, -8,
    -- layer=1 filter=106 channel=61
    9, 4, -9, 6, 7, 5, -4, 0, -6,
    -- layer=1 filter=106 channel=62
    16, 38, 6, 1, 9, 19, 3, 15, 50,
    -- layer=1 filter=106 channel=63
    -13, -31, -9, 25, 14, 0, 15, 24, 13,
    -- layer=1 filter=106 channel=64
    -7, 23, 20, 6, -3, 6, 3, 7, 1,
    -- layer=1 filter=106 channel=65
    2, 25, 21, -6, -26, -12, -19, -13, -29,
    -- layer=1 filter=106 channel=66
    -4, -15, -13, 8, 2, 10, 9, 20, 18,
    -- layer=1 filter=106 channel=67
    64, 67, 63, 42, 60, 100, -38, -18, -38,
    -- layer=1 filter=106 channel=68
    59, 11, 7, -26, 9, -10, -33, -30, -6,
    -- layer=1 filter=106 channel=69
    22, 33, 18, -9, 2, -6, 4, -10, -3,
    -- layer=1 filter=106 channel=70
    27, 64, 31, -28, 28, 74, -74, -43, -39,
    -- layer=1 filter=106 channel=71
    -20, -1, -3, -34, -23, -2, -22, -13, 6,
    -- layer=1 filter=106 channel=72
    0, 27, -3, 83, 20, 17, 8, 20, 60,
    -- layer=1 filter=106 channel=73
    -7, -2, 3, 6, 3, -10, 8, 9, 2,
    -- layer=1 filter=106 channel=74
    1, 24, -12, 2, -6, 1, -52, -14, -9,
    -- layer=1 filter=106 channel=75
    -15, -18, 6, 34, 16, -27, -26, 31, 29,
    -- layer=1 filter=106 channel=76
    24, 6, -9, 31, 0, 0, -3, -1, 1,
    -- layer=1 filter=106 channel=77
    -25, -17, -19, -38, -26, -29, -45, -47, -17,
    -- layer=1 filter=106 channel=78
    -16, -2, 2, 4, -7, -10, 0, 10, -6,
    -- layer=1 filter=106 channel=79
    15, 29, 0, -14, 0, -1, 13, 3, 22,
    -- layer=1 filter=106 channel=80
    8, -2, -4, -7, 5, -8, 4, 0, 11,
    -- layer=1 filter=106 channel=81
    -33, -25, -20, -32, -26, -23, -21, -9, 1,
    -- layer=1 filter=106 channel=82
    -18, 25, 42, -55, -36, -9, -65, -56, -59,
    -- layer=1 filter=106 channel=83
    29, 18, -10, 0, 27, 4, 7, -9, 4,
    -- layer=1 filter=106 channel=84
    23, -7, 0, 22, -4, -13, -25, -4, 2,
    -- layer=1 filter=106 channel=85
    -12, 11, 16, -23, -57, -12, -58, -34, -8,
    -- layer=1 filter=106 channel=86
    18, -9, 5, 22, 14, 6, 14, 13, 13,
    -- layer=1 filter=106 channel=87
    23, 52, 58, 89, 56, 39, -24, 32, 59,
    -- layer=1 filter=106 channel=88
    21, 16, 23, -9, -8, -6, -21, -24, -13,
    -- layer=1 filter=106 channel=89
    -29, -5, 26, -54, -42, -28, -61, -54, -50,
    -- layer=1 filter=106 channel=90
    61, 24, 2, -5, 18, 3, -35, -45, -18,
    -- layer=1 filter=106 channel=91
    -7, 29, 28, -33, -10, -11, -54, -47, -66,
    -- layer=1 filter=106 channel=92
    34, 27, -36, -30, -21, -17, -40, -5, 17,
    -- layer=1 filter=106 channel=93
    6, -2, 7, -27, -15, -3, -18, -15, -9,
    -- layer=1 filter=106 channel=94
    -8, -3, -7, 16, -12, -10, 13, 12, 1,
    -- layer=1 filter=106 channel=95
    10, -5, 0, 33, 12, -2, -19, 15, 18,
    -- layer=1 filter=106 channel=96
    0, 8, 5, 8, 13, 1, 9, 11, 19,
    -- layer=1 filter=106 channel=97
    3, -12, 2, -5, -2, 2, 6, -3, 7,
    -- layer=1 filter=106 channel=98
    -2, 7, -13, 7, 22, -7, 0, 14, 19,
    -- layer=1 filter=106 channel=99
    -25, -43, 11, -15, -88, -56, -61, -78, -23,
    -- layer=1 filter=106 channel=100
    -13, -13, -37, 7, 4, -15, 30, 23, 17,
    -- layer=1 filter=106 channel=101
    -2, 34, 43, -34, -5, -8, -46, -50, -57,
    -- layer=1 filter=106 channel=102
    11, 7, -3, 0, -9, -6, 0, -9, -7,
    -- layer=1 filter=106 channel=103
    4, -25, -15, 18, -9, 2, 18, 8, 2,
    -- layer=1 filter=106 channel=104
    -3, 30, 20, 7, -7, 4, -15, 0, -1,
    -- layer=1 filter=106 channel=105
    -4, -25, -6, 19, 7, 12, 14, 14, 22,
    -- layer=1 filter=106 channel=106
    38, 41, 20, -42, -10, -16, -58, -50, -47,
    -- layer=1 filter=106 channel=107
    8, -2, 12, -2, 0, -8, 11, 3, 0,
    -- layer=1 filter=106 channel=108
    71, 42, 20, 0, 4, -10, -46, -45, -30,
    -- layer=1 filter=106 channel=109
    9, 9, 2, -2, -5, -10, 0, 10, 6,
    -- layer=1 filter=106 channel=110
    -7, -14, 8, 5, -4, -11, 3, -5, 8,
    -- layer=1 filter=106 channel=111
    3, 0, 19, 34, 6, -12, 0, 9, -4,
    -- layer=1 filter=106 channel=112
    16, 15, 16, 17, 11, 22, -8, 0, 0,
    -- layer=1 filter=106 channel=113
    -6, 47, 13, -24, 16, 16, -25, -27, -44,
    -- layer=1 filter=106 channel=114
    0, -1, -4, -19, 16, -3, 34, -3, 0,
    -- layer=1 filter=106 channel=115
    -19, -4, -10, 3, 1, 2, -5, 2, 25,
    -- layer=1 filter=106 channel=116
    -3, 3, 9, -9, -4, 2, -4, 0, -8,
    -- layer=1 filter=106 channel=117
    18, 24, 30, 42, 31, 12, -15, -25, 3,
    -- layer=1 filter=106 channel=118
    -5, 0, -12, 25, -2, -15, -17, 8, 11,
    -- layer=1 filter=106 channel=119
    53, 14, 18, 11, 3, 7, -37, -36, -23,
    -- layer=1 filter=106 channel=120
    -44, 22, 40, -42, -44, -5, -36, -44, -18,
    -- layer=1 filter=106 channel=121
    -15, -9, -2, 21, 43, 7, 20, 44, 41,
    -- layer=1 filter=106 channel=122
    0, -6, -3, 9, 8, -2, -8, 3, 1,
    -- layer=1 filter=106 channel=123
    -30, -38, -36, 8, -7, -23, 18, 20, 26,
    -- layer=1 filter=106 channel=124
    3, -2, 3, -12, 1, -10, -3, -10, -6,
    -- layer=1 filter=106 channel=125
    25, 63, 41, -23, 32, 68, -94, -36, -37,
    -- layer=1 filter=106 channel=126
    9, 33, 9, 36, 61, 30, -7, 4, 47,
    -- layer=1 filter=106 channel=127
    1, 6, 18, 26, 21, -9, -3, 27, 14,
    -- layer=1 filter=107 channel=0
    2, 1, 5, -7, 3, -9, -4, -2, 5,
    -- layer=1 filter=107 channel=1
    2, 0, 2, 6, 7, -1, 5, -9, -10,
    -- layer=1 filter=107 channel=2
    -4, -1, -2, -6, 6, -4, -10, -8, 5,
    -- layer=1 filter=107 channel=3
    2, 1, 3, -1, 3, 6, -3, -1, 8,
    -- layer=1 filter=107 channel=4
    8, 1, 8, 2, 0, -9, 0, -11, 2,
    -- layer=1 filter=107 channel=5
    9, -8, 0, 6, -8, -4, -10, 1, -11,
    -- layer=1 filter=107 channel=6
    -7, -7, 9, -4, 2, -4, 2, 7, -1,
    -- layer=1 filter=107 channel=7
    -10, -4, 7, 0, 0, -14, 1, -8, -8,
    -- layer=1 filter=107 channel=8
    7, -7, -2, -3, -8, 0, 7, -1, -11,
    -- layer=1 filter=107 channel=9
    8, -3, -5, -3, -5, -4, 3, -8, 1,
    -- layer=1 filter=107 channel=10
    -1, 3, 6, -4, 5, 0, -4, -6, -6,
    -- layer=1 filter=107 channel=11
    -9, 4, -5, 0, 4, 8, 3, -5, -11,
    -- layer=1 filter=107 channel=12
    -8, -2, 9, -6, -9, -3, 3, -7, 1,
    -- layer=1 filter=107 channel=13
    -1, -8, -5, -4, 3, -4, 2, -5, -2,
    -- layer=1 filter=107 channel=14
    -7, 4, 0, -6, -8, -2, -8, 7, 3,
    -- layer=1 filter=107 channel=15
    -1, -4, 7, 2, -8, -6, -3, 1, -5,
    -- layer=1 filter=107 channel=16
    7, 5, -6, -11, 5, 9, 6, -2, 6,
    -- layer=1 filter=107 channel=17
    -1, -7, -4, -11, 8, -8, 0, 0, 7,
    -- layer=1 filter=107 channel=18
    7, 2, -11, -7, 0, 5, -5, 4, -2,
    -- layer=1 filter=107 channel=19
    0, -4, -7, 1, -3, 2, 2, 0, -7,
    -- layer=1 filter=107 channel=20
    0, 3, -5, -2, 3, 0, -11, -7, -10,
    -- layer=1 filter=107 channel=21
    -13, 2, 7, -9, -11, 0, 0, -10, -6,
    -- layer=1 filter=107 channel=22
    0, 5, 0, 2, 6, 2, 0, -5, -5,
    -- layer=1 filter=107 channel=23
    -10, 6, 4, -4, 1, 4, -8, 2, 7,
    -- layer=1 filter=107 channel=24
    -1, 2, 4, -7, -7, -4, 4, -2, 4,
    -- layer=1 filter=107 channel=25
    0, -7, -10, 0, 6, 3, -9, -9, -2,
    -- layer=1 filter=107 channel=26
    -2, -7, -5, 2, -3, -3, -3, -7, 2,
    -- layer=1 filter=107 channel=27
    -2, -1, 6, -2, -4, -3, -4, 5, -3,
    -- layer=1 filter=107 channel=28
    -7, -8, 3, 0, 5, 4, 0, 1, -12,
    -- layer=1 filter=107 channel=29
    -3, 9, 4, 7, 2, 5, 10, -4, -2,
    -- layer=1 filter=107 channel=30
    0, -2, -12, -2, -6, -2, -2, -5, 5,
    -- layer=1 filter=107 channel=31
    -4, -2, -2, -7, -6, -2, 8, -1, 9,
    -- layer=1 filter=107 channel=32
    -9, 6, 4, 5, -8, -3, -5, 0, -8,
    -- layer=1 filter=107 channel=33
    -3, -8, 5, 4, -8, -2, -8, 3, -4,
    -- layer=1 filter=107 channel=34
    5, -2, 2, -3, 5, 8, -9, 5, 7,
    -- layer=1 filter=107 channel=35
    1, 0, -9, 7, -12, -5, 4, -11, -10,
    -- layer=1 filter=107 channel=36
    -11, -12, -4, -6, -8, -7, 2, -7, 6,
    -- layer=1 filter=107 channel=37
    -8, -1, -9, -1, -5, 5, -5, 4, -14,
    -- layer=1 filter=107 channel=38
    0, -8, 9, -9, 0, 0, -8, -7, -2,
    -- layer=1 filter=107 channel=39
    8, -9, 1, 2, -9, -11, 0, -8, 7,
    -- layer=1 filter=107 channel=40
    2, -6, -3, -4, -9, 7, 5, 3, -11,
    -- layer=1 filter=107 channel=41
    1, 6, -1, -5, 0, -4, -11, -10, -2,
    -- layer=1 filter=107 channel=42
    9, -7, -18, -1, 4, -14, -10, 2, -15,
    -- layer=1 filter=107 channel=43
    -9, 0, -1, 5, -9, -6, 2, -5, 6,
    -- layer=1 filter=107 channel=44
    -5, 0, 7, -8, -11, -8, -6, -5, -8,
    -- layer=1 filter=107 channel=45
    -3, -9, 4, -9, 7, -1, -10, -2, 5,
    -- layer=1 filter=107 channel=46
    3, 10, -6, -6, -4, -11, -5, 4, -4,
    -- layer=1 filter=107 channel=47
    -4, 0, -2, 6, -3, 4, -11, 6, 2,
    -- layer=1 filter=107 channel=48
    2, 3, -7, 1, -3, 8, 3, -9, 5,
    -- layer=1 filter=107 channel=49
    -3, 6, 2, -2, 0, -7, -5, 2, 9,
    -- layer=1 filter=107 channel=50
    -5, -1, -7, -5, -1, 2, 5, 0, 8,
    -- layer=1 filter=107 channel=51
    -3, -4, 4, 0, -8, 5, 6, -4, -5,
    -- layer=1 filter=107 channel=52
    -2, -3, -1, -4, 8, 3, 3, 0, 6,
    -- layer=1 filter=107 channel=53
    9, -8, 8, 7, 6, -8, -8, -11, -6,
    -- layer=1 filter=107 channel=54
    10, -1, 0, 0, 3, 4, 0, 5, 6,
    -- layer=1 filter=107 channel=55
    -8, -11, 1, 6, -5, -6, 2, 10, -7,
    -- layer=1 filter=107 channel=56
    1, 2, 1, 0, -8, -5, -7, -2, 4,
    -- layer=1 filter=107 channel=57
    8, 3, -8, -7, 0, -4, 3, 1, -2,
    -- layer=1 filter=107 channel=58
    -4, -8, -8, 7, -8, 6, 8, -7, 0,
    -- layer=1 filter=107 channel=59
    9, -6, -11, 3, 7, 3, 0, 1, 2,
    -- layer=1 filter=107 channel=60
    -3, 4, 5, -7, 6, 5, -1, -4, -7,
    -- layer=1 filter=107 channel=61
    -3, -10, -1, 9, 9, 0, 0, 11, 4,
    -- layer=1 filter=107 channel=62
    3, 0, -2, -1, 6, -3, -11, -3, 0,
    -- layer=1 filter=107 channel=63
    7, 8, -1, 3, -9, 4, 8, 7, 1,
    -- layer=1 filter=107 channel=64
    1, -12, -8, -11, -8, 1, 2, -7, -1,
    -- layer=1 filter=107 channel=65
    -4, 0, -3, -5, -1, 2, -4, 2, -3,
    -- layer=1 filter=107 channel=66
    3, -2, -8, -9, -9, -3, -11, 4, -12,
    -- layer=1 filter=107 channel=67
    -1, -2, -7, -11, -7, 7, 6, -4, 0,
    -- layer=1 filter=107 channel=68
    0, -5, -3, -7, 2, -1, 8, -7, 5,
    -- layer=1 filter=107 channel=69
    -1, -9, 5, -12, -10, -6, -5, -7, -4,
    -- layer=1 filter=107 channel=70
    -1, 0, 10, -8, -3, 0, -7, 1, 5,
    -- layer=1 filter=107 channel=71
    -1, -1, -5, 3, 0, 3, 3, 4, 0,
    -- layer=1 filter=107 channel=72
    3, -8, -8, 8, 0, 0, -9, -8, -8,
    -- layer=1 filter=107 channel=73
    -9, 4, -4, 0, -6, 0, 0, -7, 7,
    -- layer=1 filter=107 channel=74
    3, 2, -2, -7, 0, -5, -1, -2, -8,
    -- layer=1 filter=107 channel=75
    0, -9, 0, -7, 2, -8, 9, -5, 0,
    -- layer=1 filter=107 channel=76
    -7, 6, -8, -9, 0, 3, -6, -4, 7,
    -- layer=1 filter=107 channel=77
    -4, 6, 6, -10, 0, 3, -8, -10, -9,
    -- layer=1 filter=107 channel=78
    1, 1, 3, -10, -6, 8, -5, 6, 1,
    -- layer=1 filter=107 channel=79
    -4, 2, 6, -10, -11, 3, 1, -5, 5,
    -- layer=1 filter=107 channel=80
    -2, -9, 3, -1, 1, 0, -9, 4, 10,
    -- layer=1 filter=107 channel=81
    3, -7, 0, -9, 0, -2, -1, 3, 5,
    -- layer=1 filter=107 channel=82
    7, -7, 8, -9, -4, 4, 0, 5, 9,
    -- layer=1 filter=107 channel=83
    2, 0, 0, -3, -8, -8, 1, 3, 8,
    -- layer=1 filter=107 channel=84
    -10, -4, -4, 2, 5, 2, 5, 0, 5,
    -- layer=1 filter=107 channel=85
    -2, 1, 3, 8, -9, -1, 3, 6, 6,
    -- layer=1 filter=107 channel=86
    9, 0, -12, -11, -12, -4, -7, -10, -4,
    -- layer=1 filter=107 channel=87
    0, -5, -2, 6, 8, -5, 5, 0, 8,
    -- layer=1 filter=107 channel=88
    -8, -10, 1, -10, 1, -11, -8, 0, -13,
    -- layer=1 filter=107 channel=89
    1, 2, -9, -8, -6, 0, -7, -6, -3,
    -- layer=1 filter=107 channel=90
    2, 6, 7, 1, 8, -5, 7, -4, 6,
    -- layer=1 filter=107 channel=91
    -3, 4, 1, -3, -9, -5, 4, 4, -6,
    -- layer=1 filter=107 channel=92
    1, 1, -1, 1, -10, 0, 5, 3, 1,
    -- layer=1 filter=107 channel=93
    3, -6, 2, 2, 0, -3, 3, 2, -1,
    -- layer=1 filter=107 channel=94
    8, -7, 5, 4, -2, 0, -2, 7, -7,
    -- layer=1 filter=107 channel=95
    0, 2, -7, 7, -2, -8, -4, 1, 0,
    -- layer=1 filter=107 channel=96
    3, 6, -7, -8, -3, -11, 8, 6, 7,
    -- layer=1 filter=107 channel=97
    -4, -9, -1, 2, -3, -2, -8, -12, -8,
    -- layer=1 filter=107 channel=98
    -12, -11, -6, 7, 7, 12, -9, -3, 6,
    -- layer=1 filter=107 channel=99
    2, 8, 7, -4, 5, -2, -3, 0, 3,
    -- layer=1 filter=107 channel=100
    3, -1, 6, 8, 4, -1, -7, -6, 2,
    -- layer=1 filter=107 channel=101
    5, -10, -2, 0, 2, 3, -1, 8, 4,
    -- layer=1 filter=107 channel=102
    4, 3, 3, 8, -7, 3, 0, 4, -9,
    -- layer=1 filter=107 channel=103
    -8, -5, 7, -9, 2, 7, -4, 0, -3,
    -- layer=1 filter=107 channel=104
    1, 6, 0, 8, 1, -4, -5, 2, -6,
    -- layer=1 filter=107 channel=105
    -1, 8, 4, -7, -6, -6, 6, 8, 6,
    -- layer=1 filter=107 channel=106
    2, 2, -3, 0, 5, 3, 4, 0, -7,
    -- layer=1 filter=107 channel=107
    -8, -1, 3, -6, -2, 2, -6, 2, 0,
    -- layer=1 filter=107 channel=108
    6, -9, 1, -12, 1, 1, 0, 0, -6,
    -- layer=1 filter=107 channel=109
    0, 6, 1, 7, 8, 0, -4, -4, 0,
    -- layer=1 filter=107 channel=110
    -6, -2, 4, -9, -5, 1, 5, -5, 5,
    -- layer=1 filter=107 channel=111
    -2, 3, 9, 2, 5, 2, -6, 4, 7,
    -- layer=1 filter=107 channel=112
    -11, 5, 6, -7, -3, -8, -1, 8, -3,
    -- layer=1 filter=107 channel=113
    -2, 0, 10, 9, -11, 1, -9, 1, 0,
    -- layer=1 filter=107 channel=114
    -1, -8, 6, -1, 0, 3, 0, 6, 0,
    -- layer=1 filter=107 channel=115
    -11, -12, 0, -8, 0, -5, 0, 1, -4,
    -- layer=1 filter=107 channel=116
    -8, -2, 5, 7, 1, 3, -8, -6, -1,
    -- layer=1 filter=107 channel=117
    -10, -9, 9, 0, -3, -4, 8, 0, 1,
    -- layer=1 filter=107 channel=118
    -5, 4, -4, -1, 4, 4, -1, -1, 6,
    -- layer=1 filter=107 channel=119
    -10, 2, 0, 8, 3, -9, 8, 3, 5,
    -- layer=1 filter=107 channel=120
    -6, -13, -11, -2, -8, 1, -10, -4, -1,
    -- layer=1 filter=107 channel=121
    -1, -1, 6, 7, -2, 5, 3, 0, -7,
    -- layer=1 filter=107 channel=122
    5, -3, -7, -5, -3, 1, -5, -2, 1,
    -- layer=1 filter=107 channel=123
    -1, -8, 2, 7, -6, 3, 6, 0, 7,
    -- layer=1 filter=107 channel=124
    -9, 3, 4, 0, -1, 0, 5, -3, 8,
    -- layer=1 filter=107 channel=125
    6, 4, 8, -6, -3, -1, -3, -3, -7,
    -- layer=1 filter=107 channel=126
    4, 1, -6, 3, 5, -4, -5, -2, -1,
    -- layer=1 filter=107 channel=127
    -5, 8, 5, 4, 2, -7, 5, -7, -2,
    -- layer=1 filter=108 channel=0
    21, -53, -9, 11, 32, -27, -36, 1, 38,
    -- layer=1 filter=108 channel=1
    -29, 45, 0, -67, -50, 59, -8, -2, -55,
    -- layer=1 filter=108 channel=2
    -28, -37, -34, -2, -47, -58, -11, -45, -86,
    -- layer=1 filter=108 channel=3
    5, -2, 3, 6, 8, 10, -9, -5, 5,
    -- layer=1 filter=108 channel=4
    -8, -9, -18, 33, 3, 23, 0, -2, 14,
    -- layer=1 filter=108 channel=5
    1, 89, 3, -51, -13, 81, 37, -38, -84,
    -- layer=1 filter=108 channel=6
    -10, -23, 7, 19, -11, -5, -23, -45, -48,
    -- layer=1 filter=108 channel=7
    -34, -90, 48, 71, 29, -51, -5, 52, 28,
    -- layer=1 filter=108 channel=8
    26, 62, -17, -63, -5, 63, 27, -37, -32,
    -- layer=1 filter=108 channel=9
    51, -37, 9, -6, 24, -45, 0, -77, 0,
    -- layer=1 filter=108 channel=10
    -11, -102, 23, 71, 49, -53, -7, 41, 71,
    -- layer=1 filter=108 channel=11
    -13, -33, -18, 4, 0, -4, -10, -15, 31,
    -- layer=1 filter=108 channel=12
    -67, 9, 23, 6, -4, -63, 2, 25, -7,
    -- layer=1 filter=108 channel=13
    38, 37, -50, -20, 23, 43, 15, -44, -15,
    -- layer=1 filter=108 channel=14
    -46, 10, 45, 104, 88, -22, 31, 56, -3,
    -- layer=1 filter=108 channel=15
    -4, 164, -7, -2, 28, 163, 14, -22, 2,
    -- layer=1 filter=108 channel=16
    22, 59, -2, -67, -9, 45, 37, -42, -61,
    -- layer=1 filter=108 channel=17
    36, -23, -86, -21, 54, 6, -30, -45, 23,
    -- layer=1 filter=108 channel=18
    11, -48, 28, 28, 35, -19, 9, 42, 17,
    -- layer=1 filter=108 channel=19
    12, -29, -45, -53, -79, -77, 36, -66, -61,
    -- layer=1 filter=108 channel=20
    -16, 29, -8, -22, -23, 16, 14, -15, -43,
    -- layer=1 filter=108 channel=21
    -26, -3, 28, -5, -35, -18, 21, 15, -26,
    -- layer=1 filter=108 channel=22
    5, 41, -53, -30, 8, 45, 0, -38, -13,
    -- layer=1 filter=108 channel=23
    -54, 13, 41, 77, -41, 14, 25, 1, -35,
    -- layer=1 filter=108 channel=24
    66, 35, -73, -75, 13, 30, 24, -105, -12,
    -- layer=1 filter=108 channel=25
    -49, -77, -7, 23, -18, -73, 15, 24, -23,
    -- layer=1 filter=108 channel=26
    41, 72, -79, -42, 10, 79, 40, -101, -16,
    -- layer=1 filter=108 channel=27
    -4, 16, 52, -4, -9, -9, 36, -2, -22,
    -- layer=1 filter=108 channel=28
    -15, -87, 28, 34, 6, -42, -24, 36, 25,
    -- layer=1 filter=108 channel=29
    1, -10, 33, 6, -4, -10, 2, 17, 14,
    -- layer=1 filter=108 channel=30
    14, -45, 26, 23, 34, -47, -14, 42, 30,
    -- layer=1 filter=108 channel=31
    -42, -2, 31, 46, 19, -26, 17, 59, -2,
    -- layer=1 filter=108 channel=32
    4, 43, -44, 25, -3, 41, 32, -21, -8,
    -- layer=1 filter=108 channel=33
    4, -10, 5, 17, 23, -24, 26, -38, -19,
    -- layer=1 filter=108 channel=34
    -46, -52, -84, -32, -63, -48, -43, -71, -86,
    -- layer=1 filter=108 channel=35
    16, 30, 3, 15, 10, 17, 1, 6, 4,
    -- layer=1 filter=108 channel=36
    1, -33, -7, -10, 1, -24, -13, 1, 43,
    -- layer=1 filter=108 channel=37
    30, 58, -34, -54, -13, 63, 47, -28, -58,
    -- layer=1 filter=108 channel=38
    15, -1, 5, 6, 16, -23, 2, -8, 0,
    -- layer=1 filter=108 channel=39
    18, 42, -48, -17, -2, 52, -4, -21, -13,
    -- layer=1 filter=108 channel=40
    -24, -20, 34, 37, 56, -36, -18, 25, 0,
    -- layer=1 filter=108 channel=41
    13, -50, -47, -4, -36, -28, 21, -75, -3,
    -- layer=1 filter=108 channel=42
    -28, -14, -16, 44, -36, -67, 14, -26, -68,
    -- layer=1 filter=108 channel=43
    14, 46, -29, -64, -24, 33, 7, -21, -50,
    -- layer=1 filter=108 channel=44
    26, 84, -50, 6, 18, 74, 35, -66, 3,
    -- layer=1 filter=108 channel=45
    37, 83, -42, -54, 23, 71, 36, -72, -26,
    -- layer=1 filter=108 channel=46
    -13, 50, 61, -51, -90, -15, 46, 2, -19,
    -- layer=1 filter=108 channel=47
    -36, 29, 24, 31, -35, 13, 6, 35, -37,
    -- layer=1 filter=108 channel=48
    21, -35, -5, 15, 34, 0, -18, -7, -3,
    -- layer=1 filter=108 channel=49
    34, 15, -2, 36, -12, -24, 29, -15, -37,
    -- layer=1 filter=108 channel=50
    5, 6, -1, -25, -1, -31, -28, -39, -14,
    -- layer=1 filter=108 channel=51
    -38, -32, 26, 45, 18, -33, -10, 5, 12,
    -- layer=1 filter=108 channel=52
    13, 15, -15, 22, -6, -1, -31, -43, 7,
    -- layer=1 filter=108 channel=53
    0, -8, -12, 8, 0, -12, -1, -11, -19,
    -- layer=1 filter=108 channel=54
    -36, -72, -21, 7, -31, -68, 32, -14, -23,
    -- layer=1 filter=108 channel=55
    -1, -9, -15, -20, 18, 46, 0, -18, 9,
    -- layer=1 filter=108 channel=56
    -3, -7, 5, 31, 5, -6, -11, -4, 4,
    -- layer=1 filter=108 channel=57
    -9, -87, 29, 66, 50, -47, -11, 38, 62,
    -- layer=1 filter=108 channel=58
    -5, -86, 16, 47, -32, -84, -22, -16, -72,
    -- layer=1 filter=108 channel=59
    9, -6, -3, -1, -22, 8, -7, -15, -9,
    -- layer=1 filter=108 channel=60
    -35, -17, -55, 33, 16, -13, 12, -29, 23,
    -- layer=1 filter=108 channel=61
    8, 4, 5, 3, -1, 3, -6, -5, 3,
    -- layer=1 filter=108 channel=62
    43, 67, -48, -63, 9, 77, 36, -44, -19,
    -- layer=1 filter=108 channel=63
    -31, -54, 23, 29, -21, -48, -18, 18, 29,
    -- layer=1 filter=108 channel=64
    -16, 9, 24, 13, -24, 0, 8, 22, -17,
    -- layer=1 filter=108 channel=65
    -4, -10, 16, 12, -11, -30, -4, -3, -19,
    -- layer=1 filter=108 channel=66
    -6, -47, 0, 5, -7, -12, -12, 1, 1,
    -- layer=1 filter=108 channel=67
    12, 9, 31, 55, 31, 10, 9, 10, -14,
    -- layer=1 filter=108 channel=68
    36, 44, -75, -27, 33, 63, 22, -95, 22,
    -- layer=1 filter=108 channel=69
    17, 115, -36, -85, 3, 121, 56, -83, -30,
    -- layer=1 filter=108 channel=70
    -35, 48, 22, 38, 23, 24, -24, 20, -25,
    -- layer=1 filter=108 channel=71
    -13, 41, 27, -1, -63, 3, 36, 6, -57,
    -- layer=1 filter=108 channel=72
    -2, -88, -38, -11, -46, -25, 12, 8, -11,
    -- layer=1 filter=108 channel=73
    7, 19, -24, 0, -7, 26, -13, -7, -10,
    -- layer=1 filter=108 channel=74
    -8, 0, -50, 11, -23, -34, -8, -37, 17,
    -- layer=1 filter=108 channel=75
    -51, 59, 61, 56, 0, -44, 6, 65, 11,
    -- layer=1 filter=108 channel=76
    -15, -25, -51, 18, 25, -19, -2, -34, 7,
    -- layer=1 filter=108 channel=77
    17, -16, -25, -12, 12, -23, 2, -14, 18,
    -- layer=1 filter=108 channel=78
    -4, -29, 22, 49, 10, -17, 15, 19, 27,
    -- layer=1 filter=108 channel=79
    31, 67, -30, -75, -19, 68, 25, -56, -42,
    -- layer=1 filter=108 channel=80
    32, 12, 25, -3, 0, 17, -2, 17, -30,
    -- layer=1 filter=108 channel=81
    33, 25, -66, -30, 18, 27, 8, -53, -37,
    -- layer=1 filter=108 channel=82
    21, 15, -16, -4, 1, 11, -4, -24, -21,
    -- layer=1 filter=108 channel=83
    47, 111, -64, -60, 43, 125, 6, -81, 2,
    -- layer=1 filter=108 channel=84
    -10, -91, -45, 14, 21, -57, -12, -23, 13,
    -- layer=1 filter=108 channel=85
    34, -49, -18, 28, -39, -22, 27, -67, -18,
    -- layer=1 filter=108 channel=86
    -12, 3, 6, 2, -7, 4, 11, 28, 15,
    -- layer=1 filter=108 channel=87
    39, -77, -4, -46, -43, -95, 17, -71, -46,
    -- layer=1 filter=108 channel=88
    1, -17, -12, 1, -1, -42, 6, -12, -56,
    -- layer=1 filter=108 channel=89
    16, 18, -3, 19, -39, -2, 4, -8, -25,
    -- layer=1 filter=108 channel=90
    50, 82, -56, -32, 34, 99, 35, -99, 6,
    -- layer=1 filter=108 channel=91
    -9, -25, 1, 36, 13, -28, -12, 10, -12,
    -- layer=1 filter=108 channel=92
    -25, 47, -22, 20, -33, 43, 0, -44, -9,
    -- layer=1 filter=108 channel=93
    9, 13, -23, -18, -8, 10, -15, -30, -25,
    -- layer=1 filter=108 channel=94
    -13, -52, 18, 44, 3, -47, -31, 20, 26,
    -- layer=1 filter=108 channel=95
    -13, -33, 17, 56, 18, -60, -26, 45, 15,
    -- layer=1 filter=108 channel=96
    -25, -46, -15, -29, -8, -32, -28, -24, -19,
    -- layer=1 filter=108 channel=97
    0, -9, -27, -16, -7, 18, -23, -10, 9,
    -- layer=1 filter=108 channel=98
    49, 32, -72, -63, 23, 73, 0, -31, 14,
    -- layer=1 filter=108 channel=99
    46, -40, -17, 24, 98, 0, -33, 4, 106,
    -- layer=1 filter=108 channel=100
    -11, -7, 23, 23, -35, -41, 8, 32, 17,
    -- layer=1 filter=108 channel=101
    -2, 1, -6, 17, 2, -22, -14, 6, -24,
    -- layer=1 filter=108 channel=102
    0, -38, 1, 27, 19, -41, -31, -14, 19,
    -- layer=1 filter=108 channel=103
    15, -26, -7, 15, 17, -26, 18, -7, 15,
    -- layer=1 filter=108 channel=104
    -14, -12, 20, 51, 2, -12, 26, 3, -7,
    -- layer=1 filter=108 channel=105
    16, -73, -35, 16, 29, -34, -31, 9, 30,
    -- layer=1 filter=108 channel=106
    3, 21, -31, 23, -5, 28, -2, -26, -28,
    -- layer=1 filter=108 channel=107
    7, 5, 8, 2, 18, 8, 5, -7, 3,
    -- layer=1 filter=108 channel=108
    52, 84, -44, -15, 28, 89, 22, -75, -19,
    -- layer=1 filter=108 channel=109
    -9, -1, 6, -4, -8, -2, 4, -7, -3,
    -- layer=1 filter=108 channel=110
    -23, 5, -8, -6, 0, -17, 0, 12, -8,
    -- layer=1 filter=108 channel=111
    50, -52, 30, 15, 83, -20, -38, 21, 45,
    -- layer=1 filter=108 channel=112
    -21, -93, -37, 36, 26, -6, -41, -23, 2,
    -- layer=1 filter=108 channel=113
    -34, -15, 5, 14, 8, -17, 27, 15, -33,
    -- layer=1 filter=108 channel=114
    21, 116, 31, -24, 8, 104, 34, -16, -49,
    -- layer=1 filter=108 channel=115
    3, -51, -11, 42, 12, -44, -4, 30, 27,
    -- layer=1 filter=108 channel=116
    5, 3, 6, -3, -8, -1, -9, 0, 6,
    -- layer=1 filter=108 channel=117
    22, -102, 7, 20, 106, 23, -72, -6, 45,
    -- layer=1 filter=108 channel=118
    3, -34, 16, 14, 48, -31, -10, 0, 31,
    -- layer=1 filter=108 channel=119
    58, 45, -86, -9, 47, 62, 33, -73, 8,
    -- layer=1 filter=108 channel=120
    -5, -57, 4, 9, -2, -23, -10, 1, 12,
    -- layer=1 filter=108 channel=121
    -10, 41, 102, 36, -41, -53, 19, 74, 28,
    -- layer=1 filter=108 channel=122
    -4, -8, 8, 2, 2, 1, 3, -7, 10,
    -- layer=1 filter=108 channel=123
    -38, -9, 69, 47, -65, -69, 22, 58, -12,
    -- layer=1 filter=108 channel=124
    17, 27, -17, 8, 6, -1, -9, -8, 8,
    -- layer=1 filter=108 channel=125
    -26, -3, 16, 45, 42, 6, -32, 6, -9,
    -- layer=1 filter=108 channel=126
    73, 46, -74, -37, 74, 109, 17, -43, 48,
    -- layer=1 filter=108 channel=127
    -7, -49, -1, 45, 10, -33, 0, 22, 39,
    -- layer=1 filter=109 channel=0
    0, -5, -11, 2, -3, 1, -2, -11, 4,
    -- layer=1 filter=109 channel=1
    -15, -13, -13, -14, -4, -6, -9, -12, -14,
    -- layer=1 filter=109 channel=2
    -16, -13, -4, -9, -10, -12, -9, 0, -1,
    -- layer=1 filter=109 channel=3
    -2, -4, 9, 8, 9, 0, 3, -9, -7,
    -- layer=1 filter=109 channel=4
    -11, 1, -2, -5, 2, -9, 5, 6, -11,
    -- layer=1 filter=109 channel=5
    -13, -13, 4, 1, -12, -8, -11, -11, -12,
    -- layer=1 filter=109 channel=6
    4, 10, 7, 0, -13, -18, 2, -4, -13,
    -- layer=1 filter=109 channel=7
    3, -6, -8, 8, -9, -16, 5, 4, -17,
    -- layer=1 filter=109 channel=8
    -14, 0, -9, 2, 6, -1, -17, -4, -11,
    -- layer=1 filter=109 channel=9
    -24, -18, 3, -2, -12, -14, 12, -5, 0,
    -- layer=1 filter=109 channel=10
    -4, -4, -8, 7, -27, -24, -10, 1, -6,
    -- layer=1 filter=109 channel=11
    2, -2, 6, -16, -10, -15, -12, -10, -11,
    -- layer=1 filter=109 channel=12
    0, 16, 10, 1, -12, -15, 1, -10, -8,
    -- layer=1 filter=109 channel=13
    3, -6, -8, -12, -9, -6, -9, -8, -16,
    -- layer=1 filter=109 channel=14
    -11, 11, -20, -7, -28, -10, 2, 3, 0,
    -- layer=1 filter=109 channel=15
    -19, -7, -7, -17, 2, -12, 0, -5, -8,
    -- layer=1 filter=109 channel=16
    -1, 3, -14, -6, 0, -2, 0, -22, -19,
    -- layer=1 filter=109 channel=17
    -8, -7, -4, 1, -14, 2, -11, -3, -11,
    -- layer=1 filter=109 channel=18
    10, 20, -1, -15, -8, -3, -4, -16, -14,
    -- layer=1 filter=109 channel=19
    -10, 3, 0, 2, -12, -3, 10, 5, 9,
    -- layer=1 filter=109 channel=20
    -5, 0, -5, -12, -16, -16, -10, -19, -16,
    -- layer=1 filter=109 channel=21
    -4, -15, -5, 0, -4, -7, -9, -8, -3,
    -- layer=1 filter=109 channel=22
    -12, -17, 1, -2, -1, -5, -25, -14, -9,
    -- layer=1 filter=109 channel=23
    -9, -5, 16, 6, 0, -3, 2, -3, -8,
    -- layer=1 filter=109 channel=24
    0, -12, -3, -6, -17, -22, -12, -1, 3,
    -- layer=1 filter=109 channel=25
    -1, -7, -3, -5, -12, -11, -15, -10, 2,
    -- layer=1 filter=109 channel=26
    -6, -11, -29, -9, -20, -28, -14, 0, -7,
    -- layer=1 filter=109 channel=27
    3, -10, 8, 10, -16, -2, 0, -1, -5,
    -- layer=1 filter=109 channel=28
    -3, -13, -9, -4, -20, -16, -4, -14, -12,
    -- layer=1 filter=109 channel=29
    6, 10, 0, -1, 8, 6, 2, -2, -2,
    -- layer=1 filter=109 channel=30
    4, -3, 14, -15, -10, -19, 6, 4, -20,
    -- layer=1 filter=109 channel=31
    6, -6, 3, -17, -25, -15, -11, 7, -6,
    -- layer=1 filter=109 channel=32
    -1, -24, -20, -18, -22, -12, -5, 0, -3,
    -- layer=1 filter=109 channel=33
    7, 1, -6, -9, -1, -5, -4, 0, 9,
    -- layer=1 filter=109 channel=34
    6, 0, 6, -4, -11, -3, 0, -10, 8,
    -- layer=1 filter=109 channel=35
    -7, -3, -10, -5, 6, -2, -1, 0, 4,
    -- layer=1 filter=109 channel=36
    -19, -3, -3, -14, 0, -6, -2, -13, -2,
    -- layer=1 filter=109 channel=37
    5, -4, -2, 4, -9, -4, -7, -5, -13,
    -- layer=1 filter=109 channel=38
    -19, -14, -13, -14, -16, -4, -21, -10, -2,
    -- layer=1 filter=109 channel=39
    -1, -12, -11, 2, 8, -1, -10, -5, 7,
    -- layer=1 filter=109 channel=40
    4, 15, -11, -14, -17, -6, -11, 4, -3,
    -- layer=1 filter=109 channel=41
    -22, -17, -11, -9, -14, -9, 3, -15, 12,
    -- layer=1 filter=109 channel=42
    1, -22, -1, -16, -17, -4, -4, -12, -4,
    -- layer=1 filter=109 channel=43
    2, -5, -2, 6, 1, 0, -8, 4, -13,
    -- layer=1 filter=109 channel=44
    -8, -12, -10, -7, -14, -23, -7, -17, -17,
    -- layer=1 filter=109 channel=45
    -15, -7, -6, -6, -12, -17, -20, -17, -6,
    -- layer=1 filter=109 channel=46
    0, 17, 10, 11, 0, -11, 9, 22, 16,
    -- layer=1 filter=109 channel=47
    6, -5, -5, -15, -10, -10, -14, -2, -6,
    -- layer=1 filter=109 channel=48
    -9, -3, -13, -19, -8, -4, -1, -14, -2,
    -- layer=1 filter=109 channel=49
    -17, -19, -19, -13, -5, -25, 2, -13, -8,
    -- layer=1 filter=109 channel=50
    7, -6, 2, -8, 0, -1, -4, -6, -11,
    -- layer=1 filter=109 channel=51
    -10, -17, -14, -13, -11, -7, -13, -4, -14,
    -- layer=1 filter=109 channel=52
    -5, 7, 4, 11, 7, 0, -2, -1, 8,
    -- layer=1 filter=109 channel=53
    -3, -7, 3, -7, 0, -4, 4, -8, 4,
    -- layer=1 filter=109 channel=54
    -3, 0, 1, -12, -11, -2, -11, 7, -7,
    -- layer=1 filter=109 channel=55
    -15, -14, -13, -7, -14, -14, -9, 1, -19,
    -- layer=1 filter=109 channel=56
    6, -5, 0, 2, -1, -4, 3, 6, 1,
    -- layer=1 filter=109 channel=57
    5, 0, -8, -12, -20, -9, -18, -6, -8,
    -- layer=1 filter=109 channel=58
    11, -12, 0, 1, -6, -10, -2, -6, -16,
    -- layer=1 filter=109 channel=59
    2, 2, -2, 3, -10, 5, 2, -7, -12,
    -- layer=1 filter=109 channel=60
    -2, -7, 7, 4, 5, 2, -11, -2, 10,
    -- layer=1 filter=109 channel=61
    0, -3, 2, 5, 7, -3, 0, 0, 3,
    -- layer=1 filter=109 channel=62
    -1, -8, -10, 6, -8, -9, -24, 0, -8,
    -- layer=1 filter=109 channel=63
    -8, -9, -7, -8, -7, -16, -11, -11, -15,
    -- layer=1 filter=109 channel=64
    2, -12, 0, 0, 2, -2, -20, -9, -14,
    -- layer=1 filter=109 channel=65
    -10, -14, -7, -13, -15, -8, -5, -7, -4,
    -- layer=1 filter=109 channel=66
    -19, -9, -2, -5, -3, -7, -6, -2, -4,
    -- layer=1 filter=109 channel=67
    7, 4, 15, 10, 7, 8, 12, 6, 5,
    -- layer=1 filter=109 channel=68
    -18, -5, -15, -13, -9, -8, -7, -23, -8,
    -- layer=1 filter=109 channel=69
    -15, 0, -5, 5, -1, -8, -12, -11, -10,
    -- layer=1 filter=109 channel=70
    1, 12, 5, 10, 0, 4, 5, -9, -5,
    -- layer=1 filter=109 channel=71
    -15, -19, -17, -7, -16, -19, -9, 0, 2,
    -- layer=1 filter=109 channel=72
    -17, -13, -4, 6, 1, -5, 5, -4, 1,
    -- layer=1 filter=109 channel=73
    -1, -5, 4, 6, -8, -2, 9, 4, -2,
    -- layer=1 filter=109 channel=74
    1, 3, 4, -6, 2, 2, -13, -17, -7,
    -- layer=1 filter=109 channel=75
    0, 8, 11, 0, -29, -3, 12, 8, -13,
    -- layer=1 filter=109 channel=76
    -17, -13, 0, 0, -22, -20, -16, -14, -10,
    -- layer=1 filter=109 channel=77
    -16, -7, -6, -7, 1, -7, 1, -6, 1,
    -- layer=1 filter=109 channel=78
    -8, -7, -9, 6, -12, -7, 8, -5, 4,
    -- layer=1 filter=109 channel=79
    -6, -9, 4, -9, -12, -11, -3, -19, -12,
    -- layer=1 filter=109 channel=80
    -1, -5, -9, -9, -1, 10, -3, 0, 4,
    -- layer=1 filter=109 channel=81
    -16, -2, -2, 1, -17, 2, 0, -5, -3,
    -- layer=1 filter=109 channel=82
    -19, -4, -15, -16, -8, -4, -8, -1, -17,
    -- layer=1 filter=109 channel=83
    -3, -8, -8, -1, 6, 9, -3, -3, -12,
    -- layer=1 filter=109 channel=84
    4, -4, -1, -6, -23, -6, 6, -4, -12,
    -- layer=1 filter=109 channel=85
    -12, -5, 1, 3, -1, -7, -15, -10, -8,
    -- layer=1 filter=109 channel=86
    -5, -8, -8, -4, -6, -11, -4, -11, -11,
    -- layer=1 filter=109 channel=87
    -16, -13, -1, -7, -10, -11, 9, 7, -3,
    -- layer=1 filter=109 channel=88
    -8, -5, -13, -4, 0, -17, 1, -5, -18,
    -- layer=1 filter=109 channel=89
    -2, -12, -20, -16, -12, -2, 1, -20, -15,
    -- layer=1 filter=109 channel=90
    -17, -8, -7, -2, -16, -11, -4, -10, -16,
    -- layer=1 filter=109 channel=91
    -7, -16, -4, -4, -7, -1, -1, -6, -2,
    -- layer=1 filter=109 channel=92
    -9, -16, -4, 0, -5, 0, -20, -10, 3,
    -- layer=1 filter=109 channel=93
    -14, -6, -13, -6, -11, -12, 0, -8, -8,
    -- layer=1 filter=109 channel=94
    -10, 6, 2, -21, -3, -13, 2, -8, -11,
    -- layer=1 filter=109 channel=95
    -5, 10, 5, -1, -17, -14, 7, -20, -15,
    -- layer=1 filter=109 channel=96
    -8, -4, 0, -6, -12, 4, -6, -3, 7,
    -- layer=1 filter=109 channel=97
    -13, -2, -7, -11, -1, -13, -10, -13, -5,
    -- layer=1 filter=109 channel=98
    -12, -4, 0, 11, -6, -1, -21, -11, -16,
    -- layer=1 filter=109 channel=99
    -10, 0, -9, -8, -9, 1, -13, 1, -7,
    -- layer=1 filter=109 channel=100
    -4, -11, 9, -7, -1, -6, -8, 1, 3,
    -- layer=1 filter=109 channel=101
    -1, -10, -9, -3, -19, -19, -6, -18, -1,
    -- layer=1 filter=109 channel=102
    0, -7, -6, -6, -16, -11, 4, -8, -9,
    -- layer=1 filter=109 channel=103
    13, 0, 15, -11, -10, -14, -4, -7, -8,
    -- layer=1 filter=109 channel=104
    -8, -11, -5, -7, 0, 3, -7, 0, -7,
    -- layer=1 filter=109 channel=105
    -21, -9, -3, -9, -13, -12, -4, -3, -3,
    -- layer=1 filter=109 channel=106
    -12, -5, -20, -6, -16, -14, -15, -13, -7,
    -- layer=1 filter=109 channel=107
    -6, 3, 11, 0, 10, -9, -7, 5, 0,
    -- layer=1 filter=109 channel=108
    -17, -12, -14, -4, -11, -15, -23, 7, -25,
    -- layer=1 filter=109 channel=109
    4, 8, 4, -5, -7, -6, 8, 2, -11,
    -- layer=1 filter=109 channel=110
    -8, 7, -7, -9, -5, -9, -2, -9, -6,
    -- layer=1 filter=109 channel=111
    -5, 7, -3, -5, -15, -6, 7, -13, -14,
    -- layer=1 filter=109 channel=112
    4, 0, -7, -16, -22, -21, -8, -5, -15,
    -- layer=1 filter=109 channel=113
    -1, -1, 0, -14, -4, -20, 1, -14, -13,
    -- layer=1 filter=109 channel=114
    -1, -2, -12, -3, -2, -5, -20, -15, 1,
    -- layer=1 filter=109 channel=115
    0, -4, -7, -13, -4, -5, 0, -6, 0,
    -- layer=1 filter=109 channel=116
    0, 2, -6, 8, -8, -7, -2, -3, 6,
    -- layer=1 filter=109 channel=117
    8, 6, 3, -1, -15, -20, -13, -17, -10,
    -- layer=1 filter=109 channel=118
    -8, 5, -5, -15, -18, -12, -14, -3, -18,
    -- layer=1 filter=109 channel=119
    -13, -9, -13, -16, -4, -14, -16, -4, -16,
    -- layer=1 filter=109 channel=120
    2, -16, 1, -17, -9, -13, -13, -4, -2,
    -- layer=1 filter=109 channel=121
    16, -1, 8, -4, -17, -3, 0, 10, 3,
    -- layer=1 filter=109 channel=122
    -5, -2, 5, -3, 2, 7, 9, -4, -9,
    -- layer=1 filter=109 channel=123
    -3, 2, -17, -12, -10, -5, -4, -7, -8,
    -- layer=1 filter=109 channel=124
    -2, -6, -8, -1, 0, 9, 4, -10, -10,
    -- layer=1 filter=109 channel=125
    0, 9, 1, 3, 1, 6, -7, -4, -9,
    -- layer=1 filter=109 channel=126
    -16, -3, -11, 5, 8, 18, -6, -11, -8,
    -- layer=1 filter=109 channel=127
    6, 13, 5, -17, -25, -1, 0, 0, -13,
    -- layer=1 filter=110 channel=0
    0, -9, -10, -2, -21, 3, 2, -11, 5,
    -- layer=1 filter=110 channel=1
    -23, -26, -30, -3, -31, -13, -2, -8, -10,
    -- layer=1 filter=110 channel=2
    -8, -8, -10, 1, -16, -11, -17, 0, -29,
    -- layer=1 filter=110 channel=3
    -7, 4, 0, 7, -11, -3, 1, -7, -14,
    -- layer=1 filter=110 channel=4
    2, -4, 2, -5, -11, -6, -2, 2, 9,
    -- layer=1 filter=110 channel=5
    -5, -30, -27, -26, -37, -31, -28, -38, -37,
    -- layer=1 filter=110 channel=6
    20, -26, 6, 7, -19, -11, -11, -40, 4,
    -- layer=1 filter=110 channel=7
    53, -24, 28, 43, 3, 30, 41, -36, 39,
    -- layer=1 filter=110 channel=8
    -29, -45, -47, -29, -45, -20, -26, -22, -25,
    -- layer=1 filter=110 channel=9
    -1, -5, 0, -18, -5, -10, -3, 21, 6,
    -- layer=1 filter=110 channel=10
    59, -19, 36, 58, -12, 53, 20, -53, 51,
    -- layer=1 filter=110 channel=11
    13, 8, 8, -10, 10, -9, 0, 8, -6,
    -- layer=1 filter=110 channel=12
    -88, -89, -32, -38, -56, -30, 25, 36, 14,
    -- layer=1 filter=110 channel=13
    -9, 30, -20, -5, 22, -26, -9, 11, -8,
    -- layer=1 filter=110 channel=14
    46, -74, -8, 14, -25, -38, 31, -34, 24,
    -- layer=1 filter=110 channel=15
    -42, 0, -46, 5, -10, -60, -3, -36, -93,
    -- layer=1 filter=110 channel=16
    7, -40, -28, -4, -47, 1, 2, -27, -19,
    -- layer=1 filter=110 channel=17
    -4, 5, -12, -13, 11, 1, -2, -10, -7,
    -- layer=1 filter=110 channel=18
    0, -24, -30, -55, -80, -59, -6, -11, -10,
    -- layer=1 filter=110 channel=19
    7, -41, -23, -27, -45, -26, -25, -48, -52,
    -- layer=1 filter=110 channel=20
    -11, 19, 6, 8, 10, -16, -4, -12, -18,
    -- layer=1 filter=110 channel=21
    -5, -19, -6, 7, -22, 14, 1, -11, 9,
    -- layer=1 filter=110 channel=22
    -10, -6, 6, -7, -28, 0, -7, -4, 4,
    -- layer=1 filter=110 channel=23
    63, 117, 0, 104, 129, 17, 97, 77, 37,
    -- layer=1 filter=110 channel=24
    1, 26, -5, -4, 29, 9, -8, 45, 2,
    -- layer=1 filter=110 channel=25
    43, -12, 10, 57, -19, 32, 33, -25, 15,
    -- layer=1 filter=110 channel=26
    -41, 44, -39, -29, 61, -45, -7, 30, -50,
    -- layer=1 filter=110 channel=27
    -9, -18, -18, 3, -12, -6, 0, -8, -4,
    -- layer=1 filter=110 channel=28
    21, -56, 29, 29, -32, 38, 32, -37, 33,
    -- layer=1 filter=110 channel=29
    -14, -30, -38, -6, -21, -14, 9, -6, -13,
    -- layer=1 filter=110 channel=30
    7, -31, -45, -85, -74, -88, -33, -34, -21,
    -- layer=1 filter=110 channel=31
    -19, -52, -13, -31, -56, -57, -38, -41, -28,
    -- layer=1 filter=110 channel=32
    -13, 75, -32, 2, 66, -66, -22, 53, -44,
    -- layer=1 filter=110 channel=33
    -12, -1, 1, -6, 0, -2, 9, -1, -20,
    -- layer=1 filter=110 channel=34
    26, 37, 24, 36, 55, 38, 36, 33, 27,
    -- layer=1 filter=110 channel=35
    -19, -8, -9, -12, -6, -3, -17, -14, -6,
    -- layer=1 filter=110 channel=36
    6, 18, 10, 11, 12, 3, 4, 6, -8,
    -- layer=1 filter=110 channel=37
    -21, -68, -23, -27, -69, -12, -24, -55, -52,
    -- layer=1 filter=110 channel=38
    -5, -1, 3, -15, -11, 11, -7, -12, 6,
    -- layer=1 filter=110 channel=39
    -11, -17, -18, -1, -8, -1, -11, -13, -13,
    -- layer=1 filter=110 channel=40
    -20, -55, -12, -56, -49, -61, -28, -63, -14,
    -- layer=1 filter=110 channel=41
    -2, 35, -24, 22, 47, -14, 3, 10, -9,
    -- layer=1 filter=110 channel=42
    -12, -12, -29, 2, -5, -4, -3, -24, -30,
    -- layer=1 filter=110 channel=43
    0, -38, 2, 30, -31, 23, 14, -22, 12,
    -- layer=1 filter=110 channel=44
    -37, 71, -65, -8, 61, -63, -28, 50, -71,
    -- layer=1 filter=110 channel=45
    -7, 19, -5, 6, 11, -26, 0, 10, 8,
    -- layer=1 filter=110 channel=46
    15, -18, -38, -15, -38, -40, -8, -50, -65,
    -- layer=1 filter=110 channel=47
    61, 102, 11, 73, 76, -11, 41, 48, -2,
    -- layer=1 filter=110 channel=48
    15, -12, -9, 12, -16, -4, 7, -11, 4,
    -- layer=1 filter=110 channel=49
    25, 13, 11, -2, 10, 0, 2, 1, 0,
    -- layer=1 filter=110 channel=50
    -18, 22, -41, -19, -14, 1, -2, -16, -11,
    -- layer=1 filter=110 channel=51
    8, -31, 6, 8, -42, 5, 11, -45, 12,
    -- layer=1 filter=110 channel=52
    12, 18, 16, -6, 6, 0, 6, 13, 2,
    -- layer=1 filter=110 channel=53
    2, 18, 9, 17, 8, 7, 13, 3, 4,
    -- layer=1 filter=110 channel=54
    15, -22, 7, 26, -40, 36, 17, -36, 2,
    -- layer=1 filter=110 channel=55
    3, 7, 0, 12, 33, 7, 4, 24, 2,
    -- layer=1 filter=110 channel=56
    -2, 4, 1, 2, 9, -2, 3, 0, 2,
    -- layer=1 filter=110 channel=57
    32, -21, 3, 20, -38, 22, 26, -55, 35,
    -- layer=1 filter=110 channel=58
    107, 140, 33, 109, 107, 40, 87, 43, 55,
    -- layer=1 filter=110 channel=59
    -18, -5, -12, -8, -10, -4, -19, 4, -12,
    -- layer=1 filter=110 channel=60
    -17, -6, -9, -10, -1, -5, -12, -1, -20,
    -- layer=1 filter=110 channel=61
    -1, -9, -4, -7, 4, 5, 3, 6, -5,
    -- layer=1 filter=110 channel=62
    -34, -78, -29, -9, -49, -10, -2, -23, -33,
    -- layer=1 filter=110 channel=63
    8, 9, -5, 6, 5, 0, 19, 7, -8,
    -- layer=1 filter=110 channel=64
    3, -18, 8, 1, -16, -9, -4, 2, 13,
    -- layer=1 filter=110 channel=65
    -2, -28, 2, 8, -25, 2, 16, 0, 9,
    -- layer=1 filter=110 channel=66
    2, 3, 4, 16, 3, -4, 9, -5, 3,
    -- layer=1 filter=110 channel=67
    1, -30, -41, -28, -42, -30, 6, -39, -37,
    -- layer=1 filter=110 channel=68
    -22, 65, -44, -22, 61, -27, -21, 62, -47,
    -- layer=1 filter=110 channel=69
    -41, 18, -3, 4, 14, -12, 10, 10, -19,
    -- layer=1 filter=110 channel=70
    20, 2, 2, 24, 15, -6, 15, -1, 12,
    -- layer=1 filter=110 channel=71
    0, -21, 13, 25, -10, 12, 18, -1, 15,
    -- layer=1 filter=110 channel=72
    14, -24, -25, -68, -57, -40, -6, -47, 8,
    -- layer=1 filter=110 channel=73
    -5, 1, 0, -9, 5, 5, 9, -6, 5,
    -- layer=1 filter=110 channel=74
    -14, 29, 27, -26, 8, 48, -14, 55, 7,
    -- layer=1 filter=110 channel=75
    -4, -31, -32, -28, -38, -73, -2, -40, -29,
    -- layer=1 filter=110 channel=76
    0, 27, -28, -5, 10, -29, -7, 32, -27,
    -- layer=1 filter=110 channel=77
    2, -17, -20, -4, 3, 10, 0, 7, 0,
    -- layer=1 filter=110 channel=78
    -1, -22, -8, -2, -1, -10, -9, 7, -17,
    -- layer=1 filter=110 channel=79
    10, -17, -11, 13, -13, 1, 23, 5, -12,
    -- layer=1 filter=110 channel=80
    -13, -12, -2, 2, -19, -11, -3, -2, -1,
    -- layer=1 filter=110 channel=81
    -2, -23, -13, 11, -11, 13, 22, 10, 26,
    -- layer=1 filter=110 channel=82
    -7, -18, -2, 8, -6, 0, 0, -5, -4,
    -- layer=1 filter=110 channel=83
    -3, 6, -32, -3, 8, -3, 4, -11, -25,
    -- layer=1 filter=110 channel=84
    -28, 3, -56, -56, -30, -94, -26, 30, -42,
    -- layer=1 filter=110 channel=85
    60, 116, 3, 107, 112, 4, 92, 53, 30,
    -- layer=1 filter=110 channel=86
    15, 11, 7, 8, -5, 4, -16, -16, -12,
    -- layer=1 filter=110 channel=87
    -9, -41, -5, -54, -33, -7, -14, -61, -51,
    -- layer=1 filter=110 channel=88
    13, -19, 0, -4, 0, -5, 0, -4, 2,
    -- layer=1 filter=110 channel=89
    -17, -12, -14, -7, 8, -12, 10, -6, -5,
    -- layer=1 filter=110 channel=90
    -29, 47, -43, -10, 72, -26, -10, 48, -46,
    -- layer=1 filter=110 channel=91
    11, -10, -7, -6, -36, -5, -2, -29, -8,
    -- layer=1 filter=110 channel=92
    -42, -3, -59, -4, 9, -86, -9, -20, -112,
    -- layer=1 filter=110 channel=93
    7, 1, -7, 9, 7, 21, 23, 12, 6,
    -- layer=1 filter=110 channel=94
    3, -25, -1, 2, -23, -4, 0, -21, 12,
    -- layer=1 filter=110 channel=95
    -8, -17, -29, -56, -60, -52, -8, 0, -13,
    -- layer=1 filter=110 channel=96
    -5, -7, -9, 12, 1, 1, -12, -1, 6,
    -- layer=1 filter=110 channel=97
    -10, -10, -5, 0, -4, 14, 2, 4, 12,
    -- layer=1 filter=110 channel=98
    -22, -54, -6, -2, -52, 19, 9, -16, 2,
    -- layer=1 filter=110 channel=99
    35, 5, 65, 17, 66, 91, 26, 53, 85,
    -- layer=1 filter=110 channel=100
    4, 13, -9, 5, 8, -8, 10, -1, -3,
    -- layer=1 filter=110 channel=101
    -3, -1, -1, 0, -13, -8, 10, 0, -4,
    -- layer=1 filter=110 channel=102
    3, -10, 12, -15, -24, 4, -14, -16, 0,
    -- layer=1 filter=110 channel=103
    -20, -20, -15, -15, -22, -24, 7, -4, -12,
    -- layer=1 filter=110 channel=104
    20, 78, -32, 62, 45, 0, 63, 9, 25,
    -- layer=1 filter=110 channel=105
    4, -25, 3, -3, -10, 20, 0, -12, 22,
    -- layer=1 filter=110 channel=106
    -14, 26, -23, -15, 25, -40, -15, 23, -25,
    -- layer=1 filter=110 channel=107
    19, 5, 18, 13, 14, 16, 14, 7, 18,
    -- layer=1 filter=110 channel=108
    -12, 66, -47, 0, 64, -50, -7, 49, -38,
    -- layer=1 filter=110 channel=109
    6, -1, 2, -3, 1, -3, 8, 2, -8,
    -- layer=1 filter=110 channel=110
    -7, -10, 3, -6, 8, -3, -2, -9, 7,
    -- layer=1 filter=110 channel=111
    11, -24, -40, -80, -104, -66, 2, -2, -14,
    -- layer=1 filter=110 channel=112
    -15, -38, -39, -15, -60, -35, 29, 35, 9,
    -- layer=1 filter=110 channel=113
    -17, -18, -12, 0, -20, -3, 0, -20, -12,
    -- layer=1 filter=110 channel=114
    -29, -49, -45, 1, -45, -43, -28, -37, -29,
    -- layer=1 filter=110 channel=115
    21, -7, 14, 28, -9, 2, 7, -16, 7,
    -- layer=1 filter=110 channel=116
    -1, -4, -4, -1, -4, 3, -11, -5, 0,
    -- layer=1 filter=110 channel=117
    -12, -64, -89, -48, -88, -74, 30, 29, 2,
    -- layer=1 filter=110 channel=118
    6, 21, -30, -51, -17, -41, 0, 19, -33,
    -- layer=1 filter=110 channel=119
    -11, 63, -43, -6, 76, -52, -2, 57, -51,
    -- layer=1 filter=110 channel=120
    17, -4, -1, 13, -14, 13, 8, -10, 7,
    -- layer=1 filter=110 channel=121
    27, -12, -8, -22, -7, -8, -9, -5, -10,
    -- layer=1 filter=110 channel=122
    -9, 10, 0, 0, -3, -8, 3, -5, -9,
    -- layer=1 filter=110 channel=123
    25, 3, 5, 6, -3, -6, 21, -16, 6,
    -- layer=1 filter=110 channel=124
    -9, 3, 2, -10, -3, -9, -13, -3, -8,
    -- layer=1 filter=110 channel=125
    -3, -8, 4, -22, 8, 13, -19, -37, 9,
    -- layer=1 filter=110 channel=126
    -82, -99, -62, -50, -50, -36, -27, -20, -45,
    -- layer=1 filter=110 channel=127
    0, -3, -27, -70, -69, -56, -15, -11, -20,
    -- layer=1 filter=111 channel=0
    -13, -5, -2, -7, -6, 2, -3, -2, 0,
    -- layer=1 filter=111 channel=1
    3, 0, 0, -8, -11, -7, -8, 1, 0,
    -- layer=1 filter=111 channel=2
    5, -13, 0, -2, -2, -9, -7, -11, -7,
    -- layer=1 filter=111 channel=3
    8, 4, -1, 9, 6, 10, 0, -5, 6,
    -- layer=1 filter=111 channel=4
    2, 3, -8, -5, -8, -3, -3, -7, 0,
    -- layer=1 filter=111 channel=5
    3, -7, 2, -10, 0, 0, -16, -8, 2,
    -- layer=1 filter=111 channel=6
    -7, -18, 3, 2, -1, -7, -13, -15, -7,
    -- layer=1 filter=111 channel=7
    -4, -11, -14, 8, 2, -7, 0, -14, -7,
    -- layer=1 filter=111 channel=8
    -7, -4, 2, -5, -2, -1, -10, -2, -6,
    -- layer=1 filter=111 channel=9
    8, -7, -12, -6, 5, -3, -8, -2, 7,
    -- layer=1 filter=111 channel=10
    0, 2, -3, 7, 4, -1, 0, -16, -6,
    -- layer=1 filter=111 channel=11
    0, -15, 0, -2, 0, -3, 0, 4, -11,
    -- layer=1 filter=111 channel=12
    3, 0, 5, 5, -6, 4, -10, -7, 8,
    -- layer=1 filter=111 channel=13
    -15, -5, 4, -15, -12, -6, -17, -13, -10,
    -- layer=1 filter=111 channel=14
    -18, -8, 0, -13, 2, -2, -4, 4, 1,
    -- layer=1 filter=111 channel=15
    0, 0, -5, 4, 7, 2, 5, -2, -2,
    -- layer=1 filter=111 channel=16
    -2, -5, -13, -9, -9, -16, 2, -3, -3,
    -- layer=1 filter=111 channel=17
    -11, 1, 2, -8, 2, -14, -11, -9, -8,
    -- layer=1 filter=111 channel=18
    1, -1, -9, -12, -12, -7, 0, -2, -8,
    -- layer=1 filter=111 channel=19
    -1, -8, -5, -5, -6, 0, 6, 0, -9,
    -- layer=1 filter=111 channel=20
    -7, 3, 0, 4, -14, 1, 3, -6, 3,
    -- layer=1 filter=111 channel=21
    -4, -9, 1, -2, -9, 4, -13, -8, 5,
    -- layer=1 filter=111 channel=22
    -8, -3, -1, -14, -1, 5, -8, -9, 1,
    -- layer=1 filter=111 channel=23
    -2, 7, -5, -8, 0, -7, 2, -1, 2,
    -- layer=1 filter=111 channel=24
    -11, -1, 3, -10, 1, -1, -3, -6, 0,
    -- layer=1 filter=111 channel=25
    -6, -9, -1, -10, -4, -3, 3, -3, 4,
    -- layer=1 filter=111 channel=26
    -14, -3, -15, -3, -5, 1, -10, 4, -17,
    -- layer=1 filter=111 channel=27
    -16, -12, -4, -5, 0, 0, -14, -2, -15,
    -- layer=1 filter=111 channel=28
    -11, -3, -8, 4, -5, -1, -11, -9, 6,
    -- layer=1 filter=111 channel=29
    0, 8, -4, -12, -1, 7, -8, -9, -11,
    -- layer=1 filter=111 channel=30
    -14, -7, -14, 9, 2, -5, -7, -14, -11,
    -- layer=1 filter=111 channel=31
    0, 5, 5, -18, -11, -8, -5, 4, 2,
    -- layer=1 filter=111 channel=32
    -15, -4, -3, -13, -9, -16, 0, 5, -5,
    -- layer=1 filter=111 channel=33
    4, -8, -10, 3, 0, -14, -9, -10, -4,
    -- layer=1 filter=111 channel=34
    -12, 4, -11, 1, 0, -1, -4, 7, -4,
    -- layer=1 filter=111 channel=35
    -4, -3, -6, -8, 3, 4, 1, 4, -5,
    -- layer=1 filter=111 channel=36
    0, -16, -9, 5, -12, -11, 3, -11, -8,
    -- layer=1 filter=111 channel=37
    5, -10, 0, -15, 0, -5, -10, -1, -3,
    -- layer=1 filter=111 channel=38
    -13, -2, -11, -7, 0, -3, -8, -2, 1,
    -- layer=1 filter=111 channel=39
    -13, 3, -2, 3, 0, 4, -9, 7, 3,
    -- layer=1 filter=111 channel=40
    -16, -20, -5, -19, -6, 9, -6, 0, 10,
    -- layer=1 filter=111 channel=41
    -10, -5, 1, -5, 1, -5, -6, 3, -9,
    -- layer=1 filter=111 channel=42
    -10, -10, 6, 2, -6, 2, -5, -1, -11,
    -- layer=1 filter=111 channel=43
    -1, -4, -15, -9, 4, -5, -10, 6, 5,
    -- layer=1 filter=111 channel=44
    -10, 1, 1, -7, 6, -3, -13, -8, -16,
    -- layer=1 filter=111 channel=45
    -9, -5, -9, -3, -11, -14, -9, -14, -15,
    -- layer=1 filter=111 channel=46
    -1, -12, 5, 1, 3, -3, -6, 8, -5,
    -- layer=1 filter=111 channel=47
    -13, -4, 0, 0, 4, 2, -12, -2, -11,
    -- layer=1 filter=111 channel=48
    -6, -10, 0, -11, -2, -10, 0, -14, -8,
    -- layer=1 filter=111 channel=49
    -6, 0, -2, 4, -13, -14, -4, -8, 1,
    -- layer=1 filter=111 channel=50
    -11, -6, 3, -4, -11, 6, 1, 0, -7,
    -- layer=1 filter=111 channel=51
    -10, -5, 1, 1, -12, -13, -12, -11, 4,
    -- layer=1 filter=111 channel=52
    2, 0, -3, 2, 7, -6, -7, -9, 4,
    -- layer=1 filter=111 channel=53
    5, -1, 0, 7, 2, -4, 2, -2, -7,
    -- layer=1 filter=111 channel=54
    3, -4, 3, -6, -5, -12, -7, 7, -9,
    -- layer=1 filter=111 channel=55
    6, -9, -15, -1, -17, -2, -1, 2, -2,
    -- layer=1 filter=111 channel=56
    -2, -11, 3, 6, -3, -1, -11, -9, 8,
    -- layer=1 filter=111 channel=57
    -2, -7, -2, -11, -12, -5, -9, -9, 4,
    -- layer=1 filter=111 channel=58
    4, 0, -8, -7, 7, -4, 0, -9, 3,
    -- layer=1 filter=111 channel=59
    -8, -7, 0, 8, -5, 0, 2, 6, 0,
    -- layer=1 filter=111 channel=60
    -6, 1, -2, -4, 8, 0, 2, -10, 3,
    -- layer=1 filter=111 channel=61
    -8, 8, 6, 3, -2, -4, -8, 2, 2,
    -- layer=1 filter=111 channel=62
    -7, -1, -6, -18, 1, -8, -4, -11, -6,
    -- layer=1 filter=111 channel=63
    -14, -4, -11, 0, -13, -13, -9, 3, -9,
    -- layer=1 filter=111 channel=64
    -9, 3, 1, -7, 5, -6, -4, -8, 3,
    -- layer=1 filter=111 channel=65
    -11, 0, 4, 1, -7, 3, -9, 0, -3,
    -- layer=1 filter=111 channel=66
    -9, -13, -16, -8, -15, -2, 2, -12, -9,
    -- layer=1 filter=111 channel=67
    2, 5, -10, -3, -10, 0, -9, 0, 0,
    -- layer=1 filter=111 channel=68
    -2, 7, -1, -9, 1, -6, -14, -2, -15,
    -- layer=1 filter=111 channel=69
    -3, -5, -9, 0, -2, -9, -3, -5, 0,
    -- layer=1 filter=111 channel=70
    3, -6, -9, -1, -6, -14, -15, -15, 6,
    -- layer=1 filter=111 channel=71
    -8, -3, -6, -17, -10, -4, -5, -10, -14,
    -- layer=1 filter=111 channel=72
    -3, 1, -12, 0, 2, -3, -11, -2, -11,
    -- layer=1 filter=111 channel=73
    3, 8, -5, 1, 7, 9, 6, 6, -2,
    -- layer=1 filter=111 channel=74
    1, -13, -14, -2, -3, -12, -12, 0, 0,
    -- layer=1 filter=111 channel=75
    -4, 4, -13, -4, -8, 0, -8, -10, -12,
    -- layer=1 filter=111 channel=76
    -5, 0, 0, -15, -9, -4, 1, -10, 6,
    -- layer=1 filter=111 channel=77
    -11, 4, -10, -3, 4, 6, 4, 8, -11,
    -- layer=1 filter=111 channel=78
    -3, -11, -7, 0, 1, 0, -2, 2, -8,
    -- layer=1 filter=111 channel=79
    -13, -4, -15, 0, 0, 2, -1, -11, -8,
    -- layer=1 filter=111 channel=80
    2, -7, 7, -6, -6, -3, -8, -9, 0,
    -- layer=1 filter=111 channel=81
    -4, -9, -2, -3, 2, 0, 3, -11, -7,
    -- layer=1 filter=111 channel=82
    2, -8, 3, -9, -3, 2, -10, -12, -1,
    -- layer=1 filter=111 channel=83
    6, 0, -8, -11, -3, -7, -11, 0, -6,
    -- layer=1 filter=111 channel=84
    1, 0, -10, -14, -2, -12, 0, -14, -13,
    -- layer=1 filter=111 channel=85
    -3, 6, -2, -9, 3, 2, -16, 4, 6,
    -- layer=1 filter=111 channel=86
    -14, -13, -10, 4, 1, -13, 4, 3, 0,
    -- layer=1 filter=111 channel=87
    4, -3, -2, -6, -11, -10, -6, 8, 8,
    -- layer=1 filter=111 channel=88
    -5, -2, 1, -8, -4, 0, -9, 0, 2,
    -- layer=1 filter=111 channel=89
    -11, -10, -5, -17, -3, -14, -5, -6, 0,
    -- layer=1 filter=111 channel=90
    5, -6, -7, 6, -13, -6, 0, -1, 1,
    -- layer=1 filter=111 channel=91
    -5, -13, 4, -12, -9, 1, -10, 0, 4,
    -- layer=1 filter=111 channel=92
    7, -5, -9, 1, -2, 2, -6, -1, 1,
    -- layer=1 filter=111 channel=93
    -9, -16, -3, 0, 0, -14, 3, -10, -14,
    -- layer=1 filter=111 channel=94
    -4, -7, -11, 2, -10, -7, 0, -14, -3,
    -- layer=1 filter=111 channel=95
    -8, 0, 5, -14, -9, -14, -6, 0, -14,
    -- layer=1 filter=111 channel=96
    0, -4, 7, 0, -2, -7, -9, 8, -1,
    -- layer=1 filter=111 channel=97
    -1, 0, -6, -13, 0, -15, -6, -5, 0,
    -- layer=1 filter=111 channel=98
    4, 7, 1, -6, -16, 2, 0, 4, -3,
    -- layer=1 filter=111 channel=99
    -13, 3, 2, -12, -1, -4, 0, 6, -4,
    -- layer=1 filter=111 channel=100
    -4, -4, -10, -2, -6, -3, 6, -5, -12,
    -- layer=1 filter=111 channel=101
    -15, -10, -15, -9, -14, -3, 0, 0, 0,
    -- layer=1 filter=111 channel=102
    1, -12, 0, 2, -11, -2, 1, 5, -12,
    -- layer=1 filter=111 channel=103
    -3, -2, -2, -15, -3, -5, 1, 2, -11,
    -- layer=1 filter=111 channel=104
    3, 4, -8, 7, 2, -6, -9, -5, -10,
    -- layer=1 filter=111 channel=105
    -3, -11, -3, 0, -10, -4, 1, -15, -14,
    -- layer=1 filter=111 channel=106
    -17, -2, -16, -11, 5, -11, -21, 6, -14,
    -- layer=1 filter=111 channel=107
    6, -5, -7, 4, -6, 5, 4, -4, -2,
    -- layer=1 filter=111 channel=108
    -1, -11, -14, 0, 5, -8, 0, -4, -4,
    -- layer=1 filter=111 channel=109
    -1, -9, 0, 7, 5, -4, -4, 10, -4,
    -- layer=1 filter=111 channel=110
    -1, -5, -5, -4, 6, 5, 3, -1, 6,
    -- layer=1 filter=111 channel=111
    -2, -4, 3, 0, 5, 0, -12, -9, -7,
    -- layer=1 filter=111 channel=112
    -5, 1, 2, -3, -3, -7, -2, -2, -2,
    -- layer=1 filter=111 channel=113
    3, -10, -10, 10, 0, -6, 7, -5, 9,
    -- layer=1 filter=111 channel=114
    -13, -1, 2, -5, -17, -1, 0, -7, 0,
    -- layer=1 filter=111 channel=115
    -16, -15, -18, -10, 0, 0, -3, -2, -14,
    -- layer=1 filter=111 channel=116
    7, 5, -2, -9, 6, 0, -1, 0, -7,
    -- layer=1 filter=111 channel=117
    -3, -3, 1, -16, 5, 0, -2, -17, -13,
    -- layer=1 filter=111 channel=118
    -6, -15, -17, 0, -9, -7, -2, -4, -1,
    -- layer=1 filter=111 channel=119
    2, 7, -11, -4, 0, 3, -17, 2, -9,
    -- layer=1 filter=111 channel=120
    -4, -12, 5, -9, -3, -12, -10, -13, -11,
    -- layer=1 filter=111 channel=121
    -15, -6, -6, -5, -12, -15, -5, -11, -4,
    -- layer=1 filter=111 channel=122
    3, 3, 6, 6, 8, -6, 7, 9, -4,
    -- layer=1 filter=111 channel=123
    -1, 1, 0, 4, -7, -16, -10, 1, -14,
    -- layer=1 filter=111 channel=124
    -2, 5, 2, -9, 7, 6, -3, -6, 2,
    -- layer=1 filter=111 channel=125
    -5, 0, -7, -14, 0, 0, 0, -4, 9,
    -- layer=1 filter=111 channel=126
    -10, 8, -10, -1, 0, -5, -5, 0, 0,
    -- layer=1 filter=111 channel=127
    -7, -13, -9, -12, 0, -8, -10, -11, -19,
    -- layer=1 filter=112 channel=0
    1, -16, -11, 0, 4, 7, -19, -3, 0,
    -- layer=1 filter=112 channel=1
    23, 25, -3, -4, -18, -25, 1, 5, -1,
    -- layer=1 filter=112 channel=2
    15, 16, 8, 20, 11, 15, -12, -14, 1,
    -- layer=1 filter=112 channel=3
    0, 4, -11, -15, -9, -1, -3, 7, 9,
    -- layer=1 filter=112 channel=4
    0, -7, 6, -7, -2, 0, 3, -10, -7,
    -- layer=1 filter=112 channel=5
    38, 47, 37, -17, -4, -24, 4, 13, -9,
    -- layer=1 filter=112 channel=6
    -30, -31, -15, -58, -76, -98, -3, -2, -12,
    -- layer=1 filter=112 channel=7
    -56, -61, 0, -16, -38, -1, -19, 23, 18,
    -- layer=1 filter=112 channel=8
    39, 27, 15, -12, -11, 5, 14, 20, 18,
    -- layer=1 filter=112 channel=9
    -24, -42, 10, -13, -2, -41, 7, -7, 21,
    -- layer=1 filter=112 channel=10
    -47, -47, -3, -6, -28, -7, -18, 17, 23,
    -- layer=1 filter=112 channel=11
    5, -12, -8, 23, 22, 13, -3, 1, 4,
    -- layer=1 filter=112 channel=12
    -23, 7, -4, -2, -35, -26, -2, 24, 31,
    -- layer=1 filter=112 channel=13
    -15, -9, -15, -52, -44, -71, 4, -5, -2,
    -- layer=1 filter=112 channel=14
    -63, -31, 21, 16, 0, -5, -4, 64, 46,
    -- layer=1 filter=112 channel=15
    16, -6, 33, -4, 30, -39, 0, -9, -3,
    -- layer=1 filter=112 channel=16
    15, 7, 7, -22, -23, -24, 11, 9, 14,
    -- layer=1 filter=112 channel=17
    15, 7, 3, -20, -22, -11, -3, -5, -15,
    -- layer=1 filter=112 channel=18
    5, 21, 13, 42, 11, 13, -35, 8, 27,
    -- layer=1 filter=112 channel=19
    0, -23, 47, 20, -9, -35, 6, -11, 11,
    -- layer=1 filter=112 channel=20
    -10, 5, 3, -59, -57, -52, -14, -2, -16,
    -- layer=1 filter=112 channel=21
    -29, -15, -43, -27, -26, -42, -19, 4, -21,
    -- layer=1 filter=112 channel=22
    10, 25, 0, -2, -13, -20, 30, 32, 24,
    -- layer=1 filter=112 channel=23
    -12, -35, -3, -28, -8, -18, 20, 11, 11,
    -- layer=1 filter=112 channel=24
    -3, -14, 12, -12, -6, 1, 24, -1, 22,
    -- layer=1 filter=112 channel=25
    -7, -23, -12, -23, -73, -15, 3, -3, 13,
    -- layer=1 filter=112 channel=26
    -12, -19, 10, 2, 0, -37, 28, 20, 37,
    -- layer=1 filter=112 channel=27
    -40, -43, -59, -10, -15, -30, -13, -9, -21,
    -- layer=1 filter=112 channel=28
    -43, -26, -33, -9, -22, -18, -3, 20, 32,
    -- layer=1 filter=112 channel=29
    -57, -47, -52, -34, -41, -21, -25, -13, -5,
    -- layer=1 filter=112 channel=30
    19, 0, 18, 27, 13, -14, -25, 3, 34,
    -- layer=1 filter=112 channel=31
    -10, 6, 14, 28, -13, -18, 4, 42, 22,
    -- layer=1 filter=112 channel=32
    -3, -27, -9, -11, -21, -48, 5, -4, 44,
    -- layer=1 filter=112 channel=33
    -7, -2, 3, 9, 8, -2, 6, 18, 3,
    -- layer=1 filter=112 channel=34
    -14, 3, -3, -5, -4, 0, -14, -2, -3,
    -- layer=1 filter=112 channel=35
    -11, -2, -14, -13, -3, -11, -2, -15, -4,
    -- layer=1 filter=112 channel=36
    2, -9, -2, 28, 29, 25, 0, -3, 14,
    -- layer=1 filter=112 channel=37
    49, 23, 27, -17, -14, 0, 10, 5, -9,
    -- layer=1 filter=112 channel=38
    -22, -11, -2, -49, -59, -55, -35, -27, -37,
    -- layer=1 filter=112 channel=39
    -6, -10, -11, -9, -11, -13, 4, 8, 2,
    -- layer=1 filter=112 channel=40
    -20, -4, -26, 19, -19, -48, 11, 30, 6,
    -- layer=1 filter=112 channel=41
    -17, -42, 12, 1, 2, -44, 12, -25, 31,
    -- layer=1 filter=112 channel=42
    14, 23, 16, -5, -14, 0, -3, -24, -24,
    -- layer=1 filter=112 channel=43
    21, 12, 10, -17, -13, -12, 18, 23, 9,
    -- layer=1 filter=112 channel=44
    -18, -40, -8, 7, -21, -19, 12, 39, 29,
    -- layer=1 filter=112 channel=45
    -19, -13, 12, -18, -4, -35, -12, -12, -8,
    -- layer=1 filter=112 channel=46
    14, 17, 104, -7, 0, -11, -15, -18, -18,
    -- layer=1 filter=112 channel=47
    -23, -43, 5, -5, -20, -30, -9, -12, 15,
    -- layer=1 filter=112 channel=48
    -4, 3, -11, -16, -12, -9, -13, -12, 8,
    -- layer=1 filter=112 channel=49
    -29, -24, -8, -28, -17, -26, -21, -23, -3,
    -- layer=1 filter=112 channel=50
    4, -3, 4, -3, 7, -9, -5, -13, 15,
    -- layer=1 filter=112 channel=51
    -5, 2, -29, -2, -22, -37, -23, -6, -1,
    -- layer=1 filter=112 channel=52
    13, 21, 3, 14, 2, 17, 0, 4, 10,
    -- layer=1 filter=112 channel=53
    2, -1, 7, -8, 3, -5, 1, -7, 6,
    -- layer=1 filter=112 channel=54
    11, -12, 7, -21, -41, -11, -11, 11, -4,
    -- layer=1 filter=112 channel=55
    -2, 0, -4, 24, 28, 30, 18, 10, 14,
    -- layer=1 filter=112 channel=56
    0, 8, 4, -8, -6, 0, 3, -11, -6,
    -- layer=1 filter=112 channel=57
    -55, -60, -16, -5, -57, -30, -12, -11, 1,
    -- layer=1 filter=112 channel=58
    -52, -103, -26, -18, -71, -41, 3, -22, -9,
    -- layer=1 filter=112 channel=59
    6, 1, -5, -8, 3, 0, 5, -10, -13,
    -- layer=1 filter=112 channel=60
    -16, -4, -22, 1, -17, 0, -1, -13, -1,
    -- layer=1 filter=112 channel=61
    1, -6, 4, 8, -8, -7, 9, -4, 4,
    -- layer=1 filter=112 channel=62
    23, 16, 14, -9, -25, -4, 5, 27, 17,
    -- layer=1 filter=112 channel=63
    -2, -5, -13, 30, 20, 21, -14, 3, 13,
    -- layer=1 filter=112 channel=64
    8, -3, -10, -2, -14, -10, -2, -10, -13,
    -- layer=1 filter=112 channel=65
    -15, -8, -22, -1, -14, -26, -6, 15, -5,
    -- layer=1 filter=112 channel=66
    -10, -6, -2, -6, 15, 4, -9, 1, -8,
    -- layer=1 filter=112 channel=67
    -47, -32, -39, -57, -56, -49, -16, -11, -8,
    -- layer=1 filter=112 channel=68
    -7, -28, -18, 0, -47, -55, 24, 0, 36,
    -- layer=1 filter=112 channel=69
    34, 7, 10, -2, 16, -26, 13, 29, 19,
    -- layer=1 filter=112 channel=70
    16, 13, 36, -24, -51, -20, 14, 8, -47,
    -- layer=1 filter=112 channel=71
    -6, -15, -14, -2, 10, 6, 6, 17, 5,
    -- layer=1 filter=112 channel=72
    -16, -11, 19, 5, 0, -32, 18, -1, 28,
    -- layer=1 filter=112 channel=73
    -3, 2, 1, -3, -6, -2, 12, 10, -6,
    -- layer=1 filter=112 channel=74
    28, -3, -3, 1, -27, -30, -18, -18, 12,
    -- layer=1 filter=112 channel=75
    -1, 4, 7, 28, -8, -20, -11, 61, 48,
    -- layer=1 filter=112 channel=76
    9, -23, -17, 3, -17, -10, -20, -29, 14,
    -- layer=1 filter=112 channel=77
    1, 1, -14, -2, 7, 2, 4, 20, 15,
    -- layer=1 filter=112 channel=78
    0, 0, 14, -6, 5, -2, -2, 17, 6,
    -- layer=1 filter=112 channel=79
    31, 13, 14, -24, -24, -13, 2, 15, 7,
    -- layer=1 filter=112 channel=80
    0, 10, -7, -6, 1, 1, -2, -1, -3,
    -- layer=1 filter=112 channel=81
    -9, -18, -8, -9, -6, 0, 27, 25, 37,
    -- layer=1 filter=112 channel=82
    -17, -14, -28, -38, -30, -27, 3, -10, -20,
    -- layer=1 filter=112 channel=83
    12, 25, 21, 11, 2, -27, 0, -3, 4,
    -- layer=1 filter=112 channel=84
    16, -2, 3, 28, 0, -2, -34, -4, 21,
    -- layer=1 filter=112 channel=85
    -5, -40, -5, -22, -52, -35, 14, -23, -14,
    -- layer=1 filter=112 channel=86
    3, 3, 0, -4, 6, 7, 5, -7, 6,
    -- layer=1 filter=112 channel=87
    13, -2, 72, 21, -4, -38, -23, -22, -12,
    -- layer=1 filter=112 channel=88
    -16, -11, -16, -23, 0, -12, -11, -14, 0,
    -- layer=1 filter=112 channel=89
    -32, -29, -26, -42, -34, -39, -25, 19, -10,
    -- layer=1 filter=112 channel=90
    -22, -29, -23, -4, -24, -50, 7, 13, 26,
    -- layer=1 filter=112 channel=91
    1, -3, -18, -29, -48, -65, -15, -24, -25,
    -- layer=1 filter=112 channel=92
    -29, -67, -24, 9, 16, -34, 27, 24, 20,
    -- layer=1 filter=112 channel=93
    1, 2, 12, -11, -1, -4, 0, 6, 0,
    -- layer=1 filter=112 channel=94
    -11, -15, -6, -13, -2, 12, -26, -11, -9,
    -- layer=1 filter=112 channel=95
    22, 12, 2, 21, 2, -6, -55, 27, 19,
    -- layer=1 filter=112 channel=96
    0, -2, 1, 8, -14, 1, -5, -6, 9,
    -- layer=1 filter=112 channel=97
    4, 0, 6, 0, -2, 0, -6, -2, 5,
    -- layer=1 filter=112 channel=98
    23, 13, 20, 3, -26, -8, 28, 31, 13,
    -- layer=1 filter=112 channel=99
    -52, -42, -14, 4, -7, -12, -13, 10, 37,
    -- layer=1 filter=112 channel=100
    1, -6, -25, 27, 12, -3, -5, -10, -9,
    -- layer=1 filter=112 channel=101
    1, -1, 0, -38, -58, -52, -35, -19, -36,
    -- layer=1 filter=112 channel=102
    2, -9, -10, -12, -26, -21, -35, -17, -24,
    -- layer=1 filter=112 channel=103
    9, 8, -7, 15, 7, -1, -10, -5, 15,
    -- layer=1 filter=112 channel=104
    -16, -21, 40, -4, -2, -10, -34, -5, -4,
    -- layer=1 filter=112 channel=105
    1, 7, 9, 4, 12, 17, -11, -6, -4,
    -- layer=1 filter=112 channel=106
    -14, -10, -19, -44, -60, -39, -44, -7, -23,
    -- layer=1 filter=112 channel=107
    9, 15, 13, 3, 3, 6, 10, 1, 7,
    -- layer=1 filter=112 channel=108
    -38, -61, -7, -17, -21, -55, 12, -1, 28,
    -- layer=1 filter=112 channel=109
    2, 5, 1, 8, -6, -9, 8, 8, 6,
    -- layer=1 filter=112 channel=110
    -9, 0, 4, 0, 0, 7, -13, -9, -1,
    -- layer=1 filter=112 channel=111
    19, 13, 5, 30, 29, 5, -46, -12, 18,
    -- layer=1 filter=112 channel=112
    29, 6, 15, 30, 10, 38, -51, 6, 19,
    -- layer=1 filter=112 channel=113
    -11, -7, -2, -5, -29, -4, 6, -35, -20,
    -- layer=1 filter=112 channel=114
    15, 7, 13, -12, 3, -29, 12, 21, 2,
    -- layer=1 filter=112 channel=115
    0, 5, 0, -5, 4, 16, -2, -7, 6,
    -- layer=1 filter=112 channel=116
    5, 7, -9, 0, -11, -9, -6, -7, -4,
    -- layer=1 filter=112 channel=117
    45, 25, 41, 37, 22, 51, -9, 2, 44,
    -- layer=1 filter=112 channel=118
    20, 22, 3, 6, 4, -15, -33, -14, 14,
    -- layer=1 filter=112 channel=119
    -7, -41, -9, -19, -34, -45, 6, -24, 21,
    -- layer=1 filter=112 channel=120
    -6, -8, -23, -6, -32, -36, -21, 4, -4,
    -- layer=1 filter=112 channel=121
    -20, -23, 3, 4, 7, -9, -6, 21, 9,
    -- layer=1 filter=112 channel=122
    -6, -9, 7, 6, -9, 3, 1, 10, -5,
    -- layer=1 filter=112 channel=123
    -27, -19, -25, 14, 4, -6, -2, 17, 10,
    -- layer=1 filter=112 channel=124
    -5, 0, -9, 2, 1, 1, 6, 1, 1,
    -- layer=1 filter=112 channel=125
    32, 30, 43, -7, -39, -27, 7, 14, 1,
    -- layer=1 filter=112 channel=126
    57, 66, 37, 41, 6, 18, 41, 16, 47,
    -- layer=1 filter=112 channel=127
    28, 23, 26, 25, 30, -5, -35, 19, 21,
    -- layer=1 filter=113 channel=0
    -15, -2, -11, -4, -1, -12, -2, -3, -6,
    -- layer=1 filter=113 channel=1
    6, 0, -11, -16, -19, -20, -16, 9, -9,
    -- layer=1 filter=113 channel=2
    11, 13, 32, 20, 15, 24, -25, -11, -12,
    -- layer=1 filter=113 channel=3
    -4, -6, -1, 7, -4, -10, 1, 8, -10,
    -- layer=1 filter=113 channel=4
    -7, 10, 10, -9, 3, -3, 2, -7, -2,
    -- layer=1 filter=113 channel=5
    3, -6, -10, -1, -3, 16, 20, 16, 8,
    -- layer=1 filter=113 channel=6
    12, 38, 60, -52, -10, -19, -82, -70, -51,
    -- layer=1 filter=113 channel=7
    0, -65, -3, -74, -103, -44, -82, -106, -85,
    -- layer=1 filter=113 channel=8
    19, 0, -9, 2, -3, -33, 7, 33, 5,
    -- layer=1 filter=113 channel=9
    36, 14, 27, -20, 5, 11, -32, -25, -1,
    -- layer=1 filter=113 channel=10
    0, -45, 5, -75, -68, -26, -58, -102, -75,
    -- layer=1 filter=113 channel=11
    2, 3, 1, 21, -2, -3, 31, 12, 21,
    -- layer=1 filter=113 channel=12
    -35, -14, -13, -4, 10, 24, -37, -64, -62,
    -- layer=1 filter=113 channel=13
    20, 39, 46, -3, -11, -7, -22, -18, -20,
    -- layer=1 filter=113 channel=14
    -16, -22, 7, -57, -28, -15, -69, -31, -55,
    -- layer=1 filter=113 channel=15
    2, 18, 34, -30, -44, -39, -18, -35, -39,
    -- layer=1 filter=113 channel=16
    0, 0, -10, -9, -16, -13, 20, 5, -10,
    -- layer=1 filter=113 channel=17
    1, 0, -7, 0, -21, -16, 1, 3, -18,
    -- layer=1 filter=113 channel=18
    27, 19, 12, -13, 8, -1, -5, -18, 28,
    -- layer=1 filter=113 channel=19
    67, 24, 22, 22, -12, -8, -24, -54, -31,
    -- layer=1 filter=113 channel=20
    30, 43, 40, -8, -4, 4, -7, -9, -8,
    -- layer=1 filter=113 channel=21
    -6, 15, 25, 0, 4, 0, -13, -16, -16,
    -- layer=1 filter=113 channel=22
    25, 38, 46, -23, -18, -23, -21, -25, -34,
    -- layer=1 filter=113 channel=23
    3, -30, -25, -49, -74, -44, -32, -24, -45,
    -- layer=1 filter=113 channel=24
    6, 2, 14, 5, 13, 27, 16, 1, 12,
    -- layer=1 filter=113 channel=25
    20, -21, 12, -33, -67, -31, -10, -41, -16,
    -- layer=1 filter=113 channel=26
    39, 7, 30, -6, -36, 5, 0, -4, 0,
    -- layer=1 filter=113 channel=27
    -47, -49, -60, -19, -19, -29, -9, -3, -11,
    -- layer=1 filter=113 channel=28
    9, -45, -2, -20, -67, -33, -16, -48, -42,
    -- layer=1 filter=113 channel=29
    -21, -27, -46, -33, -24, -15, -20, -19, -26,
    -- layer=1 filter=113 channel=30
    56, 21, 16, 1, 17, -2, -43, -47, -47,
    -- layer=1 filter=113 channel=31
    2, 5, 30, -1, 6, 0, -37, -55, -12,
    -- layer=1 filter=113 channel=32
    45, -26, 6, -17, -62, -7, -24, -63, -10,
    -- layer=1 filter=113 channel=33
    3, 4, -11, 0, 11, 12, 10, 18, 0,
    -- layer=1 filter=113 channel=34
    3, 22, 4, -15, -17, -6, 12, 4, -19,
    -- layer=1 filter=113 channel=35
    -2, -9, -2, -2, -10, -14, -8, -12, -16,
    -- layer=1 filter=113 channel=36
    9, 3, -1, 11, 1, 13, 39, 29, 30,
    -- layer=1 filter=113 channel=37
    -8, 0, -4, -10, 0, 1, 17, 13, 4,
    -- layer=1 filter=113 channel=38
    37, 32, 41, -7, 7, 14, -28, -15, -31,
    -- layer=1 filter=113 channel=39
    -23, -13, -30, -7, -19, -9, 8, 9, -6,
    -- layer=1 filter=113 channel=40
    -3, 22, 34, -50, -38, -42, -69, -64, -49,
    -- layer=1 filter=113 channel=41
    45, 8, 25, 19, -25, 3, -8, -33, 15,
    -- layer=1 filter=113 channel=42
    -2, -17, 20, 25, 32, 36, -23, -33, -20,
    -- layer=1 filter=113 channel=43
    -4, 9, -17, -8, -8, -16, -2, -1, -7,
    -- layer=1 filter=113 channel=44
    9, -52, 18, -49, -75, -40, -38, -63, 0,
    -- layer=1 filter=113 channel=45
    15, 23, 31, -15, 4, 10, -13, -15, -24,
    -- layer=1 filter=113 channel=46
    60, 54, 53, 0, 4, -3, -86, -74, -58,
    -- layer=1 filter=113 channel=47
    22, 6, 23, -32, -21, -18, -31, -36, -26,
    -- layer=1 filter=113 channel=48
    1, 14, 11, 5, 4, 0, -24, -24, -24,
    -- layer=1 filter=113 channel=49
    17, 39, 32, -1, 22, 14, -37, -20, -41,
    -- layer=1 filter=113 channel=50
    13, -17, -4, 3, -8, -7, -7, -14, -17,
    -- layer=1 filter=113 channel=51
    24, 15, 36, -9, -1, 11, -37, -31, -46,
    -- layer=1 filter=113 channel=52
    -11, 28, 15, 10, 8, -8, 4, 18, -14,
    -- layer=1 filter=113 channel=53
    -2, -9, -14, -7, -13, -17, -11, -16, -3,
    -- layer=1 filter=113 channel=54
    20, -33, 27, -10, -18, 4, 12, -31, 1,
    -- layer=1 filter=113 channel=55
    -10, -9, -6, 11, 13, 9, 37, 49, 42,
    -- layer=1 filter=113 channel=56
    -11, 2, 4, -5, -9, 3, 0, -2, -1,
    -- layer=1 filter=113 channel=57
    25, 7, 31, -17, -25, -5, -48, -80, -49,
    -- layer=1 filter=113 channel=58
    -48, -110, -39, -128, -118, -74, -75, -120, -82,
    -- layer=1 filter=113 channel=59
    2, -5, -12, 6, -2, -13, -9, 7, 3,
    -- layer=1 filter=113 channel=60
    3, -15, -22, -14, -14, -7, -4, -12, -10,
    -- layer=1 filter=113 channel=61
    -8, -11, -9, 0, -7, -2, -7, 7, 0,
    -- layer=1 filter=113 channel=62
    -5, 8, -1, -19, -27, -27, 18, 4, 8,
    -- layer=1 filter=113 channel=63
    6, 0, -13, 18, 5, 8, 29, 12, 28,
    -- layer=1 filter=113 channel=64
    -1, 6, 13, -5, 3, -6, -17, 1, -5,
    -- layer=1 filter=113 channel=65
    -5, 19, 16, -20, -4, -8, -17, -31, -17,
    -- layer=1 filter=113 channel=66
    -4, -15, -14, -6, -8, -2, 4, 8, 7,
    -- layer=1 filter=113 channel=67
    17, 15, 22, 3, 19, 35, -26, -45, -22,
    -- layer=1 filter=113 channel=68
    0, -49, 2, -63, -99, -46, -46, -97, -16,
    -- layer=1 filter=113 channel=69
    -6, 8, 24, -5, -19, 9, 0, 4, -20,
    -- layer=1 filter=113 channel=70
    39, 66, 48, 18, 60, 46, -58, -61, -63,
    -- layer=1 filter=113 channel=71
    4, 0, -11, 5, 6, 12, 11, 3, 3,
    -- layer=1 filter=113 channel=72
    69, 44, 24, 10, 1, -6, -14, -26, -3,
    -- layer=1 filter=113 channel=73
    1, 4, -8, 10, 6, 0, 0, 6, -3,
    -- layer=1 filter=113 channel=74
    15, 26, 6, -18, 20, -6, -38, -69, 45,
    -- layer=1 filter=113 channel=75
    31, 26, 0, 3, -13, -4, -46, -33, 4,
    -- layer=1 filter=113 channel=76
    6, -7, -6, -5, -20, -8, 2, -5, -6,
    -- layer=1 filter=113 channel=77
    10, 11, 3, 11, -5, 0, -9, -10, -18,
    -- layer=1 filter=113 channel=78
    -24, -33, -15, -24, -25, -20, -17, -20, -16,
    -- layer=1 filter=113 channel=79
    5, 19, -1, -5, -12, -15, 7, 0, -3,
    -- layer=1 filter=113 channel=80
    -9, -2, 3, 0, -14, 2, 2, -8, 1,
    -- layer=1 filter=113 channel=81
    -12, -18, -23, -8, -14, -27, 15, 4, 9,
    -- layer=1 filter=113 channel=82
    -1, 8, 13, 5, 13, 7, -23, -18, -27,
    -- layer=1 filter=113 channel=83
    -6, -5, 1, 0, -10, -9, 1, -8, -22,
    -- layer=1 filter=113 channel=84
    29, -3, 12, -26, -28, -31, -48, -61, 24,
    -- layer=1 filter=113 channel=85
    10, -36, -2, -62, -58, -30, -30, -68, -48,
    -- layer=1 filter=113 channel=86
    2, -3, 7, 13, 9, 8, 34, 23, 17,
    -- layer=1 filter=113 channel=87
    78, 56, 64, 18, 22, 5, -31, -37, -46,
    -- layer=1 filter=113 channel=88
    3, 1, -6, -28, -11, -27, -19, -29, -32,
    -- layer=1 filter=113 channel=89
    -3, -6, 23, -9, -4, -15, -19, -28, -22,
    -- layer=1 filter=113 channel=90
    -9, -37, -11, -41, -87, -25, -34, -54, -35,
    -- layer=1 filter=113 channel=91
    23, 51, 51, 5, 21, 21, -23, -13, -14,
    -- layer=1 filter=113 channel=92
    -33, -30, 40, -21, -17, -6, -2, -33, 34,
    -- layer=1 filter=113 channel=93
    0, 15, 8, 0, 3, 3, 0, 15, 3,
    -- layer=1 filter=113 channel=94
    9, -4, 1, 1, 0, -5, 1, -8, -3,
    -- layer=1 filter=113 channel=95
    20, 11, -9, -8, -5, -30, -65, -52, 16,
    -- layer=1 filter=113 channel=96
    1, -11, 0, -11, -3, -10, -1, -7, -9,
    -- layer=1 filter=113 channel=97
    -1, -5, -3, 4, 5, -4, 12, -1, 5,
    -- layer=1 filter=113 channel=98
    23, 50, 31, 11, 4, -23, 16, -10, 10,
    -- layer=1 filter=113 channel=99
    -36, -58, -33, -101, -56, -68, -94, -97, -98,
    -- layer=1 filter=113 channel=100
    3, -9, -22, 8, 8, 4, 24, 16, 13,
    -- layer=1 filter=113 channel=101
    17, 41, 47, 14, 9, 6, -27, -24, -16,
    -- layer=1 filter=113 channel=102
    -5, 0, 13, -20, -18, -5, -21, -28, -33,
    -- layer=1 filter=113 channel=103
    -13, -16, -17, 4, -4, -20, 2, 3, 0,
    -- layer=1 filter=113 channel=104
    40, 2, 28, -7, -29, 3, -12, -19, -40,
    -- layer=1 filter=113 channel=105
    -1, -8, -1, 6, -6, 0, 5, 8, 2,
    -- layer=1 filter=113 channel=106
    48, 43, 48, -3, 4, 23, -30, -28, -2,
    -- layer=1 filter=113 channel=107
    11, -3, 10, 0, 4, 10, 2, 4, 13,
    -- layer=1 filter=113 channel=108
    24, -59, 0, -26, -76, -50, -28, -67, -20,
    -- layer=1 filter=113 channel=109
    2, -3, -2, 7, 10, 5, -6, -4, 0,
    -- layer=1 filter=113 channel=110
    0, -6, -10, 5, 3, 1, -4, -15, -3,
    -- layer=1 filter=113 channel=111
    18, 9, -9, -8, -1, -20, -40, -35, -6,
    -- layer=1 filter=113 channel=112
    -18, -1, 6, 25, 23, 0, -28, -23, 9,
    -- layer=1 filter=113 channel=113
    12, 33, 35, -14, -20, -13, -64, -52, -53,
    -- layer=1 filter=113 channel=114
    -37, -36, -53, -11, -9, -8, 12, 12, -14,
    -- layer=1 filter=113 channel=115
    6, 20, 13, 13, 7, -3, 20, 8, -1,
    -- layer=1 filter=113 channel=116
    -6, 4, -2, 7, 7, -4, 2, -6, -5,
    -- layer=1 filter=113 channel=117
    -6, -3, 1, 7, 14, 5, -104, -64, -20,
    -- layer=1 filter=113 channel=118
    29, 23, 7, -15, -4, -11, -33, -37, 17,
    -- layer=1 filter=113 channel=119
    26, -42, -27, -31, -86, -35, -40, -83, -29,
    -- layer=1 filter=113 channel=120
    13, 37, 26, -5, 3, 7, -12, -24, -34,
    -- layer=1 filter=113 channel=121
    45, 13, 4, -8, 0, -5, 2, 1, -16,
    -- layer=1 filter=113 channel=122
    -7, -3, 4, -2, 7, 8, 3, 6, 1,
    -- layer=1 filter=113 channel=123
    26, -18, -22, 3, -2, 0, 31, 9, 8,
    -- layer=1 filter=113 channel=124
    -7, -4, -14, -6, -10, -9, -10, -1, -1,
    -- layer=1 filter=113 channel=125
    27, 59, 73, -2, 41, 39, -84, -86, -71,
    -- layer=1 filter=113 channel=126
    0, 11, -13, 10, 13, -4, -1, -11, -26,
    -- layer=1 filter=113 channel=127
    33, 16, 15, 8, 13, 2, -22, -41, 28,
    -- layer=1 filter=114 channel=0
    -5, -11, 5, -3, 1, 6, 2, -3, -2,
    -- layer=1 filter=114 channel=1
    19, 27, 0, 22, 14, -17, 13, 3, 0,
    -- layer=1 filter=114 channel=2
    16, 33, 41, 16, 11, 32, -12, 0, -8,
    -- layer=1 filter=114 channel=3
    9, -2, -1, -11, -4, 9, 8, 5, -3,
    -- layer=1 filter=114 channel=4
    4, -8, 2, -5, -1, -11, 2, 5, -4,
    -- layer=1 filter=114 channel=5
    51, 23, 1, 17, 15, -10, 43, 10, 1,
    -- layer=1 filter=114 channel=6
    -20, 2, 17, -42, -34, -62, -43, -24, -48,
    -- layer=1 filter=114 channel=7
    -25, -70, 0, -23, -62, 0, -35, -21, 4,
    -- layer=1 filter=114 channel=8
    35, 31, -4, 47, 38, -4, 27, 31, 9,
    -- layer=1 filter=114 channel=9
    41, -16, -8, -39, 35, -12, -2, 12, 17,
    -- layer=1 filter=114 channel=10
    -19, -51, 11, -29, -48, -3, -1, -14, 19,
    -- layer=1 filter=114 channel=11
    1, -23, -18, 12, -4, -2, -7, -9, 10,
    -- layer=1 filter=114 channel=12
    -28, -27, -9, -8, -4, 4, -8, -2, -10,
    -- layer=1 filter=114 channel=13
    -4, 5, -2, -31, -26, -44, -35, -26, -43,
    -- layer=1 filter=114 channel=14
    -53, -46, -10, 19, -5, 11, -19, 20, 32,
    -- layer=1 filter=114 channel=15
    29, -4, 17, -11, 30, -24, -7, -44, -31,
    -- layer=1 filter=114 channel=16
    37, 13, -10, 24, 8, -17, 17, 19, 8,
    -- layer=1 filter=114 channel=17
    0, -3, -8, -6, -13, -11, -7, -28, -20,
    -- layer=1 filter=114 channel=18
    15, -16, -9, 18, 31, -3, 5, 2, -1,
    -- layer=1 filter=114 channel=19
    65, 21, 36, -28, 1, 14, 10, -56, -40,
    -- layer=1 filter=114 channel=20
    14, 16, -4, -42, -32, -44, -40, -40, -50,
    -- layer=1 filter=114 channel=21
    -53, -17, -25, -23, -14, -9, -36, -2, -4,
    -- layer=1 filter=114 channel=22
    -23, 1, -35, -19, -28, -43, -21, -40, -20,
    -- layer=1 filter=114 channel=23
    -7, -35, -10, -27, -49, -8, -5, -8, -18,
    -- layer=1 filter=114 channel=24
    1, -19, -23, -1, 7, -1, 31, 0, 6,
    -- layer=1 filter=114 channel=25
    8, -13, -9, -32, -61, -6, 0, 4, 2,
    -- layer=1 filter=114 channel=26
    7, -18, -31, -25, 13, -45, 3, -9, -1,
    -- layer=1 filter=114 channel=27
    -39, -36, -43, -7, -35, -26, 3, 7, -6,
    -- layer=1 filter=114 channel=28
    -27, -33, -16, -25, -33, -22, 2, 18, 27,
    -- layer=1 filter=114 channel=29
    -13, 4, -5, -9, 9, -7, -1, 18, -5,
    -- layer=1 filter=114 channel=30
    57, 10, 6, 14, 55, 17, 8, 1, 14,
    -- layer=1 filter=114 channel=31
    0, -5, 5, -12, -6, -25, -24, -24, -21,
    -- layer=1 filter=114 channel=32
    17, -31, -23, -15, -18, -31, 0, 18, 34,
    -- layer=1 filter=114 channel=33
    3, -3, 14, -11, 7, -12, 1, 11, 2,
    -- layer=1 filter=114 channel=34
    -1, -4, 47, 13, 14, 19, 12, -10, -10,
    -- layer=1 filter=114 channel=35
    -11, -2, 0, -3, -10, -4, -4, -16, -8,
    -- layer=1 filter=114 channel=36
    12, 3, 2, 9, 6, 17, 14, 12, 13,
    -- layer=1 filter=114 channel=37
    53, 33, 10, 26, 10, 2, 30, 8, -11,
    -- layer=1 filter=114 channel=38
    23, 12, 15, -21, -15, -12, -36, -33, -38,
    -- layer=1 filter=114 channel=39
    19, -1, 0, 4, 11, 8, -3, -1, 5,
    -- layer=1 filter=114 channel=40
    -1, -5, -22, -21, -16, -55, -19, -41, -38,
    -- layer=1 filter=114 channel=41
    44, -30, -8, 2, 16, -22, 17, 19, 31,
    -- layer=1 filter=114 channel=42
    31, 28, 47, 10, 17, 44, -10, -24, -21,
    -- layer=1 filter=114 channel=43
    12, 8, -13, 8, 20, -2, 27, 13, 22,
    -- layer=1 filter=114 channel=44
    -27, -57, -47, -2, -13, -44, 4, -1, 13,
    -- layer=1 filter=114 channel=45
    -10, 0, 0, -2, 28, -10, -6, -10, -26,
    -- layer=1 filter=114 channel=46
    81, 47, 69, -20, 9, -8, -42, -79, -80,
    -- layer=1 filter=114 channel=47
    -20, -19, 20, -33, -46, -9, -53, 3, -9,
    -- layer=1 filter=114 channel=48
    -7, -14, -1, -13, 0, 3, -28, -25, -8,
    -- layer=1 filter=114 channel=49
    -5, -5, 14, -15, -8, 6, -45, -22, -10,
    -- layer=1 filter=114 channel=50
    9, -29, -2, -25, 0, 0, -10, -27, -14,
    -- layer=1 filter=114 channel=51
    -5, -1, 8, -5, -18, -16, -23, -30, -12,
    -- layer=1 filter=114 channel=52
    26, 14, 17, 26, 6, 6, 16, 14, 13,
    -- layer=1 filter=114 channel=53
    14, 1, 2, 3, -5, 6, 3, 14, 11,
    -- layer=1 filter=114 channel=54
    15, -10, -5, -29, -41, -6, 14, 2, 0,
    -- layer=1 filter=114 channel=55
    -13, -24, -20, 19, 3, 5, 11, -1, 25,
    -- layer=1 filter=114 channel=56
    7, 0, 8, -5, -3, 2, 2, 11, -2,
    -- layer=1 filter=114 channel=57
    -36, -68, -15, -43, -84, -30, -44, -72, -25,
    -- layer=1 filter=114 channel=58
    -18, -92, -16, -37, -113, 1, -34, -28, -28,
    -- layer=1 filter=114 channel=59
    -6, 3, -13, 4, -3, -4, 0, -17, -9,
    -- layer=1 filter=114 channel=60
    -14, -8, -20, -13, -13, -4, 1, -7, -6,
    -- layer=1 filter=114 channel=61
    -7, 5, 2, -6, 0, 4, 2, -1, -6,
    -- layer=1 filter=114 channel=62
    38, 13, -12, 16, 9, -13, 39, 6, 0,
    -- layer=1 filter=114 channel=63
    0, -25, -1, 9, 14, 15, 7, 7, 17,
    -- layer=1 filter=114 channel=64
    -2, 0, 11, 8, -6, 0, 1, 5, -9,
    -- layer=1 filter=114 channel=65
    -23, -12, -22, -9, -9, -14, -12, -10, -22,
    -- layer=1 filter=114 channel=66
    -3, -9, 2, 16, 3, 18, 6, 0, 0,
    -- layer=1 filter=114 channel=67
    -22, -34, -14, -21, -43, -17, -58, -43, -37,
    -- layer=1 filter=114 channel=68
    -26, -60, -36, -3, -17, -48, 7, -18, 4,
    -- layer=1 filter=114 channel=69
    31, 7, -18, 21, 29, -22, 26, -4, -7,
    -- layer=1 filter=114 channel=70
    17, 40, 39, 8, -12, -18, -43, -31, -48,
    -- layer=1 filter=114 channel=71
    -21, -18, -6, 0, 9, 11, 21, 29, 2,
    -- layer=1 filter=114 channel=72
    49, 25, 18, -19, 47, 5, 19, -13, -19,
    -- layer=1 filter=114 channel=73
    -2, 0, 5, -8, -8, -3, -8, -6, -5,
    -- layer=1 filter=114 channel=74
    9, -26, -34, 5, 8, -23, 2, -10, -4,
    -- layer=1 filter=114 channel=75
    20, -11, -14, 16, 26, 10, -4, 33, 1,
    -- layer=1 filter=114 channel=76
    8, -18, -3, 18, 14, 15, 28, 5, 3,
    -- layer=1 filter=114 channel=77
    -30, -19, -10, -12, -7, 5, 3, 9, 1,
    -- layer=1 filter=114 channel=78
    -4, 11, -11, -17, 2, -18, -13, 14, -8,
    -- layer=1 filter=114 channel=79
    33, 13, -14, 17, 14, -5, 15, 8, 2,
    -- layer=1 filter=114 channel=80
    -7, -1, -1, 6, -7, -1, 9, -7, -4,
    -- layer=1 filter=114 channel=81
    -20, -26, -22, -1, 12, 10, 29, 18, 15,
    -- layer=1 filter=114 channel=82
    -20, -11, 6, -23, -2, -2, -27, 0, -16,
    -- layer=1 filter=114 channel=83
    -1, 10, -20, 12, 44, -8, 17, -17, 9,
    -- layer=1 filter=114 channel=84
    19, -15, -12, 16, 36, -10, 11, 2, 8,
    -- layer=1 filter=114 channel=85
    -2, -60, -3, -52, -61, 9, -25, -42, -24,
    -- layer=1 filter=114 channel=86
    12, -5, 9, -7, -15, -9, -3, -2, -16,
    -- layer=1 filter=114 channel=87
    58, 29, 51, -32, 1, 9, -24, -60, -65,
    -- layer=1 filter=114 channel=88
    -10, -13, -10, -14, -1, -12, -20, -17, -16,
    -- layer=1 filter=114 channel=89
    -31, -35, -15, -21, -5, -17, -44, 2, -23,
    -- layer=1 filter=114 channel=90
    -22, -48, -47, -3, -14, -26, 19, 4, 1,
    -- layer=1 filter=114 channel=91
    8, 7, 7, -28, -23, -32, -48, -51, -49,
    -- layer=1 filter=114 channel=92
    3, -46, -23, -24, 10, -45, -8, 17, 5,
    -- layer=1 filter=114 channel=93
    -2, 9, 5, 5, 14, 8, 7, 8, 22,
    -- layer=1 filter=114 channel=94
    4, -3, 4, 0, -4, 2, -23, -12, -9,
    -- layer=1 filter=114 channel=95
    32, 4, 3, 21, 24, 10, 1, 17, 23,
    -- layer=1 filter=114 channel=96
    -6, -8, 7, -6, -6, -3, 0, 0, 18,
    -- layer=1 filter=114 channel=97
    7, 6, -6, 5, 3, 11, 5, 8, 3,
    -- layer=1 filter=114 channel=98
    7, 18, -18, 38, 23, -18, 21, 0, 16,
    -- layer=1 filter=114 channel=99
    -71, -48, -43, -23, 0, -11, 32, 18, 17,
    -- layer=1 filter=114 channel=100
    -17, -29, -21, 17, 3, -15, 8, -7, 2,
    -- layer=1 filter=114 channel=101
    3, 18, 11, -13, -10, -32, -36, -11, -40,
    -- layer=1 filter=114 channel=102
    6, 6, 0, 6, 6, -15, -15, -6, -30,
    -- layer=1 filter=114 channel=103
    -1, -15, -18, 0, -3, 0, -1, -28, 4,
    -- layer=1 filter=114 channel=104
    -5, 8, 4, -17, -24, 5, -16, -2, -12,
    -- layer=1 filter=114 channel=105
    -8, 5, 11, -2, 2, 2, -3, 11, 15,
    -- layer=1 filter=114 channel=106
    8, 14, 2, -44, -31, -36, -47, 6, -34,
    -- layer=1 filter=114 channel=107
    4, 0, -16, 1, 0, 0, 0, 14, 4,
    -- layer=1 filter=114 channel=108
    1, -65, -58, 3, -24, -44, 9, -11, -1,
    -- layer=1 filter=114 channel=109
    -4, -2, -3, -8, 1, -1, 8, -11, -3,
    -- layer=1 filter=114 channel=110
    6, -2, 9, 8, -7, -9, -9, 6, 0,
    -- layer=1 filter=114 channel=111
    29, -14, -8, 30, 43, 4, 6, -14, 4,
    -- layer=1 filter=114 channel=112
    -1, -11, 10, 32, 23, 2, -25, -33, 3,
    -- layer=1 filter=114 channel=113
    7, 26, 53, 5, -2, 25, -36, -71, -33,
    -- layer=1 filter=114 channel=114
    35, 0, -5, 12, 24, -11, 35, 4, -6,
    -- layer=1 filter=114 channel=115
    -9, -7, 12, -11, -7, 0, -9, -20, -4,
    -- layer=1 filter=114 channel=116
    -9, -4, -4, -8, 8, -6, -3, -6, -1,
    -- layer=1 filter=114 channel=117
    35, 12, 18, 28, 1, -9, -21, -28, 10,
    -- layer=1 filter=114 channel=118
    45, -8, 0, 16, 45, -4, 6, 1, 15,
    -- layer=1 filter=114 channel=119
    10, -57, -37, -26, -23, -42, 16, -28, 17,
    -- layer=1 filter=114 channel=120
    -15, -16, -8, -17, -17, -8, -8, -3, 0,
    -- layer=1 filter=114 channel=121
    15, -12, -5, -1, 0, 18, 1, 18, -9,
    -- layer=1 filter=114 channel=122
    0, -9, 9, -6, 2, 1, 0, 4, 2,
    -- layer=1 filter=114 channel=123
    -5, -18, -17, 1, 3, 11, 11, 11, 0,
    -- layer=1 filter=114 channel=124
    1, 11, -3, -12, 0, 4, -1, -1, 0,
    -- layer=1 filter=114 channel=125
    33, 45, 72, 9, 11, 4, -34, -49, -57,
    -- layer=1 filter=114 channel=126
    25, 26, -2, 50, 39, -4, 29, 0, 42,
    -- layer=1 filter=114 channel=127
    43, 4, 12, 30, 53, 11, 20, 0, 25,
    -- layer=1 filter=115 channel=0
    4, 1, 4, 9, 7, -1, 11, 5, 14,
    -- layer=1 filter=115 channel=1
    -1, -4, -2, -4, -17, 7, 2, -25, 18,
    -- layer=1 filter=115 channel=2
    26, 12, 5, 22, 4, -1, -6, -1, -1,
    -- layer=1 filter=115 channel=3
    -15, -9, -4, 6, -3, -7, -14, -3, -4,
    -- layer=1 filter=115 channel=4
    2, -4, -8, 5, -4, -5, -5, 0, 8,
    -- layer=1 filter=115 channel=5
    -4, -10, -12, -6, -16, 10, -7, -30, -4,
    -- layer=1 filter=115 channel=6
    -28, -16, -8, -10, -11, -4, -15, 1, -3,
    -- layer=1 filter=115 channel=7
    -13, 18, 4, -17, 22, -6, 6, 14, -7,
    -- layer=1 filter=115 channel=8
    0, 3, -5, -7, -9, -1, 11, -18, 5,
    -- layer=1 filter=115 channel=9
    7, -13, 6, -20, 7, 16, 9, -4, -2,
    -- layer=1 filter=115 channel=10
    -12, 18, 5, -1, 0, 6, 5, 13, -15,
    -- layer=1 filter=115 channel=11
    -25, -22, -26, -18, -31, -13, -26, -30, -19,
    -- layer=1 filter=115 channel=12
    9, -16, 0, -34, -26, -58, -11, -15, -25,
    -- layer=1 filter=115 channel=13
    -10, -7, -3, -6, -6, 11, 12, 1, 4,
    -- layer=1 filter=115 channel=14
    -14, 9, -1, -20, 2, -13, 20, 0, 5,
    -- layer=1 filter=115 channel=15
    3, -20, -20, -7, -17, 5, 4, -47, -12,
    -- layer=1 filter=115 channel=16
    -1, 6, -6, 5, 1, 2, 0, -16, 8,
    -- layer=1 filter=115 channel=17
    -4, -12, -11, 8, 7, -1, -6, -7, -5,
    -- layer=1 filter=115 channel=18
    -25, -21, -27, 0, -17, -8, -21, -32, -12,
    -- layer=1 filter=115 channel=19
    -5, -19, 0, 16, 8, 44, 29, 41, 26,
    -- layer=1 filter=115 channel=20
    -3, -5, 9, -1, 0, 2, 2, 8, 7,
    -- layer=1 filter=115 channel=21
    -8, -2, 10, 0, 10, -10, -11, 0, 6,
    -- layer=1 filter=115 channel=22
    -9, -8, -9, -10, -3, -12, 3, -4, 3,
    -- layer=1 filter=115 channel=23
    4, -31, 15, -23, -18, 10, 2, -16, 15,
    -- layer=1 filter=115 channel=24
    -5, 8, 1, -13, 8, 14, 0, 15, 5,
    -- layer=1 filter=115 channel=25
    -6, 21, -5, -5, 2, 6, 12, 20, 1,
    -- layer=1 filter=115 channel=26
    7, -8, -19, 2, -1, -3, 19, 9, -1,
    -- layer=1 filter=115 channel=27
    14, 22, 12, 21, 24, 13, -2, -3, 3,
    -- layer=1 filter=115 channel=28
    -11, 25, 16, -11, 21, -4, -1, 4, 10,
    -- layer=1 filter=115 channel=29
    17, 19, 8, 12, 6, 5, -3, -1, -3,
    -- layer=1 filter=115 channel=30
    -22, -14, -6, 10, 9, 16, 25, 11, 21,
    -- layer=1 filter=115 channel=31
    -13, -29, -6, -23, -25, -18, -35, -22, -5,
    -- layer=1 filter=115 channel=32
    -6, -3, 14, -9, 11, 5, 1, -5, -11,
    -- layer=1 filter=115 channel=33
    -2, 0, -10, -17, -8, 0, -3, -6, 0,
    -- layer=1 filter=115 channel=34
    -19, -24, 11, -12, -13, 10, -26, -3, 9,
    -- layer=1 filter=115 channel=35
    20, 11, 1, 2, 16, -1, 11, 7, 4,
    -- layer=1 filter=115 channel=36
    -32, -35, -40, -23, -34, -25, -22, -24, -22,
    -- layer=1 filter=115 channel=37
    3, 6, -2, -6, -6, 14, -2, -9, -15,
    -- layer=1 filter=115 channel=38
    -4, 6, -6, 12, 16, 2, 14, 13, 5,
    -- layer=1 filter=115 channel=39
    0, -9, -7, -11, -2, -3, -4, -8, 5,
    -- layer=1 filter=115 channel=40
    -19, -6, -9, -10, -7, -5, -15, -3, -2,
    -- layer=1 filter=115 channel=41
    4, 14, 19, -13, 5, 7, 22, -7, 2,
    -- layer=1 filter=115 channel=42
    21, 8, -6, 29, 7, -6, -13, -3, -18,
    -- layer=1 filter=115 channel=43
    -1, 25, 0, 0, 4, 21, 7, -15, 12,
    -- layer=1 filter=115 channel=44
    12, 15, 0, -13, 15, -8, 23, 8, -3,
    -- layer=1 filter=115 channel=45
    1, 12, -9, -6, 1, 10, 0, 2, -5,
    -- layer=1 filter=115 channel=46
    -4, -14, -27, -10, -4, -3, 6, 1, 16,
    -- layer=1 filter=115 channel=47
    -8, -14, 17, -23, -3, 21, -15, 1, 5,
    -- layer=1 filter=115 channel=48
    -8, -3, 2, -7, 4, 6, -10, 3, 5,
    -- layer=1 filter=115 channel=49
    1, 1, 21, 3, 4, 17, -5, 4, 0,
    -- layer=1 filter=115 channel=50
    -11, -11, -10, 2, -8, 0, -2, -7, -7,
    -- layer=1 filter=115 channel=51
    -5, 7, 1, 4, 10, 5, -3, 11, 5,
    -- layer=1 filter=115 channel=52
    11, 14, 9, -3, 7, 8, 1, -2, 2,
    -- layer=1 filter=115 channel=53
    10, 2, -1, 15, 14, 7, 8, 14, 3,
    -- layer=1 filter=115 channel=54
    5, 33, 4, 10, -14, 1, 11, 5, -2,
    -- layer=1 filter=115 channel=55
    -23, -19, -12, -21, -20, -20, -25, -23, -16,
    -- layer=1 filter=115 channel=56
    5, 3, 0, -4, 9, -5, 0, 4, -11,
    -- layer=1 filter=115 channel=57
    -23, 3, -6, -12, -4, -6, 0, 14, -17,
    -- layer=1 filter=115 channel=58
    -7, 3, 2, -11, -3, 31, -21, 34, -3,
    -- layer=1 filter=115 channel=59
    0, -2, 13, 1, 12, -5, 6, 11, 1,
    -- layer=1 filter=115 channel=60
    0, 0, -7, -11, -15, 2, -12, 5, -13,
    -- layer=1 filter=115 channel=61
    -5, -14, 3, -16, -11, -1, -3, -1, 1,
    -- layer=1 filter=115 channel=62
    14, 9, -13, 5, -8, 19, 10, -2, 6,
    -- layer=1 filter=115 channel=63
    -22, -2, -16, -1, -5, 3, 0, 0, -2,
    -- layer=1 filter=115 channel=64
    2, 2, 8, -11, -2, 1, 8, 11, 5,
    -- layer=1 filter=115 channel=65
    0, 10, 6, 3, 4, -6, 11, 2, 15,
    -- layer=1 filter=115 channel=66
    2, -6, 4, 1, -6, 13, -1, -2, 4,
    -- layer=1 filter=115 channel=67
    -29, -25, -19, -32, -37, -27, -52, -53, -43,
    -- layer=1 filter=115 channel=68
    0, 12, -2, 0, 11, 0, 9, 11, -11,
    -- layer=1 filter=115 channel=69
    7, -4, -21, -9, -21, -3, -5, -31, -9,
    -- layer=1 filter=115 channel=70
    -37, -32, -2, -28, -39, -13, -44, -38, -18,
    -- layer=1 filter=115 channel=71
    4, 9, 6, 13, 2, 10, -8, 5, -1,
    -- layer=1 filter=115 channel=72
    -3, -31, -14, 2, -8, 22, 15, 0, 20,
    -- layer=1 filter=115 channel=73
    2, -6, 4, 4, -7, -7, 2, 0, 7,
    -- layer=1 filter=115 channel=74
    -7, -16, -9, 0, 19, 0, 11, -4, -8,
    -- layer=1 filter=115 channel=75
    -12, -21, -16, -12, 21, -10, -7, -8, -11,
    -- layer=1 filter=115 channel=76
    5, 12, 0, 2, 14, -8, 11, 2, -8,
    -- layer=1 filter=115 channel=77
    -17, -8, -11, -5, -7, -8, -5, 0, -6,
    -- layer=1 filter=115 channel=78
    1, 9, 7, 12, 2, 8, 1, 11, -1,
    -- layer=1 filter=115 channel=79
    9, 10, -5, 1, -17, 15, 11, -7, 11,
    -- layer=1 filter=115 channel=80
    -7, -5, -8, 0, 7, 6, 6, -6, 0,
    -- layer=1 filter=115 channel=81
    11, 14, 16, -9, 7, 12, -14, 10, 1,
    -- layer=1 filter=115 channel=82
    -8, 3, 9, -1, 6, 10, -6, 9, 8,
    -- layer=1 filter=115 channel=83
    15, -2, -2, -11, 13, 2, 1, -15, -13,
    -- layer=1 filter=115 channel=84
    -6, 0, 8, 20, 6, 13, -2, 4, 0,
    -- layer=1 filter=115 channel=85
    -21, -10, 4, -15, -2, 31, -13, 8, 13,
    -- layer=1 filter=115 channel=86
    -15, -19, -11, -23, -15, -19, -5, -16, -17,
    -- layer=1 filter=115 channel=87
    -25, -15, -17, -12, -16, 26, 16, -8, 1,
    -- layer=1 filter=115 channel=88
    -17, -11, 3, -16, -12, 0, -9, -2, -13,
    -- layer=1 filter=115 channel=89
    0, -4, 14, -10, 17, 13, -6, 4, 3,
    -- layer=1 filter=115 channel=90
    -1, -8, -28, -8, -2, -8, 13, 0, -6,
    -- layer=1 filter=115 channel=91
    4, -6, 5, -5, 8, -1, -1, 16, 7,
    -- layer=1 filter=115 channel=92
    6, 11, 1, -22, 19, -36, 15, 0, -42,
    -- layer=1 filter=115 channel=93
    8, 19, 4, -1, 8, 0, -1, 1, 11,
    -- layer=1 filter=115 channel=94
    -6, -9, 9, 11, 0, 10, 10, -4, 13,
    -- layer=1 filter=115 channel=95
    -18, -3, 0, 17, 18, 21, 14, 0, -2,
    -- layer=1 filter=115 channel=96
    6, -15, 0, 3, 5, 1, 6, 4, -6,
    -- layer=1 filter=115 channel=97
    -3, -7, -7, 8, 13, -7, 13, 10, 5,
    -- layer=1 filter=115 channel=98
    -6, 4, 3, 3, 4, 15, 13, -11, 0,
    -- layer=1 filter=115 channel=99
    -6, 7, -25, 11, -6, -8, 24, 19, 0,
    -- layer=1 filter=115 channel=100
    -12, -28, -26, -35, -8, -12, -11, -12, -11,
    -- layer=1 filter=115 channel=101
    1, -2, -5, 8, 16, -2, 12, 13, 7,
    -- layer=1 filter=115 channel=102
    2, -9, 4, 11, 6, 12, 8, -1, 7,
    -- layer=1 filter=115 channel=103
    -31, -17, -6, -23, -17, -7, -34, -20, -20,
    -- layer=1 filter=115 channel=104
    3, -16, -4, 6, -13, 10, -1, -10, 5,
    -- layer=1 filter=115 channel=105
    -10, 3, 11, 2, 8, 6, -4, -5, 8,
    -- layer=1 filter=115 channel=106
    6, 0, 5, 1, -4, -3, 13, 12, -5,
    -- layer=1 filter=115 channel=107
    -10, -3, 11, 2, 3, -6, -1, -5, 1,
    -- layer=1 filter=115 channel=108
    14, 4, 10, -10, 2, 3, 0, -4, -19,
    -- layer=1 filter=115 channel=109
    -6, 4, 5, 1, 3, 0, 3, -5, 8,
    -- layer=1 filter=115 channel=110
    1, 0, -3, 6, 3, 1, 1, -3, 13,
    -- layer=1 filter=115 channel=111
    -6, -3, -15, 31, -3, 36, 11, 16, 0,
    -- layer=1 filter=115 channel=112
    -20, -10, 2, 2, 2, 1, -4, 0, -12,
    -- layer=1 filter=115 channel=113
    -16, -13, -3, 18, 13, 14, -15, 7, 10,
    -- layer=1 filter=115 channel=114
    -29, -18, -32, -28, -42, -16, -32, -67, -37,
    -- layer=1 filter=115 channel=115
    -5, -14, -11, -10, -2, -1, -14, -7, -23,
    -- layer=1 filter=115 channel=116
    4, 8, 11, -8, 3, -10, 3, -14, 5,
    -- layer=1 filter=115 channel=117
    -5, 4, -2, 15, -11, -8, -12, 14, -9,
    -- layer=1 filter=115 channel=118
    -11, 7, -5, 20, 21, 13, 17, 14, 9,
    -- layer=1 filter=115 channel=119
    -3, 11, -9, 0, 6, -1, 7, 5, -15,
    -- layer=1 filter=115 channel=120
    -10, 1, 8, -2, 8, 9, -1, -6, 14,
    -- layer=1 filter=115 channel=121
    -3, -25, -23, -8, -29, -5, 7, -15, -18,
    -- layer=1 filter=115 channel=122
    -3, -4, 4, 1, -9, 1, -1, 0, 4,
    -- layer=1 filter=115 channel=123
    -6, -33, -20, -28, -8, -12, -11, -1, -23,
    -- layer=1 filter=115 channel=124
    -6, -9, -2, -12, 2, -5, 0, 7, -10,
    -- layer=1 filter=115 channel=125
    -24, -12, -6, -3, -10, 0, -11, -17, -4,
    -- layer=1 filter=115 channel=126
    -1, 3, -1, -9, 4, 22, 26, 1, -4,
    -- layer=1 filter=115 channel=127
    -18, -10, -12, 9, 6, 12, 19, 2, -1,
    -- layer=1 filter=116 channel=0
    -5, -5, -5, 7, -1, 7, -1, -7, -10,
    -- layer=1 filter=116 channel=1
    1, -4, 0, 9, -8, 5, -1, -1, 4,
    -- layer=1 filter=116 channel=2
    -4, -4, 7, -4, -10, 0, 5, 3, -7,
    -- layer=1 filter=116 channel=3
    4, -4, -4, 1, 9, 8, -8, -7, -4,
    -- layer=1 filter=116 channel=4
    -7, -5, -7, 4, 3, 5, 2, 8, 0,
    -- layer=1 filter=116 channel=5
    -5, -7, -2, -11, 6, -3, 0, -10, 0,
    -- layer=1 filter=116 channel=6
    4, -2, 7, -5, 0, 4, 0, -2, 0,
    -- layer=1 filter=116 channel=7
    -9, -5, 14, 0, -2, -6, 5, -6, 5,
    -- layer=1 filter=116 channel=8
    4, 5, -2, -9, -4, 0, -8, -7, 2,
    -- layer=1 filter=116 channel=9
    -5, 7, -1, -11, 1, -7, 8, -6, -4,
    -- layer=1 filter=116 channel=10
    -13, -9, -12, 4, 5, -12, -8, -5, -8,
    -- layer=1 filter=116 channel=11
    0, -8, -6, -2, 10, 2, 1, -4, -7,
    -- layer=1 filter=116 channel=12
    -4, -1, -6, 2, -4, -9, 0, -3, -7,
    -- layer=1 filter=116 channel=13
    5, 5, -8, -9, -12, -8, -12, -11, -6,
    -- layer=1 filter=116 channel=14
    -9, 0, 0, -13, -6, -10, 0, 4, -2,
    -- layer=1 filter=116 channel=15
    -6, 4, 8, 1, 3, -3, -6, -11, -2,
    -- layer=1 filter=116 channel=16
    9, 9, 0, 0, -4, -8, -4, -12, 8,
    -- layer=1 filter=116 channel=17
    5, -5, 5, 0, 7, -6, -6, -3, -2,
    -- layer=1 filter=116 channel=18
    -1, -6, 3, -5, 6, -6, 3, 10, 3,
    -- layer=1 filter=116 channel=19
    -7, 7, 0, 2, 0, 0, -7, -5, 0,
    -- layer=1 filter=116 channel=20
    -6, -4, -7, 3, -11, 7, 6, -6, -10,
    -- layer=1 filter=116 channel=21
    2, -17, 5, 2, -7, -2, 1, -9, 6,
    -- layer=1 filter=116 channel=22
    -3, -5, 4, -5, -7, -6, -9, -9, -9,
    -- layer=1 filter=116 channel=23
    0, 6, -1, -5, -8, 0, -2, 0, -10,
    -- layer=1 filter=116 channel=24
    1, -1, -10, 0, -6, -3, -5, 4, 0,
    -- layer=1 filter=116 channel=25
    6, -1, 5, 0, -6, -6, 3, -5, 6,
    -- layer=1 filter=116 channel=26
    -6, -2, -7, -11, -7, 3, -2, -5, -1,
    -- layer=1 filter=116 channel=27
    0, 6, -6, -1, -8, -8, -5, -7, -14,
    -- layer=1 filter=116 channel=28
    -6, -12, 1, -10, 6, 3, -7, -10, -8,
    -- layer=1 filter=116 channel=29
    7, 5, -1, 0, -6, 3, -8, -7, -7,
    -- layer=1 filter=116 channel=30
    -14, 7, -8, -8, -8, -7, -11, 12, 13,
    -- layer=1 filter=116 channel=31
    5, -9, -3, 3, -5, -1, -7, 6, -10,
    -- layer=1 filter=116 channel=32
    -8, 3, 2, -5, 3, 3, -6, -5, 3,
    -- layer=1 filter=116 channel=33
    5, 5, 3, 2, 10, -7, 0, 7, 1,
    -- layer=1 filter=116 channel=34
    -3, -10, 6, 0, -9, 1, 4, 8, 7,
    -- layer=1 filter=116 channel=35
    1, -6, -11, -12, -7, -3, 6, -11, -4,
    -- layer=1 filter=116 channel=36
    -3, -2, 6, -7, -3, 1, 0, 1, 1,
    -- layer=1 filter=116 channel=37
    1, 0, 4, -1, -7, -12, 0, -12, -8,
    -- layer=1 filter=116 channel=38
    -1, 5, 4, -3, -2, -8, 3, 0, 7,
    -- layer=1 filter=116 channel=39
    -9, -4, 7, 6, 6, -6, -7, -4, 3,
    -- layer=1 filter=116 channel=40
    -1, -9, -11, 6, -1, -2, 5, 1, -9,
    -- layer=1 filter=116 channel=41
    8, 1, 2, 5, 1, -6, 3, -4, 5,
    -- layer=1 filter=116 channel=42
    -6, 0, -7, -7, 3, 6, -1, 1, -12,
    -- layer=1 filter=116 channel=43
    0, 8, -4, 9, -3, -4, -1, -11, 7,
    -- layer=1 filter=116 channel=44
    -12, -11, -11, 2, 8, -2, 2, -5, -1,
    -- layer=1 filter=116 channel=45
    -4, -1, -1, -8, -8, -7, -11, -6, -11,
    -- layer=1 filter=116 channel=46
    -6, -8, 4, -11, -10, -1, 8, -8, 5,
    -- layer=1 filter=116 channel=47
    -11, -7, 1, 5, -7, -14, -8, 0, 1,
    -- layer=1 filter=116 channel=48
    -8, -12, -8, -4, 2, -10, -8, -12, -10,
    -- layer=1 filter=116 channel=49
    -5, 7, -8, -5, -8, -13, -5, -5, 5,
    -- layer=1 filter=116 channel=50
    2, -10, 3, 3, 0, -11, 2, 0, -5,
    -- layer=1 filter=116 channel=51
    -5, 4, -10, -10, 7, -4, 3, -1, -11,
    -- layer=1 filter=116 channel=52
    -1, 3, -3, -5, 8, 3, -8, -8, 5,
    -- layer=1 filter=116 channel=53
    6, 3, -8, -7, -3, -9, 0, 6, 8,
    -- layer=1 filter=116 channel=54
    -8, -2, 3, 4, -1, 0, 6, -4, -5,
    -- layer=1 filter=116 channel=55
    -4, -5, -13, 1, 5, -9, -16, -13, -3,
    -- layer=1 filter=116 channel=56
    0, 6, -3, 3, -4, -10, 7, 5, 3,
    -- layer=1 filter=116 channel=57
    6, 0, 2, -8, -10, -3, -4, -9, -10,
    -- layer=1 filter=116 channel=58
    8, -1, 3, -10, 5, 2, 1, 0, -7,
    -- layer=1 filter=116 channel=59
    -6, -9, 6, 1, -3, -6, -12, 0, -5,
    -- layer=1 filter=116 channel=60
    -6, -5, 4, 5, -4, 2, -2, 8, 5,
    -- layer=1 filter=116 channel=61
    0, 8, 3, -3, 1, -4, -1, 0, -3,
    -- layer=1 filter=116 channel=62
    -2, 0, -5, 7, -6, 3, 1, -7, -10,
    -- layer=1 filter=116 channel=63
    -8, 2, -3, -7, -7, 4, -1, -9, -11,
    -- layer=1 filter=116 channel=64
    -9, 8, 6, -5, 7, -1, 3, -2, 7,
    -- layer=1 filter=116 channel=65
    0, -3, 4, -1, 7, 0, -2, -7, -6,
    -- layer=1 filter=116 channel=66
    -6, -10, -10, -1, -2, 2, -9, 1, 7,
    -- layer=1 filter=116 channel=67
    0, -1, -5, -2, -9, 2, 0, -10, -10,
    -- layer=1 filter=116 channel=68
    -2, -11, -3, -4, -8, -6, 1, -1, -10,
    -- layer=1 filter=116 channel=69
    -7, 11, 7, -3, 1, 8, -5, -8, -13,
    -- layer=1 filter=116 channel=70
    0, 0, 0, 2, -13, -4, -1, 4, 5,
    -- layer=1 filter=116 channel=71
    4, 2, 2, -5, -3, -5, -10, -6, 0,
    -- layer=1 filter=116 channel=72
    -2, 0, 3, -10, 1, 4, -9, -9, 6,
    -- layer=1 filter=116 channel=73
    2, 5, -2, 9, -3, -1, 6, 0, 7,
    -- layer=1 filter=116 channel=74
    -4, 3, 7, -1, -6, 2, 2, 2, -10,
    -- layer=1 filter=116 channel=75
    7, -1, -2, 5, -1, -1, 9, -6, -3,
    -- layer=1 filter=116 channel=76
    -11, -11, 0, 2, -8, 8, -6, -2, 5,
    -- layer=1 filter=116 channel=77
    -2, 5, -1, -10, -5, 0, -7, 7, 4,
    -- layer=1 filter=116 channel=78
    0, -2, -4, -6, 5, -9, -9, 3, -1,
    -- layer=1 filter=116 channel=79
    5, -10, 7, -9, 5, -7, -8, 4, -9,
    -- layer=1 filter=116 channel=80
    7, -4, 12, 3, -5, 5, 4, -1, 10,
    -- layer=1 filter=116 channel=81
    -4, 9, -2, 0, -7, 8, -4, -5, 0,
    -- layer=1 filter=116 channel=82
    4, 4, -1, -1, -5, -9, -2, -8, 2,
    -- layer=1 filter=116 channel=83
    -5, -1, -11, 8, -8, 0, -1, 5, 0,
    -- layer=1 filter=116 channel=84
    -5, 11, 0, 3, 5, 9, -8, 0, -7,
    -- layer=1 filter=116 channel=85
    7, -9, -10, -5, -6, 0, 5, 6, -10,
    -- layer=1 filter=116 channel=86
    4, 1, 2, 4, -1, 0, 7, -9, 2,
    -- layer=1 filter=116 channel=87
    -8, -11, -10, -10, -11, -7, -10, -7, 3,
    -- layer=1 filter=116 channel=88
    1, 5, 2, -12, 6, 8, 4, 1, 1,
    -- layer=1 filter=116 channel=89
    8, 6, -12, -3, -8, -6, 7, -10, -9,
    -- layer=1 filter=116 channel=90
    -5, 3, 2, -11, -11, -10, 6, 3, 4,
    -- layer=1 filter=116 channel=91
    -11, 3, -11, -2, -8, 5, -12, 0, -5,
    -- layer=1 filter=116 channel=92
    -5, 6, -2, 2, -3, 4, 9, -8, -4,
    -- layer=1 filter=116 channel=93
    5, 4, -6, -5, 3, 0, -7, -11, -8,
    -- layer=1 filter=116 channel=94
    2, 3, -8, -4, 2, 7, 5, -2, -3,
    -- layer=1 filter=116 channel=95
    7, -6, -2, -7, -4, 4, 10, 10, -10,
    -- layer=1 filter=116 channel=96
    -5, 9, -1, -1, 6, 8, -11, 5, -12,
    -- layer=1 filter=116 channel=97
    2, -7, -9, 0, -7, 1, -6, 4, -2,
    -- layer=1 filter=116 channel=98
    8, -2, -4, -4, -8, -9, -3, 0, 0,
    -- layer=1 filter=116 channel=99
    -7, -10, 0, -11, -6, -5, 4, 7, -10,
    -- layer=1 filter=116 channel=100
    1, 5, 0, 6, -5, 3, 6, -11, -5,
    -- layer=1 filter=116 channel=101
    -11, -4, 4, -3, 6, 6, 0, 3, -11,
    -- layer=1 filter=116 channel=102
    -2, 3, 4, 0, -6, -9, -7, 1, -7,
    -- layer=1 filter=116 channel=103
    -1, 4, 8, -6, -2, 2, 5, 0, 2,
    -- layer=1 filter=116 channel=104
    -5, -3, -4, 3, -10, 2, 0, -6, -11,
    -- layer=1 filter=116 channel=105
    -10, -5, -1, 8, -6, -9, 5, -10, 2,
    -- layer=1 filter=116 channel=106
    -5, 6, -8, -7, -7, -9, -6, -10, -6,
    -- layer=1 filter=116 channel=107
    8, 5, 0, -7, -10, 2, 3, -8, 5,
    -- layer=1 filter=116 channel=108
    1, 4, -7, -3, -10, -12, -10, -20, -9,
    -- layer=1 filter=116 channel=109
    3, 3, 4, 0, -2, 0, 6, 9, -3,
    -- layer=1 filter=116 channel=110
    -8, -7, 7, -7, 6, 7, -2, 0, 6,
    -- layer=1 filter=116 channel=111
    -4, 2, -2, -7, 0, 2, 2, 10, -5,
    -- layer=1 filter=116 channel=112
    6, 0, 4, 4, 0, 6, -11, -1, -10,
    -- layer=1 filter=116 channel=113
    -1, -11, 3, 7, 7, -5, 8, 0, -6,
    -- layer=1 filter=116 channel=114
    12, 9, -1, -10, 6, 0, 3, -10, 1,
    -- layer=1 filter=116 channel=115
    -9, -7, -6, 0, 6, 5, -11, -8, -5,
    -- layer=1 filter=116 channel=116
    4, -1, -6, -10, -10, 10, -9, 0, 9,
    -- layer=1 filter=116 channel=117
    -4, -1, -8, -4, 8, -7, -4, 2, 1,
    -- layer=1 filter=116 channel=118
    -8, 0, -11, 3, -3, 5, 10, 4, 5,
    -- layer=1 filter=116 channel=119
    -1, 6, 0, -11, -15, 8, -15, 6, 6,
    -- layer=1 filter=116 channel=120
    3, -10, -14, -11, -9, 3, -13, -1, -13,
    -- layer=1 filter=116 channel=121
    3, 4, 8, -1, -15, -8, 6, 5, 5,
    -- layer=1 filter=116 channel=122
    9, 0, 5, 2, -1, -6, 0, -3, 10,
    -- layer=1 filter=116 channel=123
    5, -4, 2, -13, 6, -9, 0, 5, -8,
    -- layer=1 filter=116 channel=124
    9, -1, 4, -3, -9, 1, -1, -1, -3,
    -- layer=1 filter=116 channel=125
    4, -14, -15, -12, -10, 1, 3, -4, -8,
    -- layer=1 filter=116 channel=126
    -8, 8, 8, -3, -11, -1, -10, -3, -5,
    -- layer=1 filter=116 channel=127
    -11, -8, -8, -8, -7, 8, 1, 4, -12,
    -- layer=1 filter=117 channel=0
    -5, 0, 10, -19, 18, 14, -17, 3, 4,
    -- layer=1 filter=117 channel=1
    -35, -44, -51, 1, -63, -53, -25, 29, 11,
    -- layer=1 filter=117 channel=2
    -36, -48, -58, -6, -10, -27, 14, -14, 6,
    -- layer=1 filter=117 channel=3
    -9, -9, -10, -1, -6, 1, 2, -11, 3,
    -- layer=1 filter=117 channel=4
    1, -3, -6, -5, 5, 10, 5, -6, 6,
    -- layer=1 filter=117 channel=5
    -72, -80, -97, -33, -125, -89, 1, 37, 36,
    -- layer=1 filter=117 channel=6
    29, 11, 21, 32, -22, 9, 31, 0, -27,
    -- layer=1 filter=117 channel=7
    33, 49, -100, 40, 51, -100, 22, 93, -40,
    -- layer=1 filter=117 channel=8
    -68, -117, -135, -43, -130, -92, -1, 42, 26,
    -- layer=1 filter=117 channel=9
    -95, -49, -50, 35, -13, -6, 3, 16, 26,
    -- layer=1 filter=117 channel=10
    38, 59, -83, 18, 58, -47, 50, 96, -9,
    -- layer=1 filter=117 channel=11
    5, -9, -6, 6, 0, 5, -5, -4, 9,
    -- layer=1 filter=117 channel=12
    -48, -19, -28, 16, 12, 21, -6, 16, 31,
    -- layer=1 filter=117 channel=13
    -20, -9, 18, -7, -9, 20, -11, -19, 18,
    -- layer=1 filter=117 channel=14
    27, 28, -80, 70, 88, -45, -14, 115, -71,
    -- layer=1 filter=117 channel=15
    -35, -78, 21, -39, -43, -9, 1, -10, -25,
    -- layer=1 filter=117 channel=16
    -100, -111, -141, -46, -112, -107, 15, 53, 23,
    -- layer=1 filter=117 channel=17
    -19, -2, 1, -15, -7, 22, -22, -7, 17,
    -- layer=1 filter=117 channel=18
    -5, -52, -64, 20, 28, 19, 20, 27, 17,
    -- layer=1 filter=117 channel=19
    -80, -104, -92, -33, -63, -74, 30, -32, -51,
    -- layer=1 filter=117 channel=20
    -13, -9, 32, -31, -21, 12, -17, -26, 3,
    -- layer=1 filter=117 channel=21
    -9, -38, -44, 19, -24, -37, -7, 13, -13,
    -- layer=1 filter=117 channel=22
    -32, -15, -7, -12, -30, 0, -16, -2, 1,
    -- layer=1 filter=117 channel=23
    54, -1, 1, 70, -17, -19, 25, 5, -55,
    -- layer=1 filter=117 channel=24
    -33, -30, -21, -16, -21, -17, 6, 19, 26,
    -- layer=1 filter=117 channel=25
    25, 0, -93, -13, 9, -99, 32, 58, -11,
    -- layer=1 filter=117 channel=26
    -58, -51, 24, -41, -55, 5, -30, -75, 26,
    -- layer=1 filter=117 channel=27
    -10, 0, -22, 3, 4, -6, 7, 12, 8,
    -- layer=1 filter=117 channel=28
    4, 42, -76, 13, 47, -59, 13, 82, -14,
    -- layer=1 filter=117 channel=29
    -8, 6, -11, -6, 4, -1, -37, -21, -12,
    -- layer=1 filter=117 channel=30
    -19, -73, -135, 12, 31, -3, 23, 1, -10,
    -- layer=1 filter=117 channel=31
    -33, -43, -49, 1, 8, -6, 18, 33, -34,
    -- layer=1 filter=117 channel=32
    -29, -90, -3, -10, -97, -1, -14, -81, 23,
    -- layer=1 filter=117 channel=33
    7, -2, -7, 2, -11, -15, -12, -1, -7,
    -- layer=1 filter=117 channel=34
    18, 9, 9, 12, -11, 2, 18, 12, 19,
    -- layer=1 filter=117 channel=35
    -2, -16, -2, -7, 1, -16, -2, -7, -7,
    -- layer=1 filter=117 channel=36
    12, 9, 12, 19, 31, 9, 6, 0, 19,
    -- layer=1 filter=117 channel=37
    -72, -140, -134, -97, -125, -126, 20, 30, 30,
    -- layer=1 filter=117 channel=38
    -8, -12, 28, -12, -25, -2, 0, -12, -6,
    -- layer=1 filter=117 channel=39
    -11, -9, -26, -19, -5, -5, -19, -12, -7,
    -- layer=1 filter=117 channel=40
    -46, -17, -57, -4, 0, -30, 37, 22, -45,
    -- layer=1 filter=117 channel=41
    -6, -8, -10, 24, -24, -21, 4, -36, -2,
    -- layer=1 filter=117 channel=42
    -19, -31, -59, 25, 7, -39, 41, -18, 1,
    -- layer=1 filter=117 channel=43
    -46, -34, -110, -32, -81, -92, 15, 48, 22,
    -- layer=1 filter=117 channel=44
    -57, -47, 5, -45, -91, 10, -20, -66, 47,
    -- layer=1 filter=117 channel=45
    -26, -25, 8, -10, -24, -7, -12, -15, 24,
    -- layer=1 filter=117 channel=46
    -23, -87, -17, 7, -36, -66, 69, -10, -14,
    -- layer=1 filter=117 channel=47
    38, -56, -6, 41, -64, -45, 37, 26, -44,
    -- layer=1 filter=117 channel=48
    15, -11, 6, 0, -5, 1, -4, 7, -16,
    -- layer=1 filter=117 channel=49
    -24, -6, -7, 15, -4, -5, 14, 6, -2,
    -- layer=1 filter=117 channel=50
    -11, 1, -5, 1, -10, 11, 9, -2, -3,
    -- layer=1 filter=117 channel=51
    12, 20, -10, -4, 29, -14, 12, 33, -20,
    -- layer=1 filter=117 channel=52
    -2, 6, 7, 15, 18, -1, -24, -13, -1,
    -- layer=1 filter=117 channel=53
    -10, -12, -1, -8, -14, -4, -5, -13, 10,
    -- layer=1 filter=117 channel=54
    12, -12, -84, -40, 2, -77, 54, 50, 17,
    -- layer=1 filter=117 channel=55
    28, -6, -1, 21, 11, -4, 21, 2, -4,
    -- layer=1 filter=117 channel=56
    7, 0, -7, 0, -3, 8, 6, 4, 0,
    -- layer=1 filter=117 channel=57
    17, 35, -98, -8, 32, -70, 49, 56, -27,
    -- layer=1 filter=117 channel=58
    69, -7, -69, 55, 6, -69, 69, 78, -80,
    -- layer=1 filter=117 channel=59
    -4, 0, -4, -4, -2, -8, -7, -11, -3,
    -- layer=1 filter=117 channel=60
    4, -4, 6, 13, 12, 0, 7, -4, 4,
    -- layer=1 filter=117 channel=61
    -5, 7, 0, 6, 0, 9, -5, 0, -2,
    -- layer=1 filter=117 channel=62
    -115, -154, -112, -102, -140, -128, 10, 21, 17,
    -- layer=1 filter=117 channel=63
    9, 5, 4, 35, 22, 13, 2, 6, 11,
    -- layer=1 filter=117 channel=64
    -3, -5, 6, -8, -14, -10, -8, -2, -12,
    -- layer=1 filter=117 channel=65
    -27, 2, -2, -25, -2, -2, -21, -11, -11,
    -- layer=1 filter=117 channel=66
    18, 24, 1, 8, 10, 4, -8, 5, 6,
    -- layer=1 filter=117 channel=67
    -15, -3, -1, 12, 0, -4, -8, -11, -23,
    -- layer=1 filter=117 channel=68
    -80, -42, -14, -60, -71, 8, -32, -60, 67,
    -- layer=1 filter=117 channel=69
    -55, -92, -36, -39, -93, -53, -1, 26, 18,
    -- layer=1 filter=117 channel=70
    20, -6, 7, 32, -12, 1, 28, 3, -47,
    -- layer=1 filter=117 channel=71
    7, 16, -10, 18, -9, -16, 16, 14, -6,
    -- layer=1 filter=117 channel=72
    -49, -62, -51, 16, -2, 3, 21, -2, -7,
    -- layer=1 filter=117 channel=73
    -7, 7, -6, 5, 9, 2, -1, -4, -5,
    -- layer=1 filter=117 channel=74
    -54, -1, -11, -30, -16, 21, -5, -10, 63,
    -- layer=1 filter=117 channel=75
    12, -49, -52, 76, 70, 42, 32, 55, -10,
    -- layer=1 filter=117 channel=76
    -8, -19, 1, -20, -6, 13, -7, -24, 17,
    -- layer=1 filter=117 channel=77
    9, -13, -15, -7, -18, -15, 0, 13, 0,
    -- layer=1 filter=117 channel=78
    24, 20, 7, 10, 25, -15, 4, 31, 2,
    -- layer=1 filter=117 channel=79
    -61, -129, -94, -66, -119, -108, 15, 13, 1,
    -- layer=1 filter=117 channel=80
    -9, -12, -11, -4, -4, 0, -1, -10, 5,
    -- layer=1 filter=117 channel=81
    13, -3, -34, -1, 0, -24, 48, 21, 6,
    -- layer=1 filter=117 channel=82
    -19, -30, -15, 1, -25, -20, -1, -28, -14,
    -- layer=1 filter=117 channel=83
    -8, -24, -9, -21, -16, 9, 3, 11, 32,
    -- layer=1 filter=117 channel=84
    -73, -91, -63, -8, 3, 21, 19, -21, 42,
    -- layer=1 filter=117 channel=85
    61, -8, -3, 39, -27, -22, 57, 4, -40,
    -- layer=1 filter=117 channel=86
    6, 11, 15, -3, 8, 10, -12, 18, -4,
    -- layer=1 filter=117 channel=87
    -59, -31, -37, 19, -47, -6, 50, -7, -39,
    -- layer=1 filter=117 channel=88
    -2, 12, 5, 12, 15, 5, 17, 20, 4,
    -- layer=1 filter=117 channel=89
    -32, -23, -4, -12, -28, -8, -22, -37, -5,
    -- layer=1 filter=117 channel=90
    -61, -67, -10, -49, -66, 8, -20, -47, 35,
    -- layer=1 filter=117 channel=91
    -6, -1, 7, -5, -7, -9, -2, -7, -5,
    -- layer=1 filter=117 channel=92
    -29, -40, 4, -36, -52, -18, -42, -23, 1,
    -- layer=1 filter=117 channel=93
    8, 3, 5, -13, 3, -3, -8, 0, 7,
    -- layer=1 filter=117 channel=94
    -6, 19, 20, -4, 25, 6, -6, 17, -1,
    -- layer=1 filter=117 channel=95
    -59, -122, -83, -1, -11, 16, -2, 3, 11,
    -- layer=1 filter=117 channel=96
    4, -4, 13, 13, 14, 1, 3, 19, 23,
    -- layer=1 filter=117 channel=97
    0, 10, 11, -14, -6, 8, -8, 10, 19,
    -- layer=1 filter=117 channel=98
    -63, -40, -87, -51, -60, -66, 18, 37, -4,
    -- layer=1 filter=117 channel=99
    -26, 72, -12, -39, 81, 12, 7, 45, 21,
    -- layer=1 filter=117 channel=100
    0, -19, -10, 17, 10, -3, -8, -7, -6,
    -- layer=1 filter=117 channel=101
    -15, -1, 9, -24, -11, 6, -19, -16, 9,
    -- layer=1 filter=117 channel=102
    -2, 4, 13, -17, 21, 24, -24, 3, 14,
    -- layer=1 filter=117 channel=103
    9, 6, 6, 5, 8, 2, -2, 0, -4,
    -- layer=1 filter=117 channel=104
    28, -16, -19, 23, -3, -7, -2, 13, -38,
    -- layer=1 filter=117 channel=105
    11, 28, 13, -4, 19, 1, 5, 22, 2,
    -- layer=1 filter=117 channel=106
    -43, -33, 11, -43, -50, 17, -33, -53, 9,
    -- layer=1 filter=117 channel=107
    10, 13, 14, -3, 5, 6, 9, 2, 15,
    -- layer=1 filter=117 channel=108
    -60, -129, 0, -57, -139, -3, -44, -95, 14,
    -- layer=1 filter=117 channel=109
    1, 2, -7, 5, -3, 0, -7, -1, -10,
    -- layer=1 filter=117 channel=110
    6, 10, 6, 9, 25, -1, 2, 11, 11,
    -- layer=1 filter=117 channel=111
    -15, -64, -79, 15, 41, 19, 39, 38, 16,
    -- layer=1 filter=117 channel=112
    -19, -38, -31, 29, 23, 20, 38, 32, 19,
    -- layer=1 filter=117 channel=113
    -11, -36, -26, 19, -16, -40, 7, -34, -7,
    -- layer=1 filter=117 channel=114
    -53, -71, -88, -7, -52, -71, 39, 25, 30,
    -- layer=1 filter=117 channel=115
    5, 30, -4, 1, 26, -9, 8, 40, 12,
    -- layer=1 filter=117 channel=116
    0, 3, 0, 4, 9, 4, -5, 8, 8,
    -- layer=1 filter=117 channel=117
    -20, -54, -34, 37, 31, 2, 51, 81, 7,
    -- layer=1 filter=117 channel=118
    -42, -68, -37, -11, 9, 36, 31, -5, 47,
    -- layer=1 filter=117 channel=119
    -46, -76, -23, -53, -120, -5, -20, -98, 18,
    -- layer=1 filter=117 channel=120
    15, -5, -33, -2, -8, -36, 13, 31, -20,
    -- layer=1 filter=117 channel=121
    -4, -46, -39, 44, 32, 5, 1, 1, -63,
    -- layer=1 filter=117 channel=122
    7, 8, -8, 3, 2, 0, -6, 1, -3,
    -- layer=1 filter=117 channel=123
    36, 5, -16, 65, 38, 9, 27, 24, -18,
    -- layer=1 filter=117 channel=124
    -7, -15, 1, -13, 2, 0, 0, 9, -2,
    -- layer=1 filter=117 channel=125
    21, 28, 23, 19, -1, 3, 32, -4, -30,
    -- layer=1 filter=117 channel=126
    -67, -76, -64, -35, -95, -77, 0, 12, -19,
    -- layer=1 filter=117 channel=127
    -37, -100, -82, 7, 10, 18, 21, 10, 26,
    -- layer=1 filter=118 channel=0
    1, 3, -11, -4, -6, 6, -3, 7, 7,
    -- layer=1 filter=118 channel=1
    -1, 1, 1, 1, -11, 2, 7, -1, -8,
    -- layer=1 filter=118 channel=2
    -7, 3, -6, 6, -7, 4, 2, -1, 11,
    -- layer=1 filter=118 channel=3
    -11, -1, -8, 0, -7, 3, -5, -1, 0,
    -- layer=1 filter=118 channel=4
    -9, 8, 5, 1, -10, -3, 1, -1, 7,
    -- layer=1 filter=118 channel=5
    6, -6, -13, 3, -7, -10, -4, 4, -3,
    -- layer=1 filter=118 channel=6
    -4, 4, 0, -5, -7, -3, -1, -4, -9,
    -- layer=1 filter=118 channel=7
    -7, -15, 5, -2, 1, 3, 3, -1, 0,
    -- layer=1 filter=118 channel=8
    0, -8, 6, 4, 7, -2, 2, 6, -2,
    -- layer=1 filter=118 channel=9
    -5, 3, -5, -9, 4, 4, -4, 4, 0,
    -- layer=1 filter=118 channel=10
    3, -5, 0, -13, 3, 0, -2, -3, -5,
    -- layer=1 filter=118 channel=11
    -3, -9, -3, 9, 0, 0, -10, 4, 3,
    -- layer=1 filter=118 channel=12
    2, -4, 8, -6, 6, 1, -3, -8, 5,
    -- layer=1 filter=118 channel=13
    1, 6, 4, -6, -1, -5, 4, 3, 3,
    -- layer=1 filter=118 channel=14
    -7, -9, 4, -3, -7, -9, -10, -7, -8,
    -- layer=1 filter=118 channel=15
    1, -5, 0, -4, -10, -2, 0, 2, -6,
    -- layer=1 filter=118 channel=16
    3, -5, 6, -6, 1, 0, 0, -3, 7,
    -- layer=1 filter=118 channel=17
    -10, -5, -3, -6, -8, -11, -11, 5, -10,
    -- layer=1 filter=118 channel=18
    -2, -11, -12, 3, -2, -4, 8, -11, 8,
    -- layer=1 filter=118 channel=19
    8, -10, 7, 1, -4, -11, 4, -7, 0,
    -- layer=1 filter=118 channel=20
    0, -9, -10, 0, 2, 6, -12, -5, -3,
    -- layer=1 filter=118 channel=21
    -10, 9, 0, 6, 1, 1, -3, 5, -5,
    -- layer=1 filter=118 channel=22
    -11, 3, 3, 7, -4, 3, 0, 0, -11,
    -- layer=1 filter=118 channel=23
    -11, -11, -8, -6, -2, -12, -11, -7, -3,
    -- layer=1 filter=118 channel=24
    1, -8, -5, -1, 2, -5, -10, -9, 0,
    -- layer=1 filter=118 channel=25
    7, -4, 3, 0, -4, -7, 0, 1, -5,
    -- layer=1 filter=118 channel=26
    -5, 4, -8, 6, -2, -10, -6, -12, 0,
    -- layer=1 filter=118 channel=27
    7, 5, 0, -3, 4, -2, -4, -5, 0,
    -- layer=1 filter=118 channel=28
    1, -2, -6, 1, -4, -11, -6, 8, 1,
    -- layer=1 filter=118 channel=29
    -8, 3, -4, -3, -11, -10, 0, -1, -2,
    -- layer=1 filter=118 channel=30
    -3, 1, -10, -4, -7, -4, 1, -7, 1,
    -- layer=1 filter=118 channel=31
    5, -7, -5, 0, -8, -9, 2, -7, -7,
    -- layer=1 filter=118 channel=32
    -9, -2, 1, -9, -4, 8, -4, -4, -3,
    -- layer=1 filter=118 channel=33
    9, -7, -5, 3, 0, 6, 4, 6, 3,
    -- layer=1 filter=118 channel=34
    4, -8, 2, -6, 6, -5, 1, -6, -4,
    -- layer=1 filter=118 channel=35
    -13, 1, -2, 4, 2, -10, -12, -12, -6,
    -- layer=1 filter=118 channel=36
    -5, -9, 4, -7, -3, -6, -4, 7, -9,
    -- layer=1 filter=118 channel=37
    9, -9, 6, 1, -4, 1, 0, -7, 0,
    -- layer=1 filter=118 channel=38
    3, 0, 4, 5, 0, -6, 0, 9, -6,
    -- layer=1 filter=118 channel=39
    -1, 4, 3, -2, -11, -1, -3, -4, 5,
    -- layer=1 filter=118 channel=40
    2, 1, -1, 8, -3, -6, -3, -9, 7,
    -- layer=1 filter=118 channel=41
    -5, -4, -11, 1, -6, -11, -7, -3, -8,
    -- layer=1 filter=118 channel=42
    -3, 9, 7, 4, 2, 0, -9, 1, -5,
    -- layer=1 filter=118 channel=43
    -10, 4, -12, 1, 1, -5, 5, -2, -7,
    -- layer=1 filter=118 channel=44
    -2, 4, 3, -7, -12, -6, 2, 5, 7,
    -- layer=1 filter=118 channel=45
    6, -7, -8, -9, -10, 9, -10, 1, -8,
    -- layer=1 filter=118 channel=46
    2, 1, -4, 7, 2, -4, -11, -3, -5,
    -- layer=1 filter=118 channel=47
    0, -4, -12, -3, -13, -11, -4, 2, 0,
    -- layer=1 filter=118 channel=48
    -3, -1, 2, 0, -7, -8, -12, 0, 3,
    -- layer=1 filter=118 channel=49
    -4, 0, 2, 7, 4, -4, 6, -6, -9,
    -- layer=1 filter=118 channel=50
    6, -1, -6, 0, 2, -2, 0, -8, 6,
    -- layer=1 filter=118 channel=51
    0, -12, -8, -13, 5, -7, 0, 4, -4,
    -- layer=1 filter=118 channel=52
    5, 8, -11, -12, -2, -3, 3, 6, -5,
    -- layer=1 filter=118 channel=53
    7, 3, -8, -9, 7, 3, 1, 1, -2,
    -- layer=1 filter=118 channel=54
    -2, 0, -3, 3, -3, -10, -7, -13, -6,
    -- layer=1 filter=118 channel=55
    -9, 4, 0, -3, 0, 4, -1, 7, 0,
    -- layer=1 filter=118 channel=56
    1, 7, -9, -12, 3, 6, 1, -10, -3,
    -- layer=1 filter=118 channel=57
    3, 8, -3, -5, 0, -4, -8, -4, 5,
    -- layer=1 filter=118 channel=58
    4, 8, -8, 7, -9, 4, -2, 4, 2,
    -- layer=1 filter=118 channel=59
    -7, -2, 2, 9, 6, -6, -11, -8, -2,
    -- layer=1 filter=118 channel=60
    0, 5, -9, 9, -3, -10, -1, 2, -5,
    -- layer=1 filter=118 channel=61
    0, 6, -1, -3, 1, 8, -5, 0, -11,
    -- layer=1 filter=118 channel=62
    -8, 0, 7, -5, -8, -10, 5, 5, -8,
    -- layer=1 filter=118 channel=63
    -1, -8, 6, -7, 4, -1, -2, 2, 0,
    -- layer=1 filter=118 channel=64
    -5, 3, 6, -11, -3, 6, -12, -11, -8,
    -- layer=1 filter=118 channel=65
    2, 0, -4, 2, -6, -6, -1, -2, -9,
    -- layer=1 filter=118 channel=66
    -4, -6, 0, -1, -10, 1, 4, 1, -7,
    -- layer=1 filter=118 channel=67
    5, -5, 6, -5, 0, -11, 9, 9, -9,
    -- layer=1 filter=118 channel=68
    -7, -1, -5, 6, -8, 7, 0, -12, -7,
    -- layer=1 filter=118 channel=69
    -4, -8, 0, -10, 0, -8, -1, 1, 5,
    -- layer=1 filter=118 channel=70
    3, -4, 3, -2, 8, -7, -7, 9, -6,
    -- layer=1 filter=118 channel=71
    -10, -2, 1, 0, -10, 5, 0, 5, -8,
    -- layer=1 filter=118 channel=72
    -2, -2, 5, 3, 1, 1, -9, -2, 4,
    -- layer=1 filter=118 channel=73
    -7, -8, -3, 7, -1, 5, -2, 2, -4,
    -- layer=1 filter=118 channel=74
    0, -1, 0, 4, -8, -3, 7, -8, -9,
    -- layer=1 filter=118 channel=75
    -3, -8, -2, 7, 2, 11, -9, 6, 5,
    -- layer=1 filter=118 channel=76
    3, -6, 8, 8, -2, 7, 5, 7, -11,
    -- layer=1 filter=118 channel=77
    3, -2, 5, -4, 4, 0, 6, 7, 1,
    -- layer=1 filter=118 channel=78
    0, 2, 4, -7, -11, 4, 0, 8, -7,
    -- layer=1 filter=118 channel=79
    -7, -1, -8, 2, -7, 0, -3, 0, -3,
    -- layer=1 filter=118 channel=80
    0, -5, -13, -6, -10, -1, -3, 6, -1,
    -- layer=1 filter=118 channel=81
    -9, 4, 8, 4, -3, 3, -4, -11, -9,
    -- layer=1 filter=118 channel=82
    0, 0, 1, -12, 8, -10, -9, 1, 5,
    -- layer=1 filter=118 channel=83
    6, 5, -6, -11, 3, -8, 4, -5, -6,
    -- layer=1 filter=118 channel=84
    -12, 5, 2, -5, 1, 6, -9, 6, 7,
    -- layer=1 filter=118 channel=85
    9, 7, 1, -5, -8, -8, 1, 3, -8,
    -- layer=1 filter=118 channel=86
    7, -2, -7, -6, -10, -1, -11, -11, 0,
    -- layer=1 filter=118 channel=87
    -1, 4, -11, -10, 1, 4, -5, -9, 5,
    -- layer=1 filter=118 channel=88
    -9, 0, -8, -8, -1, 0, -11, 3, -4,
    -- layer=1 filter=118 channel=89
    0, -1, 3, -12, 6, 0, -9, 8, -9,
    -- layer=1 filter=118 channel=90
    0, -7, -3, 3, 7, -2, 5, 4, 4,
    -- layer=1 filter=118 channel=91
    -4, -4, 7, -7, 8, 6, -2, -2, 6,
    -- layer=1 filter=118 channel=92
    -5, -6, 0, -8, 7, -4, 8, 3, -6,
    -- layer=1 filter=118 channel=93
    3, -2, -7, 7, 5, 2, -5, -2, -7,
    -- layer=1 filter=118 channel=94
    4, 5, -1, -7, 7, -2, 2, 8, 3,
    -- layer=1 filter=118 channel=95
    -6, 6, -13, 5, -12, 5, -2, 8, -10,
    -- layer=1 filter=118 channel=96
    -10, -1, -8, -12, 4, 5, 1, -5, -7,
    -- layer=1 filter=118 channel=97
    4, 4, 7, 4, -1, -10, -2, -3, -4,
    -- layer=1 filter=118 channel=98
    -10, -4, 3, -12, -6, -7, -4, -12, 6,
    -- layer=1 filter=118 channel=99
    6, 4, -5, 5, -10, -9, -9, 1, -10,
    -- layer=1 filter=118 channel=100
    0, 3, 0, 8, 5, -8, 7, 0, -2,
    -- layer=1 filter=118 channel=101
    4, -6, 8, -2, 6, -10, -7, 5, 6,
    -- layer=1 filter=118 channel=102
    -10, 7, 4, -10, -5, -6, 3, 7, 6,
    -- layer=1 filter=118 channel=103
    7, -6, -2, 0, -8, 4, -3, 7, 1,
    -- layer=1 filter=118 channel=104
    -5, 1, 1, -12, -10, 7, -10, -7, -7,
    -- layer=1 filter=118 channel=105
    0, 3, 7, 5, -1, 8, -9, 0, 5,
    -- layer=1 filter=118 channel=106
    -6, -1, 5, 7, -2, 1, 2, -8, -6,
    -- layer=1 filter=118 channel=107
    4, -5, -3, 3, -6, -4, -11, -9, 1,
    -- layer=1 filter=118 channel=108
    -6, -10, -8, -3, -1, 2, 2, -6, -2,
    -- layer=1 filter=118 channel=109
    9, 10, 1, -9, 7, 8, 10, -1, 8,
    -- layer=1 filter=118 channel=110
    -4, 2, -4, -6, 3, 2, -4, -11, 0,
    -- layer=1 filter=118 channel=111
    7, -3, -2, -14, -11, -7, 5, 6, -5,
    -- layer=1 filter=118 channel=112
    -6, -7, -5, 6, -5, 1, 4, -7, -9,
    -- layer=1 filter=118 channel=113
    -2, -2, 1, -8, -8, 4, 3, -13, -11,
    -- layer=1 filter=118 channel=114
    -11, -3, -2, 0, 2, 8, -2, 3, -3,
    -- layer=1 filter=118 channel=115
    1, 0, 8, 0, 5, 0, 0, -9, 0,
    -- layer=1 filter=118 channel=116
    11, -9, 9, 6, -7, -10, 2, -8, -9,
    -- layer=1 filter=118 channel=117
    7, 1, -10, 6, 0, -8, -4, 6, -3,
    -- layer=1 filter=118 channel=118
    8, 1, 5, 8, -2, 2, 7, -3, -2,
    -- layer=1 filter=118 channel=119
    -10, -3, -9, -5, 2, 5, 10, -1, 1,
    -- layer=1 filter=118 channel=120
    -12, 0, 6, -7, 3, -6, -7, -7, -12,
    -- layer=1 filter=118 channel=121
    -4, 0, -4, -10, 4, -7, 2, -4, -12,
    -- layer=1 filter=118 channel=122
    -6, -4, 8, -4, -8, 1, -8, 2, -10,
    -- layer=1 filter=118 channel=123
    5, 3, -12, 5, -9, 0, 4, -4, -3,
    -- layer=1 filter=118 channel=124
    0, -2, -12, -11, 1, -12, 3, -3, 0,
    -- layer=1 filter=118 channel=125
    -1, -4, -7, -10, 2, 8, 1, -3, 1,
    -- layer=1 filter=118 channel=126
    -2, 7, 3, 7, -9, -11, -4, 0, -4,
    -- layer=1 filter=118 channel=127
    -11, -5, -9, -6, 4, -1, 3, 2, -10,
    -- layer=1 filter=119 channel=0
    7, -5, -11, 7, -10, -1, 4, -3, 1,
    -- layer=1 filter=119 channel=1
    -9, -6, -9, -4, 8, 6, 5, -8, 0,
    -- layer=1 filter=119 channel=2
    -1, -1, -10, 8, 0, -8, -10, -7, -13,
    -- layer=1 filter=119 channel=3
    -10, -6, 4, 7, -6, -8, -7, -1, -6,
    -- layer=1 filter=119 channel=4
    -4, -6, 5, 3, 0, 0, 5, -11, 1,
    -- layer=1 filter=119 channel=5
    8, -5, -7, -7, -3, -3, 0, -6, 2,
    -- layer=1 filter=119 channel=6
    0, -4, -1, -9, 5, 4, -1, 6, -10,
    -- layer=1 filter=119 channel=7
    10, -8, 0, 0, -9, 4, -5, -4, -7,
    -- layer=1 filter=119 channel=8
    10, 9, -5, -7, -6, 4, 7, 10, -7,
    -- layer=1 filter=119 channel=9
    -8, 1, -8, 6, -5, -4, 2, -5, -8,
    -- layer=1 filter=119 channel=10
    6, -5, 0, 7, -8, -12, -3, -7, -13,
    -- layer=1 filter=119 channel=11
    -4, -1, -7, 0, 0, -12, -2, -3, -2,
    -- layer=1 filter=119 channel=12
    -9, 3, -6, 3, 0, 1, -1, -9, 0,
    -- layer=1 filter=119 channel=13
    -2, 9, -8, 2, 6, -5, 1, 0, 9,
    -- layer=1 filter=119 channel=14
    1, -9, -7, 0, -1, -7, 6, -11, -11,
    -- layer=1 filter=119 channel=15
    -6, -10, 6, 3, -6, -5, -3, 8, -6,
    -- layer=1 filter=119 channel=16
    8, 2, 10, 1, 2, 3, -2, 0, 1,
    -- layer=1 filter=119 channel=17
    8, -11, 3, 0, -11, -9, 6, -8, -11,
    -- layer=1 filter=119 channel=18
    -4, -3, 5, 5, -6, -11, 0, -6, 8,
    -- layer=1 filter=119 channel=19
    -10, -7, 3, -9, 8, 6, -10, 7, 6,
    -- layer=1 filter=119 channel=20
    -4, -3, -10, -1, -2, -11, 0, 8, 7,
    -- layer=1 filter=119 channel=21
    0, -5, -3, -12, 2, 9, 0, -6, -10,
    -- layer=1 filter=119 channel=22
    -8, -10, 4, -2, -1, -8, 1, 0, -10,
    -- layer=1 filter=119 channel=23
    4, -12, -4, -4, -1, -12, 0, -12, -11,
    -- layer=1 filter=119 channel=24
    1, 8, 2, 0, 5, -12, 0, 7, -4,
    -- layer=1 filter=119 channel=25
    -2, 3, -2, 2, -10, 0, -5, -11, 5,
    -- layer=1 filter=119 channel=26
    2, -2, -12, 0, 7, 0, -7, 3, -3,
    -- layer=1 filter=119 channel=27
    6, 5, -4, -1, 0, 4, -9, -3, 9,
    -- layer=1 filter=119 channel=28
    6, 6, -3, 1, 5, 0, -9, 3, -6,
    -- layer=1 filter=119 channel=29
    -7, -6, -1, -3, 10, 7, -2, 6, -5,
    -- layer=1 filter=119 channel=30
    5, 12, 2, -4, 6, 5, 4, -7, -9,
    -- layer=1 filter=119 channel=31
    6, -7, 0, 6, 1, 6, -5, -10, -5,
    -- layer=1 filter=119 channel=32
    1, 4, 3, -3, -1, 0, -6, 6, 7,
    -- layer=1 filter=119 channel=33
    -2, -8, -2, 2, 5, -11, -2, 6, -5,
    -- layer=1 filter=119 channel=34
    -5, 6, -10, -11, -8, 6, -5, -8, -7,
    -- layer=1 filter=119 channel=35
    0, -3, 0, -9, 4, -10, -2, 8, 10,
    -- layer=1 filter=119 channel=36
    -8, -11, -3, -6, -1, -10, -8, -10, -8,
    -- layer=1 filter=119 channel=37
    -10, 0, 2, -3, 4, -12, -7, -4, 0,
    -- layer=1 filter=119 channel=38
    -7, -8, 8, 0, -13, 0, 7, 3, -8,
    -- layer=1 filter=119 channel=39
    3, -11, -3, 0, -11, -6, -8, 0, 6,
    -- layer=1 filter=119 channel=40
    -9, -10, 4, -3, 1, 8, -2, -6, -13,
    -- layer=1 filter=119 channel=41
    2, 10, -5, -14, 6, 2, -8, 0, -9,
    -- layer=1 filter=119 channel=42
    7, -7, -7, 0, 0, -9, 1, 6, -2,
    -- layer=1 filter=119 channel=43
    -8, -11, -11, -2, 8, -12, 8, -3, -8,
    -- layer=1 filter=119 channel=44
    -14, -1, -8, -8, -2, 7, 7, -6, -11,
    -- layer=1 filter=119 channel=45
    -7, 7, 4, -11, -10, 7, -10, -3, 8,
    -- layer=1 filter=119 channel=46
    3, -8, -4, -5, 4, -3, 6, 3, -6,
    -- layer=1 filter=119 channel=47
    4, 8, 1, -7, 2, -3, 5, -7, -10,
    -- layer=1 filter=119 channel=48
    4, -6, 0, -3, 4, -12, 0, -4, 5,
    -- layer=1 filter=119 channel=49
    -5, 4, -10, 7, 4, -11, -9, -4, -12,
    -- layer=1 filter=119 channel=50
    -4, -11, 0, 11, -8, 5, 0, -7, 4,
    -- layer=1 filter=119 channel=51
    4, -13, -8, -7, 7, -7, -10, -9, 0,
    -- layer=1 filter=119 channel=52
    -5, -3, 8, 5, 3, 4, 7, -9, 9,
    -- layer=1 filter=119 channel=53
    -6, -2, 2, -9, -12, 2, -5, 0, -11,
    -- layer=1 filter=119 channel=54
    3, 0, -3, 5, -4, -2, -9, 0, 4,
    -- layer=1 filter=119 channel=55
    -7, 0, -1, -7, -6, -7, -10, -8, -4,
    -- layer=1 filter=119 channel=56
    0, -4, 4, 3, 8, 7, 6, -8, 0,
    -- layer=1 filter=119 channel=57
    8, 2, -10, 0, -1, -1, -2, 6, -5,
    -- layer=1 filter=119 channel=58
    -9, -9, -5, 0, -5, -10, 7, -5, -4,
    -- layer=1 filter=119 channel=59
    -3, 0, 5, 7, -8, -9, 3, 8, -12,
    -- layer=1 filter=119 channel=60
    0, -8, 3, -6, -9, 9, 7, 3, 7,
    -- layer=1 filter=119 channel=61
    1, -2, -8, -2, 8, -7, 4, -6, 1,
    -- layer=1 filter=119 channel=62
    0, 0, 11, 9, -2, -8, 5, -3, 5,
    -- layer=1 filter=119 channel=63
    7, -6, 2, -2, 9, -6, -6, -2, -2,
    -- layer=1 filter=119 channel=64
    -8, -11, 3, 4, 2, -10, 2, -12, -12,
    -- layer=1 filter=119 channel=65
    2, 0, 4, -6, 0, -7, -5, 0, 0,
    -- layer=1 filter=119 channel=66
    5, -9, 3, -10, 3, 0, 4, -10, 5,
    -- layer=1 filter=119 channel=67
    -9, -4, 0, -2, 9, 8, 0, -1, 2,
    -- layer=1 filter=119 channel=68
    -12, 7, -2, 4, -5, -9, 2, 7, -1,
    -- layer=1 filter=119 channel=69
    -7, -9, 0, -2, 3, 4, -13, -2, -4,
    -- layer=1 filter=119 channel=70
    2, 9, 1, -4, -9, 7, -3, 0, -2,
    -- layer=1 filter=119 channel=71
    -5, 4, -3, 1, 3, 0, 4, -2, 1,
    -- layer=1 filter=119 channel=72
    -9, 1, 5, 4, -12, 1, 9, -11, -1,
    -- layer=1 filter=119 channel=73
    4, 4, -3, 4, 8, -6, -8, 4, -10,
    -- layer=1 filter=119 channel=74
    -7, 5, -2, -1, -11, 7, -8, -9, -9,
    -- layer=1 filter=119 channel=75
    -9, -9, -1, 5, -2, -4, -8, -7, 6,
    -- layer=1 filter=119 channel=76
    0, -7, -13, 0, -11, 6, -5, -7, 3,
    -- layer=1 filter=119 channel=77
    4, 7, -8, -3, -8, 4, 4, 7, 5,
    -- layer=1 filter=119 channel=78
    5, -2, 7, 3, -6, -6, 0, 7, 0,
    -- layer=1 filter=119 channel=79
    2, 6, 9, 5, -11, -9, -3, -7, 1,
    -- layer=1 filter=119 channel=80
    6, 8, -8, 3, -8, 3, 7, 4, 0,
    -- layer=1 filter=119 channel=81
    4, -5, -8, 7, -9, 2, -8, -3, 1,
    -- layer=1 filter=119 channel=82
    1, 2, -6, -3, 8, -8, -5, 0, -8,
    -- layer=1 filter=119 channel=83
    -11, -10, -12, 3, -7, 2, -4, 4, 5,
    -- layer=1 filter=119 channel=84
    -2, 6, -7, 1, -6, 1, -3, -7, 0,
    -- layer=1 filter=119 channel=85
    -3, 1, 3, -5, 1, -2, -8, 6, 7,
    -- layer=1 filter=119 channel=86
    10, -7, 2, 0, -12, -2, 1, -6, 6,
    -- layer=1 filter=119 channel=87
    -5, 6, 5, 7, -11, 7, -6, -10, -3,
    -- layer=1 filter=119 channel=88
    -7, -6, -11, -3, 8, -3, -8, 6, 6,
    -- layer=1 filter=119 channel=89
    -3, -10, 1, -6, 4, -3, 6, -10, -4,
    -- layer=1 filter=119 channel=90
    -4, 0, -3, -14, 5, 1, -12, -2, -7,
    -- layer=1 filter=119 channel=91
    -5, -11, -8, 3, -3, -3, 5, 7, 1,
    -- layer=1 filter=119 channel=92
    2, 5, 0, -6, 4, 3, 1, 0, -6,
    -- layer=1 filter=119 channel=93
    -9, -7, 0, 7, -5, -8, -4, -8, -7,
    -- layer=1 filter=119 channel=94
    -6, 2, 3, 7, -9, -9, -7, 0, 6,
    -- layer=1 filter=119 channel=95
    -10, 8, 4, -13, -4, 6, -2, 0, 3,
    -- layer=1 filter=119 channel=96
    4, -4, -11, -4, 6, -3, 8, -7, -1,
    -- layer=1 filter=119 channel=97
    -8, 7, -2, 4, 8, 3, -10, 2, 7,
    -- layer=1 filter=119 channel=98
    2, -7, 0, -5, -8, -4, -8, -10, -5,
    -- layer=1 filter=119 channel=99
    1, 3, 0, 5, -10, -10, -12, 6, -3,
    -- layer=1 filter=119 channel=100
    -1, -5, -10, 6, -13, 6, -6, -6, -8,
    -- layer=1 filter=119 channel=101
    -3, -6, 6, 0, -7, 3, -9, -1, -7,
    -- layer=1 filter=119 channel=102
    4, 0, -8, 3, 0, -2, 0, -6, -5,
    -- layer=1 filter=119 channel=103
    -3, -1, 1, 6, -9, -10, 5, 0, 3,
    -- layer=1 filter=119 channel=104
    -4, -9, 5, 3, 6, -12, 7, 4, -4,
    -- layer=1 filter=119 channel=105
    8, -6, -5, 4, -1, 6, -1, 2, -4,
    -- layer=1 filter=119 channel=106
    -7, -7, -4, 1, -6, 7, -6, -5, -7,
    -- layer=1 filter=119 channel=107
    -8, 3, 7, -7, -1, 8, -8, -2, -8,
    -- layer=1 filter=119 channel=108
    4, -4, 0, -6, 0, -8, 1, -5, -6,
    -- layer=1 filter=119 channel=109
    7, -4, -10, 1, 1, -4, 2, 5, 4,
    -- layer=1 filter=119 channel=110
    -9, -5, -4, 8, -12, 2, -7, 9, 4,
    -- layer=1 filter=119 channel=111
    4, -9, 5, -5, -11, -1, -5, 3, 3,
    -- layer=1 filter=119 channel=112
    -6, -1, -10, 7, -6, -11, 1, -11, -1,
    -- layer=1 filter=119 channel=113
    3, -12, -9, 7, -4, 3, -2, -8, -5,
    -- layer=1 filter=119 channel=114
    1, -10, 4, -7, 5, -9, -5, -3, 8,
    -- layer=1 filter=119 channel=115
    -9, 4, -9, -6, -9, -4, 6, -8, 1,
    -- layer=1 filter=119 channel=116
    -3, -5, 0, 4, -9, 3, -9, 0, -5,
    -- layer=1 filter=119 channel=117
    -4, -7, 6, -5, -1, -7, -7, -2, 6,
    -- layer=1 filter=119 channel=118
    -7, -4, -1, 5, 5, -8, 3, -9, 9,
    -- layer=1 filter=119 channel=119
    4, -4, -4, -5, -4, -1, 0, -5, -3,
    -- layer=1 filter=119 channel=120
    0, -12, 5, -12, 7, -1, 5, 3, 3,
    -- layer=1 filter=119 channel=121
    -12, -8, 6, -2, -13, 1, 0, 0, -4,
    -- layer=1 filter=119 channel=122
    -9, 0, -5, 1, -4, -3, -9, -7, -6,
    -- layer=1 filter=119 channel=123
    -5, -7, 4, -7, 2, -5, -6, -4, -3,
    -- layer=1 filter=119 channel=124
    5, -1, -10, -3, 1, -12, 1, -5, 8,
    -- layer=1 filter=119 channel=125
    0, -6, -1, 0, -6, -11, -7, 1, 0,
    -- layer=1 filter=119 channel=126
    3, 9, -2, 0, -3, -4, 3, 2, -7,
    -- layer=1 filter=119 channel=127
    -7, 0, -7, -14, -8, 5, -5, -7, 6,
    -- layer=1 filter=120 channel=0
    -14, -22, -23, -4, -9, -11, 19, 18, 10,
    -- layer=1 filter=120 channel=1
    12, -25, -17, 32, 17, -8, 20, 16, 2,
    -- layer=1 filter=120 channel=2
    -8, -4, 7, -4, 23, 12, 15, 5, -9,
    -- layer=1 filter=120 channel=3
    8, -3, -8, -3, 2, -8, 0, -9, -15,
    -- layer=1 filter=120 channel=4
    0, 5, -2, -10, -10, 3, 10, -11, 0,
    -- layer=1 filter=120 channel=5
    40, -2, 19, 23, 20, 12, 19, 34, 28,
    -- layer=1 filter=120 channel=6
    -57, -77, -44, -58, -69, -92, -51, -50, -57,
    -- layer=1 filter=120 channel=7
    6, 11, -5, -21, -17, -25, -32, -49, -45,
    -- layer=1 filter=120 channel=8
    27, -17, 21, 37, 36, 18, 49, 32, 19,
    -- layer=1 filter=120 channel=9
    -2, -48, 8, -17, -10, -10, -33, -18, -21,
    -- layer=1 filter=120 channel=10
    16, -5, 15, -10, -16, -17, -20, -42, -32,
    -- layer=1 filter=120 channel=11
    -21, -12, -1, -5, -24, -8, -8, 0, 14,
    -- layer=1 filter=120 channel=12
    -5, -64, -52, -31, -41, -50, -20, 32, -6,
    -- layer=1 filter=120 channel=13
    -16, -18, -20, -7, -18, -21, 20, 18, -2,
    -- layer=1 filter=120 channel=14
    -1, 24, 6, 7, 1, 5, -16, 7, -30,
    -- layer=1 filter=120 channel=15
    23, 3, 5, 0, 18, -25, -2, 16, 6,
    -- layer=1 filter=120 channel=16
    27, 24, 25, 32, 23, 2, 36, 42, 27,
    -- layer=1 filter=120 channel=17
    -22, -23, -33, 23, 16, 10, 19, 23, 27,
    -- layer=1 filter=120 channel=18
    -11, -56, -9, -8, 4, -26, -17, -4, 1,
    -- layer=1 filter=120 channel=19
    24, 39, 68, 55, 59, 35, 51, 47, 37,
    -- layer=1 filter=120 channel=20
    -27, -15, -35, 6, 0, -11, 23, 26, 11,
    -- layer=1 filter=120 channel=21
    -6, -2, -13, 6, -1, 5, 13, 12, 26,
    -- layer=1 filter=120 channel=22
    -36, -58, -46, -6, 0, -13, 26, 34, 2,
    -- layer=1 filter=120 channel=23
    38, 57, 10, 22, 51, 3, -20, -9, 4,
    -- layer=1 filter=120 channel=24
    0, 6, 12, 9, -7, 0, 7, 14, 17,
    -- layer=1 filter=120 channel=25
    -3, 17, 23, 14, -12, -12, 6, 10, -10,
    -- layer=1 filter=120 channel=26
    19, 24, 22, 0, 12, -6, -25, 5, -20,
    -- layer=1 filter=120 channel=27
    -32, -31, -28, -52, -57, -52, -26, -24, -15,
    -- layer=1 filter=120 channel=28
    5, -4, 18, -7, -16, -22, 9, -1, -16,
    -- layer=1 filter=120 channel=29
    -2, -18, -5, -25, -23, 0, 10, 16, 34,
    -- layer=1 filter=120 channel=30
    2, -53, -4, 24, 10, 0, -1, 23, 15,
    -- layer=1 filter=120 channel=31
    -48, -75, -59, -30, -28, -32, -27, -23, -41,
    -- layer=1 filter=120 channel=32
    12, 25, 35, -20, 11, -18, -29, -28, -25,
    -- layer=1 filter=120 channel=33
    -36, -37, -40, -25, -32, -25, -17, -15, -16,
    -- layer=1 filter=120 channel=34
    -54, -32, 5, -6, -24, -2, -28, -28, -14,
    -- layer=1 filter=120 channel=35
    1, 5, 7, 2, 0, 11, 1, 22, 15,
    -- layer=1 filter=120 channel=36
    -8, -7, 7, -9, -13, 2, -4, 0, 15,
    -- layer=1 filter=120 channel=37
    25, 25, 29, 30, 22, 8, 31, 42, 19,
    -- layer=1 filter=120 channel=38
    -10, -21, -19, -2, -6, -26, 16, 18, 20,
    -- layer=1 filter=120 channel=39
    -8, -17, -10, 10, 3, 12, -5, 16, 10,
    -- layer=1 filter=120 channel=40
    -29, -47, -7, -21, -8, -49, -27, -30, -41,
    -- layer=1 filter=120 channel=41
    13, 15, 31, -38, 12, -3, -21, 3, -4,
    -- layer=1 filter=120 channel=42
    -16, -2, -7, 17, 32, 22, 14, -1, 0,
    -- layer=1 filter=120 channel=43
    10, 11, 19, 18, 3, -7, 11, 37, 0,
    -- layer=1 filter=120 channel=44
    19, 21, 34, 1, -9, -6, -6, -38, -1,
    -- layer=1 filter=120 channel=45
    13, -17, -4, 8, -2, -12, 11, 0, 6,
    -- layer=1 filter=120 channel=46
    23, 40, 32, 32, 9, 20, 48, 24, 23,
    -- layer=1 filter=120 channel=47
    29, 43, -8, -9, 34, -23, -57, -5, -18,
    -- layer=1 filter=120 channel=48
    -9, -16, -38, -17, -3, -12, 9, 14, 31,
    -- layer=1 filter=120 channel=49
    -4, -13, -30, -31, 0, -18, 1, 3, -5,
    -- layer=1 filter=120 channel=50
    -5, -18, 7, -13, -13, 3, 17, 1, 7,
    -- layer=1 filter=120 channel=51
    -12, -18, -17, -9, -1, -10, -2, 8, -3,
    -- layer=1 filter=120 channel=52
    12, -4, 10, 3, -5, 1, -7, 4, -13,
    -- layer=1 filter=120 channel=53
    9, 27, 0, 12, 1, -13, 20, 7, 11,
    -- layer=1 filter=120 channel=54
    8, 25, 30, 10, -3, -7, 14, 22, -8,
    -- layer=1 filter=120 channel=55
    10, 10, 4, -2, 4, 7, -5, 10, 18,
    -- layer=1 filter=120 channel=56
    4, 3, -7, 7, -10, 1, 8, 6, -14,
    -- layer=1 filter=120 channel=57
    -3, -23, 3, -23, -21, -10, -18, -22, -16,
    -- layer=1 filter=120 channel=58
    22, 30, -5, -11, 10, -4, -44, -41, -14,
    -- layer=1 filter=120 channel=59
    -5, -14, -15, -17, -12, -14, 15, 0, -8,
    -- layer=1 filter=120 channel=60
    29, 26, 5, 24, 16, 2, 21, 6, 1,
    -- layer=1 filter=120 channel=61
    0, -9, -11, 5, -7, -1, -1, -9, -7,
    -- layer=1 filter=120 channel=62
    20, 12, 30, 48, 33, 25, 50, 40, 20,
    -- layer=1 filter=120 channel=63
    -17, 4, -12, -21, -23, -2, -2, -7, 19,
    -- layer=1 filter=120 channel=64
    -25, -19, -23, -1, -9, -9, 10, 4, -3,
    -- layer=1 filter=120 channel=65
    -31, -27, -23, -14, -3, -8, 17, 20, 3,
    -- layer=1 filter=120 channel=66
    -5, -9, -18, -11, 0, 0, 14, 10, 22,
    -- layer=1 filter=120 channel=67
    -37, -45, -28, -53, -53, -38, -35, -6, -7,
    -- layer=1 filter=120 channel=68
    14, 28, 42, 3, -19, -11, -14, -45, -16,
    -- layer=1 filter=120 channel=69
    39, 25, 32, 5, 25, -12, 18, 41, 9,
    -- layer=1 filter=120 channel=70
    -24, -54, -59, -35, -18, -34, -42, -39, -59,
    -- layer=1 filter=120 channel=71
    -17, -6, 8, 7, 0, -7, 10, 4, 17,
    -- layer=1 filter=120 channel=72
    5, -30, 15, 6, 0, -9, 6, 15, -28,
    -- layer=1 filter=120 channel=73
    -17, -13, -11, -8, 4, 3, -13, -9, 2,
    -- layer=1 filter=120 channel=74
    0, -12, 4, -10, -24, -37, -10, -28, -31,
    -- layer=1 filter=120 channel=75
    -28, -40, -25, -8, -15, 4, -24, 27, -13,
    -- layer=1 filter=120 channel=76
    -6, 9, 18, 0, -14, 0, -6, 17, 8,
    -- layer=1 filter=120 channel=77
    -10, -22, -12, -10, 1, 5, 22, 15, 14,
    -- layer=1 filter=120 channel=78
    2, 3, 7, -13, -11, -17, 5, 2, 2,
    -- layer=1 filter=120 channel=79
    8, 12, 16, 16, 24, 9, 31, 40, 14,
    -- layer=1 filter=120 channel=80
    -10, 0, -1, 9, 5, 15, 17, 7, 18,
    -- layer=1 filter=120 channel=81
    -2, -12, -2, 1, 12, 23, 19, 13, 5,
    -- layer=1 filter=120 channel=82
    -15, -30, -31, -2, 1, -10, 10, 23, 18,
    -- layer=1 filter=120 channel=83
    12, -10, -4, 13, 7, -5, 8, 5, -5,
    -- layer=1 filter=120 channel=84
    0, -11, 1, 18, -8, -32, -48, -24, -33,
    -- layer=1 filter=120 channel=85
    33, 33, 9, -14, 23, -6, -67, -17, -12,
    -- layer=1 filter=120 channel=86
    -6, -9, -9, 1, 6, 17, 12, 16, 26,
    -- layer=1 filter=120 channel=87
    0, -2, -4, 19, 11, 28, 59, 26, 19,
    -- layer=1 filter=120 channel=88
    -27, -4, -30, -19, -9, 0, 4, 16, 0,
    -- layer=1 filter=120 channel=89
    -18, -19, -19, -14, -7, 0, 16, 22, 4,
    -- layer=1 filter=120 channel=90
    16, 20, 14, 0, 9, 4, 5, -3, -5,
    -- layer=1 filter=120 channel=91
    -24, -24, -34, -20, -13, -28, 4, 6, 1,
    -- layer=1 filter=120 channel=92
    -35, 15, -15, -23, -1, -36, 32, -8, -1,
    -- layer=1 filter=120 channel=93
    -8, -18, -3, -3, 1, -2, 18, 20, 13,
    -- layer=1 filter=120 channel=94
    -10, -17, -21, 2, -11, -7, 14, 12, 12,
    -- layer=1 filter=120 channel=95
    -23, -36, 3, 8, 7, -2, -14, 1, -13,
    -- layer=1 filter=120 channel=96
    -10, -13, -2, -1, -3, 3, 7, -10, -3,
    -- layer=1 filter=120 channel=97
    -16, -13, -16, 1, 12, 9, 19, 21, 13,
    -- layer=1 filter=120 channel=98
    -12, -28, 0, 31, 3, 18, 32, 30, 6,
    -- layer=1 filter=120 channel=99
    64, 34, 49, 30, 12, -11, 26, -15, -46,
    -- layer=1 filter=120 channel=100
    -19, -22, 0, -18, -17, -15, 2, 2, 0,
    -- layer=1 filter=120 channel=101
    -15, -35, -40, -9, -7, -16, 18, 15, -5,
    -- layer=1 filter=120 channel=102
    -7, -30, -15, -3, -19, -10, 21, 19, 21,
    -- layer=1 filter=120 channel=103
    -22, -47, -14, -10, -42, -32, -28, -21, -8,
    -- layer=1 filter=120 channel=104
    26, 11, 13, -2, 18, 1, -35, 13, 15,
    -- layer=1 filter=120 channel=105
    -17, -17, -16, -6, -2, 3, 21, 2, 19,
    -- layer=1 filter=120 channel=106
    -10, -12, -17, -14, 0, -20, -6, -7, 5,
    -- layer=1 filter=120 channel=107
    -23, -11, -19, 1, -21, -24, -9, -15, -18,
    -- layer=1 filter=120 channel=108
    19, 25, 20, -25, 20, -3, -1, -19, -21,
    -- layer=1 filter=120 channel=109
    -1, -5, -4, -4, 8, -3, -5, 0, -5,
    -- layer=1 filter=120 channel=110
    -6, -24, -21, -4, -11, 2, 5, 17, 1,
    -- layer=1 filter=120 channel=111
    15, -50, -12, 24, 26, -10, 2, 2, 5,
    -- layer=1 filter=120 channel=112
    -22, -39, -22, 23, 10, 10, -14, 8, 7,
    -- layer=1 filter=120 channel=113
    -58, -16, -20, -28, -9, -13, -2, -4, 12,
    -- layer=1 filter=120 channel=114
    43, 18, 38, 23, 31, 3, 20, 43, 36,
    -- layer=1 filter=120 channel=115
    -25, -9, -3, -12, -1, 7, 29, 15, 12,
    -- layer=1 filter=120 channel=116
    0, 4, 8, 7, 0, 9, -5, 2, 10,
    -- layer=1 filter=120 channel=117
    38, -8, 2, 48, 46, 32, 26, 17, 41,
    -- layer=1 filter=120 channel=118
    -15, -33, 7, 13, -5, -28, -15, -10, -18,
    -- layer=1 filter=120 channel=119
    6, 24, 42, -17, -2, -24, -40, -17, -32,
    -- layer=1 filter=120 channel=120
    -7, -15, -20, 3, -3, 1, 2, 15, 1,
    -- layer=1 filter=120 channel=121
    15, 2, 6, 18, 28, 36, 35, 22, 8,
    -- layer=1 filter=120 channel=122
    7, 1, -3, -9, -7, -10, 1, -8, 0,
    -- layer=1 filter=120 channel=123
    -3, 2, 9, -6, -2, 22, -5, 0, -2,
    -- layer=1 filter=120 channel=124
    9, -7, 0, 14, 7, 0, 8, 19, 11,
    -- layer=1 filter=120 channel=125
    4, -25, -36, 0, 11, -13, -54, -46, -16,
    -- layer=1 filter=120 channel=126
    13, -12, 18, 60, 47, 30, 40, 38, 5,
    -- layer=1 filter=120 channel=127
    -31, -48, -6, 12, 14, -9, -1, 11, -9,
    -- layer=1 filter=121 channel=0
    2, 9, -1, -11, 1, 7, -4, -10, -10,
    -- layer=1 filter=121 channel=1
    -23, -34, -24, -49, -44, -38, -3, 7, 14,
    -- layer=1 filter=121 channel=2
    -44, -27, 0, -2, 14, 17, -16, 18, 32,
    -- layer=1 filter=121 channel=3
    -4, 8, 3, 8, 9, 8, 4, 11, 10,
    -- layer=1 filter=121 channel=4
    6, 6, 2, -6, 0, 9, -3, 0, 7,
    -- layer=1 filter=121 channel=5
    -81, -111, -67, -101, -126, -84, 21, 26, 29,
    -- layer=1 filter=121 channel=6
    -9, 1, -19, 0, -1, -5, -3, -10, 3,
    -- layer=1 filter=121 channel=7
    -10, -110, -112, -24, -154, -159, -40, -133, -112,
    -- layer=1 filter=121 channel=8
    -70, -140, -63, -120, -136, -140, 5, 28, 35,
    -- layer=1 filter=121 channel=9
    -11, -16, -7, -39, 0, -24, 10, -45, 4,
    -- layer=1 filter=121 channel=10
    -5, -78, -115, -4, -130, -142, -15, -113, -82,
    -- layer=1 filter=121 channel=11
    10, 14, 10, 16, 15, -15, -3, -17, -22,
    -- layer=1 filter=121 channel=12
    -24, -25, -28, -18, -48, -2, 12, -20, 24,
    -- layer=1 filter=121 channel=13
    -4, 23, 10, 0, -4, 12, 4, 1, -2,
    -- layer=1 filter=121 channel=14
    -23, -44, -22, -26, -36, -35, -45, -46, -71,
    -- layer=1 filter=121 channel=15
    -50, -13, -34, -23, -61, -62, -21, -5, -3,
    -- layer=1 filter=121 channel=16
    -60, -106, -62, -68, -106, -82, 24, 33, 29,
    -- layer=1 filter=121 channel=17
    9, 8, 0, -15, 0, -16, -2, -9, -6,
    -- layer=1 filter=121 channel=18
    13, -3, 10, 3, -10, 10, -9, -24, -1,
    -- layer=1 filter=121 channel=19
    -68, -51, -65, -40, -57, -15, 21, 20, 35,
    -- layer=1 filter=121 channel=20
    3, 21, 13, 2, 0, -8, 11, 8, 7,
    -- layer=1 filter=121 channel=21
    -5, -15, -7, 6, 12, 8, 26, 23, 29,
    -- layer=1 filter=121 channel=22
    8, -5, 15, -26, -10, -16, -20, -14, 0,
    -- layer=1 filter=121 channel=23
    -26, -46, -18, -47, -57, -43, -18, -65, 0,
    -- layer=1 filter=121 channel=24
    -1, 0, 15, 12, 27, 31, 52, 59, 47,
    -- layer=1 filter=121 channel=25
    -24, -81, -120, -33, -141, -134, -4, -57, -37,
    -- layer=1 filter=121 channel=26
    32, 27, 23, -10, 12, 13, -8, 15, -5,
    -- layer=1 filter=121 channel=27
    -8, -1, -30, -8, -7, -27, 14, 0, -3,
    -- layer=1 filter=121 channel=28
    0, -35, -43, 6, -61, -68, -11, -58, -48,
    -- layer=1 filter=121 channel=29
    -9, -20, -33, -1, -6, -8, -18, -11, -6,
    -- layer=1 filter=121 channel=30
    19, -16, -19, -5, -8, 12, 14, -39, -14,
    -- layer=1 filter=121 channel=31
    -19, -22, -44, 16, -7, 20, 36, 12, 10,
    -- layer=1 filter=121 channel=32
    39, 1, 14, -1, -2, 10, -31, -13, 13,
    -- layer=1 filter=121 channel=33
    8, 6, 2, -3, 14, 16, -7, -7, -9,
    -- layer=1 filter=121 channel=34
    -18, -19, 3, -26, -26, 7, -12, -21, -21,
    -- layer=1 filter=121 channel=35
    -16, -8, -13, 1, -10, -8, -6, -9, -7,
    -- layer=1 filter=121 channel=36
    35, 9, 5, 28, 2, 2, -1, -2, -10,
    -- layer=1 filter=121 channel=37
    -110, -109, -79, -100, -112, -93, 22, 39, 41,
    -- layer=1 filter=121 channel=38
    16, 6, 19, 8, 21, 0, 24, 13, 1,
    -- layer=1 filter=121 channel=39
    -30, -20, -28, -26, -25, -23, -2, -2, -12,
    -- layer=1 filter=121 channel=40
    -16, -24, -16, 1, 0, 3, 8, 1, 0,
    -- layer=1 filter=121 channel=41
    53, 7, -39, 27, -35, 10, 55, -36, 33,
    -- layer=1 filter=121 channel=42
    -31, -36, 2, -10, 7, 34, -24, -20, 10,
    -- layer=1 filter=121 channel=43
    -42, -76, -82, -68, -76, -69, 11, 12, 15,
    -- layer=1 filter=121 channel=44
    -9, 6, 13, -12, 3, 12, -44, -14, -5,
    -- layer=1 filter=121 channel=45
    -2, -10, 18, -4, 10, 1, 0, 35, 28,
    -- layer=1 filter=121 channel=46
    -95, -86, -78, -62, -46, 7, 42, 71, 62,
    -- layer=1 filter=121 channel=47
    -7, -40, -34, -42, -53, 3, -9, -30, 32,
    -- layer=1 filter=121 channel=48
    13, 4, -5, 4, 0, 12, 14, 9, 3,
    -- layer=1 filter=121 channel=49
    -21, -17, -3, -11, 1, 13, -3, -1, 23,
    -- layer=1 filter=121 channel=50
    0, -1, 3, -10, 0, -7, 8, -7, 10,
    -- layer=1 filter=121 channel=51
    6, -14, -14, 9, 5, -1, 0, 17, 2,
    -- layer=1 filter=121 channel=52
    -2, 0, 6, 3, 4, 5, -8, 0, 0,
    -- layer=1 filter=121 channel=53
    -3, -2, 1, -3, -14, -9, -16, -11, -16,
    -- layer=1 filter=121 channel=54
    -74, -60, -89, -10, -109, -79, 12, -19, -7,
    -- layer=1 filter=121 channel=55
    13, -3, 15, 28, 16, 9, 17, 27, 9,
    -- layer=1 filter=121 channel=56
    -10, -4, -3, -10, -4, -7, 0, -13, -3,
    -- layer=1 filter=121 channel=57
    -25, -67, -75, 5, -77, -73, -15, -98, -50,
    -- layer=1 filter=121 channel=58
    -69, -119, -129, -59, -117, -104, -11, -82, -46,
    -- layer=1 filter=121 channel=59
    0, -3, -12, 2, 1, -14, 0, -11, 0,
    -- layer=1 filter=121 channel=60
    -12, 1, -15, 3, 0, 0, -21, -10, -12,
    -- layer=1 filter=121 channel=61
    -10, 0, -5, -5, 9, -1, 5, -1, -11,
    -- layer=1 filter=121 channel=62
    -102, -132, -85, -109, -143, -120, 0, 16, 1,
    -- layer=1 filter=121 channel=63
    27, 17, 1, 9, 0, 5, 1, -13, -17,
    -- layer=1 filter=121 channel=64
    -5, 8, 7, -7, 0, -11, 2, -1, -13,
    -- layer=1 filter=121 channel=65
    17, 11, 9, 10, 7, -6, 23, 13, 3,
    -- layer=1 filter=121 channel=66
    15, 2, -4, 4, 3, 1, 1, -13, -4,
    -- layer=1 filter=121 channel=67
    13, 0, 9, -1, 17, 7, 28, 7, 0,
    -- layer=1 filter=121 channel=68
    -7, 22, 31, -8, 14, 11, -21, 8, -10,
    -- layer=1 filter=121 channel=69
    -38, -59, -31, -37, -67, -50, 18, 40, 28,
    -- layer=1 filter=121 channel=70
    -51, -51, -36, -16, -20, 0, 12, -19, -1,
    -- layer=1 filter=121 channel=71
    -3, 2, -12, 20, 7, 14, 39, 46, 38,
    -- layer=1 filter=121 channel=72
    13, -2, -22, -32, -46, -18, 8, -58, -16,
    -- layer=1 filter=121 channel=73
    4, 0, 5, 2, 4, -4, 6, 3, -10,
    -- layer=1 filter=121 channel=74
    7, 10, 0, 6, 18, 16, -12, -1, -50,
    -- layer=1 filter=121 channel=75
    -33, -1, -27, -29, -42, -27, -21, -30, -19,
    -- layer=1 filter=121 channel=76
    16, 10, -1, 1, -8, -12, -15, -14, -33,
    -- layer=1 filter=121 channel=77
    -4, -7, 6, 7, 9, 5, 21, 37, 23,
    -- layer=1 filter=121 channel=78
    7, 6, -8, 11, -8, 2, -2, -5, -6,
    -- layer=1 filter=121 channel=79
    -58, -71, -49, -76, -109, -95, 7, 23, 25,
    -- layer=1 filter=121 channel=80
    1, 7, -1, -3, 6, 8, -1, 9, 7,
    -- layer=1 filter=121 channel=81
    -18, -12, -10, 4, 7, 11, 41, 44, 33,
    -- layer=1 filter=121 channel=82
    -13, -4, 9, -2, 13, 14, 16, 18, 9,
    -- layer=1 filter=121 channel=83
    -30, -23, -24, -4, -37, -43, 3, -2, 4,
    -- layer=1 filter=121 channel=84
    29, 6, 21, -2, 11, 34, -1, -18, -10,
    -- layer=1 filter=121 channel=85
    -22, -25, -16, -35, -44, -29, 1, -58, -14,
    -- layer=1 filter=121 channel=86
    16, 21, 2, 14, 4, -3, 11, 3, 0,
    -- layer=1 filter=121 channel=87
    -33, -22, -32, -29, -8, -27, 72, 3, 28,
    -- layer=1 filter=121 channel=88
    -26, -11, -13, -14, -11, 8, 0, 2, 8,
    -- layer=1 filter=121 channel=89
    5, 19, 7, 6, 22, 18, 26, 30, 31,
    -- layer=1 filter=121 channel=90
    -16, -6, 2, -24, -20, -6, -29, 3, -12,
    -- layer=1 filter=121 channel=91
    19, 9, -1, 9, 19, 3, 10, -5, 0,
    -- layer=1 filter=121 channel=92
    12, -22, -44, 68, 26, -29, 16, -14, 0,
    -- layer=1 filter=121 channel=93
    5, 24, 9, 4, 6, 9, 31, 20, 10,
    -- layer=1 filter=121 channel=94
    21, 18, 4, 0, -4, -2, -3, -12, -14,
    -- layer=1 filter=121 channel=95
    12, 3, 10, -8, 0, 13, -28, -28, -12,
    -- layer=1 filter=121 channel=96
    5, -2, 2, 11, -7, 8, 9, 2, 3,
    -- layer=1 filter=121 channel=97
    24, 20, 10, 17, 7, -8, 13, -5, -13,
    -- layer=1 filter=121 channel=98
    -13, -45, -46, -54, -101, -111, -3, -20, -10,
    -- layer=1 filter=121 channel=99
    -1, -19, 4, 12, -24, -36, -11, -19, -38,
    -- layer=1 filter=121 channel=100
    14, 2, -1, 13, 7, -23, 2, -23, -4,
    -- layer=1 filter=121 channel=101
    9, 5, 12, 15, 6, 10, 14, 8, 2,
    -- layer=1 filter=121 channel=102
    17, 18, 1, 5, 13, 4, -7, -20, -15,
    -- layer=1 filter=121 channel=103
    12, 6, -1, 13, 13, -18, 0, -1, -4,
    -- layer=1 filter=121 channel=104
    8, -11, -25, -19, 6, 2, 5, -44, -10,
    -- layer=1 filter=121 channel=105
    9, 20, 18, 14, 13, 0, 11, 0, -14,
    -- layer=1 filter=121 channel=106
    16, 18, 21, 18, 20, 34, 2, 13, 9,
    -- layer=1 filter=121 channel=107
    3, 10, -2, 15, 9, 13, 11, 0, 14,
    -- layer=1 filter=121 channel=108
    -10, 0, 8, -17, -20, -6, -29, -7, 1,
    -- layer=1 filter=121 channel=109
    2, 0, 0, 8, -8, -7, 10, 8, 0,
    -- layer=1 filter=121 channel=110
    9, 6, -4, 1, 0, -14, 3, 2, -13,
    -- layer=1 filter=121 channel=111
    10, -11, 9, 7, 12, 32, -11, -19, -2,
    -- layer=1 filter=121 channel=112
    -32, -15, -7, 0, 3, 14, -37, 1, -20,
    -- layer=1 filter=121 channel=113
    -35, -33, -33, -28, -24, -17, -13, -42, -28,
    -- layer=1 filter=121 channel=114
    -90, -88, -85, -68, -47, -52, 18, 38, 17,
    -- layer=1 filter=121 channel=115
    24, -3, 12, 17, 8, 0, 8, -17, -1,
    -- layer=1 filter=121 channel=116
    5, 0, -3, -10, -4, 6, -5, 6, 0,
    -- layer=1 filter=121 channel=117
    -42, -66, -24, -30, -28, -10, -23, -18, -5,
    -- layer=1 filter=121 channel=118
    36, 13, 2, 5, 32, 26, 19, -12, 0,
    -- layer=1 filter=121 channel=119
    9, 0, 14, -14, -14, 15, -19, -13, -1,
    -- layer=1 filter=121 channel=120
    -12, -1, -4, -11, -8, -7, 18, 10, 10,
    -- layer=1 filter=121 channel=121
    -13, -4, -18, 12, -16, 12, 29, -3, 2,
    -- layer=1 filter=121 channel=122
    0, 8, -2, -6, -5, 0, 6, 5, -4,
    -- layer=1 filter=121 channel=123
    24, 10, 4, 8, 3, 20, 24, 2, 11,
    -- layer=1 filter=121 channel=124
    10, 0, -5, 6, -4, 1, 2, -6, 12,
    -- layer=1 filter=121 channel=125
    -60, -61, -27, -30, -29, -21, -2, -34, -4,
    -- layer=1 filter=121 channel=126
    -45, -71, -44, -80, -104, -92, -23, -33, -4,
    -- layer=1 filter=121 channel=127
    15, -3, -10, 13, 18, 32, -5, -17, -7,
    -- layer=1 filter=122 channel=0
    -8, 9, 3, 2, -7, -7, -5, -10, 1,
    -- layer=1 filter=122 channel=1
    60, 21, 4, -13, -5, -33, -47, -41, -39,
    -- layer=1 filter=122 channel=2
    -8, 0, -6, -38, -29, -64, 0, -33, -44,
    -- layer=1 filter=122 channel=3
    8, 6, 6, 3, 10, 10, 3, 11, 0,
    -- layer=1 filter=122 channel=4
    4, 5, 1, 7, 8, 6, 4, 7, 0,
    -- layer=1 filter=122 channel=5
    45, 12, 16, -40, -36, -39, -52, -29, -4,
    -- layer=1 filter=122 channel=6
    20, 15, 30, 22, 12, 19, -28, -25, -33,
    -- layer=1 filter=122 channel=7
    1, 9, 29, -36, -14, -17, -15, -29, 2,
    -- layer=1 filter=122 channel=8
    36, 3, -3, -10, -20, -27, -51, -22, -6,
    -- layer=1 filter=122 channel=9
    -16, -1, 8, -22, -41, -42, 2, -40, -11,
    -- layer=1 filter=122 channel=10
    -1, 17, 22, -27, -6, -12, -20, -29, 7,
    -- layer=1 filter=122 channel=11
    -9, -6, -8, 1, 14, 18, 14, 15, 0,
    -- layer=1 filter=122 channel=12
    -74, -30, -18, 15, -25, -21, -54, -23, -57,
    -- layer=1 filter=122 channel=13
    21, 40, 38, 0, -12, 4, -25, -27, -25,
    -- layer=1 filter=122 channel=14
    -33, 4, 39, -39, 15, -7, -26, -13, -11,
    -- layer=1 filter=122 channel=15
    -10, -8, -15, -63, -54, -48, -30, -37, -47,
    -- layer=1 filter=122 channel=16
    22, -12, -5, -34, -37, -18, -30, -29, 4,
    -- layer=1 filter=122 channel=17
    13, 19, 32, -2, -1, -6, -32, -17, -22,
    -- layer=1 filter=122 channel=18
    18, 24, 9, 28, 23, 28, 32, 25, 18,
    -- layer=1 filter=122 channel=19
    -21, -5, 8, -9, -23, -3, 26, 10, 18,
    -- layer=1 filter=122 channel=20
    26, 21, 26, -11, -3, -1, -46, -33, -26,
    -- layer=1 filter=122 channel=21
    15, 13, 6, -38, -28, -16, -58, -43, -62,
    -- layer=1 filter=122 channel=22
    29, 24, 34, 0, -7, -5, -32, -16, -23,
    -- layer=1 filter=122 channel=23
    -13, -19, -2, -62, -42, -47, -40, -55, -42,
    -- layer=1 filter=122 channel=24
    -14, -19, 9, -15, -35, -17, -13, -40, -13,
    -- layer=1 filter=122 channel=25
    22, -10, 8, -64, -60, -44, -12, -55, -4,
    -- layer=1 filter=122 channel=26
    13, 6, 25, -11, -10, 6, -7, -38, -10,
    -- layer=1 filter=122 channel=27
    -44, -42, -43, -27, -28, -29, -27, 0, -10,
    -- layer=1 filter=122 channel=28
    11, 19, 25, -41, -34, -11, -37, -33, -10,
    -- layer=1 filter=122 channel=29
    -20, -22, 0, 0, -8, -10, -23, -18, -16,
    -- layer=1 filter=122 channel=30
    26, 3, 14, 37, 34, 20, 34, 23, 15,
    -- layer=1 filter=122 channel=31
    2, -3, 5, 53, 33, 45, -1, 17, 3,
    -- layer=1 filter=122 channel=32
    -4, -20, 16, 15, -20, 2, 2, -32, -12,
    -- layer=1 filter=122 channel=33
    -5, 1, 5, -1, 0, 18, 0, -9, -1,
    -- layer=1 filter=122 channel=34
    -24, -19, -10, 18, -1, 3, -13, -1, 5,
    -- layer=1 filter=122 channel=35
    -3, -10, -10, -11, -20, -5, -1, -9, -10,
    -- layer=1 filter=122 channel=36
    7, -2, 3, 18, 23, 22, 6, 16, 25,
    -- layer=1 filter=122 channel=37
    28, 5, 23, -22, -28, 16, -16, -23, 4,
    -- layer=1 filter=122 channel=38
    31, 17, 28, -9, -7, 9, -19, -22, -12,
    -- layer=1 filter=122 channel=39
    -10, -13, 4, -2, -1, 4, -28, -12, 6,
    -- layer=1 filter=122 channel=40
    27, 11, 36, 19, 16, 31, -9, 13, -2,
    -- layer=1 filter=122 channel=41
    -4, -3, 0, -12, -64, -16, 23, -41, 0,
    -- layer=1 filter=122 channel=42
    -19, -29, -21, -10, -26, -32, -11, -28, -40,
    -- layer=1 filter=122 channel=43
    35, 2, -11, -18, -22, -14, -44, -14, -5,
    -- layer=1 filter=122 channel=44
    -13, -14, 17, -34, -44, 1, -16, -51, -26,
    -- layer=1 filter=122 channel=45
    15, -1, 16, -40, -30, -18, -55, -43, -22,
    -- layer=1 filter=122 channel=46
    -34, -51, 21, -24, -18, -3, 14, 7, 18,
    -- layer=1 filter=122 channel=47
    -19, -3, 4, -4, -38, -40, -20, -45, -26,
    -- layer=1 filter=122 channel=48
    22, 7, 25, -14, -19, -11, -39, -35, -34,
    -- layer=1 filter=122 channel=49
    -18, -2, -9, 4, 7, 0, -3, -38, -14,
    -- layer=1 filter=122 channel=50
    17, 8, 12, -5, -14, 2, -17, -9, -7,
    -- layer=1 filter=122 channel=51
    5, 30, 32, -33, 10, -1, -51, -25, -32,
    -- layer=1 filter=122 channel=52
    -13, -3, -3, 0, -6, 6, 0, 4, 0,
    -- layer=1 filter=122 channel=53
    0, -2, -17, -13, -12, -9, 5, -16, -4,
    -- layer=1 filter=122 channel=54
    11, -18, -9, -58, -47, -26, 11, -35, 21,
    -- layer=1 filter=122 channel=55
    -13, -26, -2, 15, 6, 7, 5, 19, 26,
    -- layer=1 filter=122 channel=56
    4, -5, 0, 7, 5, 2, 10, -3, 3,
    -- layer=1 filter=122 channel=57
    5, 25, 36, 0, 22, 9, -3, 3, 21,
    -- layer=1 filter=122 channel=58
    -55, 8, -17, -78, -58, -68, -27, -89, -5,
    -- layer=1 filter=122 channel=59
    5, -11, 0, 7, -3, -8, -4, -10, 6,
    -- layer=1 filter=122 channel=60
    -8, -6, -18, 2, 2, -19, 4, -12, 4,
    -- layer=1 filter=122 channel=61
    7, 6, 9, 0, 7, -4, 14, 12, -9,
    -- layer=1 filter=122 channel=62
    35, 3, -2, -19, -30, 2, -28, -25, -8,
    -- layer=1 filter=122 channel=63
    -11, 3, 1, 12, 9, 16, 8, 16, 0,
    -- layer=1 filter=122 channel=64
    0, 9, 18, 8, -11, 8, -12, -23, -8,
    -- layer=1 filter=122 channel=65
    4, 2, 25, -5, -15, 1, -23, -23, -18,
    -- layer=1 filter=122 channel=66
    -2, -8, 4, 0, 9, 5, -2, -4, -9,
    -- layer=1 filter=122 channel=67
    14, 29, -3, 35, 20, 48, -68, -70, -29,
    -- layer=1 filter=122 channel=68
    1, -20, 10, -26, -46, 7, -37, -66, -30,
    -- layer=1 filter=122 channel=69
    -7, -15, 0, -67, -61, -31, -38, -41, -33,
    -- layer=1 filter=122 channel=70
    -3, -20, -21, 40, 33, 43, -23, -11, -15,
    -- layer=1 filter=122 channel=71
    -10, -12, -7, -26, -12, -11, -11, -6, -25,
    -- layer=1 filter=122 channel=72
    -3, -17, 13, 0, -11, -18, 33, 17, 25,
    -- layer=1 filter=122 channel=73
    -5, 0, -9, 1, -2, -8, 5, -7, 0,
    -- layer=1 filter=122 channel=74
    33, -21, 0, 4, 15, 22, -11, -33, -6,
    -- layer=1 filter=122 channel=75
    -13, -19, 6, -6, -31, -24, 7, 3, -5,
    -- layer=1 filter=122 channel=76
    14, 0, 13, 0, 4, -2, 9, -14, -15,
    -- layer=1 filter=122 channel=77
    15, -2, 14, -16, -11, -21, -37, -33, -24,
    -- layer=1 filter=122 channel=78
    -6, 2, 7, -7, 6, 3, 0, -5, 9,
    -- layer=1 filter=122 channel=79
    12, -6, -3, -29, -45, -7, -20, -30, 1,
    -- layer=1 filter=122 channel=80
    5, 6, 8, 8, 0, 8, -1, 0, -5,
    -- layer=1 filter=122 channel=81
    -12, -27, -18, -9, -10, -17, -2, -21, -11,
    -- layer=1 filter=122 channel=82
    26, 14, 22, 1, -22, -5, -36, -43, -44,
    -- layer=1 filter=122 channel=83
    -5, -11, 1, -32, -16, -25, -38, -39, -26,
    -- layer=1 filter=122 channel=84
    45, 15, 30, 27, 11, 28, 32, 10, -8,
    -- layer=1 filter=122 channel=85
    -28, 4, 0, -34, -36, -47, -13, -51, -6,
    -- layer=1 filter=122 channel=86
    8, 15, 12, 7, 12, 8, -10, 2, 17,
    -- layer=1 filter=122 channel=87
    -33, -26, 23, 19, -12, -1, 22, 1, 21,
    -- layer=1 filter=122 channel=88
    -4, 0, -3, -12, -19, -25, -38, -28, -27,
    -- layer=1 filter=122 channel=89
    3, 22, 18, -5, -22, 2, -31, -31, -43,
    -- layer=1 filter=122 channel=90
    -38, -43, 10, -68, -98, -36, -66, -90, -34,
    -- layer=1 filter=122 channel=91
    26, 29, 34, 6, 0, 13, -17, -11, -23,
    -- layer=1 filter=122 channel=92
    -27, -76, -21, -104, -65, -28, -39, -72, -70,
    -- layer=1 filter=122 channel=93
    12, 7, 6, -7, -19, -20, -24, -15, -17,
    -- layer=1 filter=122 channel=94
    4, 16, 14, 2, 18, 10, -15, -7, 0,
    -- layer=1 filter=122 channel=95
    38, 8, 28, 30, 9, 41, 41, 28, 22,
    -- layer=1 filter=122 channel=96
    -2, 10, 14, 17, 0, 0, 1, 21, 5,
    -- layer=1 filter=122 channel=97
    -5, 10, 12, 0, -5, 4, -8, -18, -14,
    -- layer=1 filter=122 channel=98
    45, 0, -2, -14, -37, -14, -57, -31, -2,
    -- layer=1 filter=122 channel=99
    1, -9, 15, -50, -20, -28, -73, -49, -19,
    -- layer=1 filter=122 channel=100
    -10, -7, 2, -6, 11, 10, 5, 7, -9,
    -- layer=1 filter=122 channel=101
    33, 30, 29, 0, 12, 8, -36, -25, -35,
    -- layer=1 filter=122 channel=102
    30, 31, 32, 6, 16, 24, -18, -26, -16,
    -- layer=1 filter=122 channel=103
    -14, -17, 1, 3, -1, 12, -9, -3, 0,
    -- layer=1 filter=122 channel=104
    -17, 7, 0, -10, -6, -32, -2, -22, 4,
    -- layer=1 filter=122 channel=105
    1, 12, 9, 3, 15, 4, -1, -6, -7,
    -- layer=1 filter=122 channel=106
    30, 29, 35, 10, 7, 16, -17, -33, -25,
    -- layer=1 filter=122 channel=107
    -2, 1, 5, -5, -6, 1, 15, -5, -3,
    -- layer=1 filter=122 channel=108
    -34, -31, 3, -76, -103, -24, -40, -97, -50,
    -- layer=1 filter=122 channel=109
    4, 0, -8, 2, 0, -2, -8, 0, 6,
    -- layer=1 filter=122 channel=110
    -4, -2, -2, 2, 7, -2, -9, -1, 5,
    -- layer=1 filter=122 channel=111
    33, 20, 11, 25, 31, 25, 11, 11, -6,
    -- layer=1 filter=122 channel=112
    21, 7, 5, 32, -3, 24, -3, -4, -16,
    -- layer=1 filter=122 channel=113
    -7, 9, 7, 7, 10, 5, 0, 4, 1,
    -- layer=1 filter=122 channel=114
    -7, -22, -21, -31, -19, -29, -27, -27, -10,
    -- layer=1 filter=122 channel=115
    22, 24, 8, 12, 10, 15, -1, 0, 18,
    -- layer=1 filter=122 channel=116
    0, -10, -2, 4, 7, -9, 0, -3, 1,
    -- layer=1 filter=122 channel=117
    7, 10, 14, 2, 11, 29, -23, -18, -12,
    -- layer=1 filter=122 channel=118
    38, 16, 16, 28, 27, 26, 26, 4, -3,
    -- layer=1 filter=122 channel=119
    -7, -24, 10, -19, -40, -18, -11, -66, -33,
    -- layer=1 filter=122 channel=120
    17, 2, 24, -44, -36, -18, -42, -55, -34,
    -- layer=1 filter=122 channel=121
    -13, -22, 4, 20, -3, 7, 22, 11, 16,
    -- layer=1 filter=122 channel=122
    3, 6, -4, -6, -4, -5, -6, 0, 9,
    -- layer=1 filter=122 channel=123
    -17, -27, -15, -3, 1, 0, 19, 11, 10,
    -- layer=1 filter=122 channel=124
    -9, -18, -2, -6, -1, -3, -15, -11, 0,
    -- layer=1 filter=122 channel=125
    0, 3, -9, 20, 49, 40, -33, -20, -4,
    -- layer=1 filter=122 channel=126
    41, -4, 16, 13, -4, -1, -55, -53, -39,
    -- layer=1 filter=122 channel=127
    37, 18, 35, 34, 35, 37, 35, 33, 21,
    -- layer=1 filter=123 channel=0
    2, 10, 3, -4, 5, 11, -2, 6, 11,
    -- layer=1 filter=123 channel=1
    -11, 0, -8, 1, -17, 7, 10, -14, 0,
    -- layer=1 filter=123 channel=2
    19, 1, 9, 31, 12, 22, 15, 21, 4,
    -- layer=1 filter=123 channel=3
    -7, 7, 7, 1, 0, -7, -8, 3, -3,
    -- layer=1 filter=123 channel=4
    -7, -6, -10, -5, -9, 1, 0, 4, -2,
    -- layer=1 filter=123 channel=5
    2, 7, 7, -20, -10, -5, 14, -3, -2,
    -- layer=1 filter=123 channel=6
    -5, -11, 7, -33, -34, -33, -51, -39, -23,
    -- layer=1 filter=123 channel=7
    -26, -66, -60, -37, -103, -74, -39, -77, -81,
    -- layer=1 filter=123 channel=8
    4, 0, -6, 2, -6, 8, 11, 9, 10,
    -- layer=1 filter=123 channel=9
    -33, -38, -34, -31, -41, 1, 0, -6, 10,
    -- layer=1 filter=123 channel=10
    -14, -37, -43, -6, -83, -46, -29, -71, -80,
    -- layer=1 filter=123 channel=11
    -18, 1, 0, 7, -4, -10, -17, -14, -18,
    -- layer=1 filter=123 channel=12
    -32, -28, -21, -28, -33, -12, 27, 14, 15,
    -- layer=1 filter=123 channel=13
    -1, 2, 3, -8, -5, -3, 0, 7, 8,
    -- layer=1 filter=123 channel=14
    8, -29, -23, 20, -42, -22, 28, -29, -59,
    -- layer=1 filter=123 channel=15
    -5, -11, -2, -3, -27, -16, -30, -23, -33,
    -- layer=1 filter=123 channel=16
    20, 11, 5, 12, 2, 4, 8, 11, 17,
    -- layer=1 filter=123 channel=17
    -30, -16, -12, -14, -15, -14, -10, -12, 2,
    -- layer=1 filter=123 channel=18
    -6, 10, 18, 15, 2, 10, 20, 3, 6,
    -- layer=1 filter=123 channel=19
    0, 13, 46, 54, 30, 32, -12, -14, 25,
    -- layer=1 filter=123 channel=20
    -4, -11, 4, -10, -3, -1, 15, 1, 17,
    -- layer=1 filter=123 channel=21
    -3, -5, -15, 4, -6, -8, 14, 8, 4,
    -- layer=1 filter=123 channel=22
    1, -23, -10, 2, -2, -1, 32, 16, 24,
    -- layer=1 filter=123 channel=23
    -9, -71, -26, -43, -46, -45, -49, -83, -43,
    -- layer=1 filter=123 channel=24
    7, 3, 6, 3, 2, 2, 14, 21, 27,
    -- layer=1 filter=123 channel=25
    -3, -23, -12, -7, -39, -17, -7, -10, -1,
    -- layer=1 filter=123 channel=26
    -3, -24, -4, 6, -47, -21, -5, -12, 4,
    -- layer=1 filter=123 channel=27
    -44, -18, -44, -17, -27, -18, -12, -24, -8,
    -- layer=1 filter=123 channel=28
    -2, 0, -33, -9, -39, -34, 21, -29, -24,
    -- layer=1 filter=123 channel=29
    -52, -49, -52, -28, -34, -40, -32, -33, -27,
    -- layer=1 filter=123 channel=30
    12, 28, 40, 30, 11, 13, 44, 20, 14,
    -- layer=1 filter=123 channel=31
    17, -1, 17, 7, 8, 30, 22, 5, 10,
    -- layer=1 filter=123 channel=32
    -40, -66, -11, -54, -92, -35, -30, -89, -45,
    -- layer=1 filter=123 channel=33
    9, 10, 3, -22, 8, 4, -6, 0, -7,
    -- layer=1 filter=123 channel=34
    -15, -25, -20, -6, 6, -5, -35, -33, -18,
    -- layer=1 filter=123 channel=35
    11, 6, 6, -1, 3, 7, 8, 10, 6,
    -- layer=1 filter=123 channel=36
    -7, 2, 8, -9, -7, 0, -15, -15, -18,
    -- layer=1 filter=123 channel=37
    28, 12, 14, -17, -2, 0, 3, -12, -4,
    -- layer=1 filter=123 channel=38
    2, -2, 1, 13, 4, 10, 14, 14, 15,
    -- layer=1 filter=123 channel=39
    -6, 0, 10, -33, -32, -18, 1, -3, 0,
    -- layer=1 filter=123 channel=40
    18, 0, 22, -19, -14, -8, 0, -9, 6,
    -- layer=1 filter=123 channel=41
    -42, -55, 22, -68, -88, -21, -24, -103, -30,
    -- layer=1 filter=123 channel=42
    11, 8, 13, 37, 12, 28, 14, 10, 4,
    -- layer=1 filter=123 channel=43
    21, -2, 2, 2, -14, 0, 17, -3, -3,
    -- layer=1 filter=123 channel=44
    -58, -81, -41, -50, -96, -49, -37, -78, -64,
    -- layer=1 filter=123 channel=45
    -11, -9, -4, -7, -3, 9, 0, -20, -6,
    -- layer=1 filter=123 channel=46
    34, 48, 23, 66, 31, 31, 23, 11, 7,
    -- layer=1 filter=123 channel=47
    6, -67, 8, -39, -51, -38, -24, -66, -42,
    -- layer=1 filter=123 channel=48
    10, 12, 7, 0, 4, -6, 3, 9, 11,
    -- layer=1 filter=123 channel=49
    25, 6, 27, 4, 17, 20, -1, -10, 3,
    -- layer=1 filter=123 channel=50
    -7, -9, -15, 2, -7, -9, 3, 18, -4,
    -- layer=1 filter=123 channel=51
    19, 16, 10, 8, 7, -17, 18, 14, -13,
    -- layer=1 filter=123 channel=52
    0, 9, 24, 15, 15, 16, 8, 0, 11,
    -- layer=1 filter=123 channel=53
    4, 6, 0, 13, 8, 5, 20, 11, 5,
    -- layer=1 filter=123 channel=54
    16, 1, 0, 34, -16, -20, -11, -36, -11,
    -- layer=1 filter=123 channel=55
    -3, 9, 21, 3, 3, 8, -6, 2, 16,
    -- layer=1 filter=123 channel=56
    -9, 8, 1, -1, -7, 5, 5, 2, 2,
    -- layer=1 filter=123 channel=57
    -8, -17, -6, 9, -15, -1, 10, -25, -31,
    -- layer=1 filter=123 channel=58
    -18, -79, 3, -63, -66, -43, -88, -80, -83,
    -- layer=1 filter=123 channel=59
    0, -4, 0, 5, -4, -5, -6, -9, 7,
    -- layer=1 filter=123 channel=60
    10, 7, -8, -2, 3, 5, -3, -2, 13,
    -- layer=1 filter=123 channel=61
    3, -4, 5, 5, 8, 8, -5, 4, 11,
    -- layer=1 filter=123 channel=62
    14, -15, 14, 14, 4, 9, 12, -2, 21,
    -- layer=1 filter=123 channel=63
    -15, 5, -3, 13, 6, 1, 0, -14, -9,
    -- layer=1 filter=123 channel=64
    6, -9, -5, 0, -5, -3, 10, 6, -12,
    -- layer=1 filter=123 channel=65
    -2, 11, -4, -2, 8, -15, -2, 7, 7,
    -- layer=1 filter=123 channel=66
    -5, -3, 0, 7, -2, 15, -15, -10, 2,
    -- layer=1 filter=123 channel=67
    -8, -11, -3, -24, -33, -51, -62, -54, -57,
    -- layer=1 filter=123 channel=68
    -79, -65, -42, -82, -122, -60, -72, -98, -63,
    -- layer=1 filter=123 channel=69
    21, -14, 28, 4, -17, 0, 5, -13, 0,
    -- layer=1 filter=123 channel=70
    20, 24, 27, 8, -1, 17, -27, -40, -46,
    -- layer=1 filter=123 channel=71
    10, 1, 1, 18, 5, 15, 1, 13, 0,
    -- layer=1 filter=123 channel=72
    -1, 15, 34, 25, 13, 32, 23, -2, 31,
    -- layer=1 filter=123 channel=73
    -2, -11, -2, 3, -7, 3, 0, 5, 4,
    -- layer=1 filter=123 channel=74
    -30, 7, -6, -13, -13, -6, -10, -21, 0,
    -- layer=1 filter=123 channel=75
    -15, -21, -23, 19, 6, 26, 25, 12, 10,
    -- layer=1 filter=123 channel=76
    -21, -2, 0, -13, -17, -21, -9, 0, -10,
    -- layer=1 filter=123 channel=77
    -7, 10, 1, 14, 6, 10, 3, 5, 11,
    -- layer=1 filter=123 channel=78
    -29, -17, -11, -7, -14, -17, -6, -19, -15,
    -- layer=1 filter=123 channel=79
    26, -1, 14, 0, 1, 0, 8, 3, 10,
    -- layer=1 filter=123 channel=80
    -6, -10, -6, -8, -11, -4, -9, -13, -13,
    -- layer=1 filter=123 channel=81
    9, 4, 3, 4, 5, -10, -3, 14, -5,
    -- layer=1 filter=123 channel=82
    12, 9, 6, 9, 6, 7, 12, 13, 3,
    -- layer=1 filter=123 channel=83
    -7, -36, -16, 1, -20, -17, 8, -12, -1,
    -- layer=1 filter=123 channel=84
    1, 30, 23, -11, 15, 9, 26, 6, 26,
    -- layer=1 filter=123 channel=85
    4, -56, -2, -45, -17, -12, -54, -67, -42,
    -- layer=1 filter=123 channel=86
    -4, 9, 11, 4, 1, 12, -13, -12, 3,
    -- layer=1 filter=123 channel=87
    11, 13, 14, 37, 31, 28, 30, 4, 13,
    -- layer=1 filter=123 channel=88
    2, -10, -7, -16, 8, -18, 0, -9, 1,
    -- layer=1 filter=123 channel=89
    18, 10, -3, -12, 5, 5, 12, 16, 6,
    -- layer=1 filter=123 channel=90
    -68, -108, -55, -47, -102, -48, -52, -101, -65,
    -- layer=1 filter=123 channel=91
    9, 20, 9, 4, -4, 14, 21, 13, 8,
    -- layer=1 filter=123 channel=92
    -30, -53, 7, -91, -40, -33, -26, -63, -20,
    -- layer=1 filter=123 channel=93
    14, 4, 16, 5, 15, 9, 3, 24, 12,
    -- layer=1 filter=123 channel=94
    -18, -12, 0, -18, -18, -12, -7, -4, 1,
    -- layer=1 filter=123 channel=95
    1, 24, 18, 5, 5, 19, 18, 17, 26,
    -- layer=1 filter=123 channel=96
    -26, -1, -11, -15, -10, -3, -24, -17, 1,
    -- layer=1 filter=123 channel=97
    -12, 6, -4, -5, 4, 6, 7, 7, 4,
    -- layer=1 filter=123 channel=98
    22, -10, 14, 15, -7, 14, 17, 9, 2,
    -- layer=1 filter=123 channel=99
    -40, -10, -36, -8, -38, -66, 12, -74, -68,
    -- layer=1 filter=123 channel=100
    -8, 3, -9, 9, 12, 6, 1, -7, 1,
    -- layer=1 filter=123 channel=101
    21, 15, 3, 9, 11, 4, 8, 12, 8,
    -- layer=1 filter=123 channel=102
    -16, -9, -7, -22, -14, -8, -15, -4, -4,
    -- layer=1 filter=123 channel=103
    -33, -8, -25, -4, 18, -2, -4, -16, 0,
    -- layer=1 filter=123 channel=104
    10, 1, 12, -14, -2, -28, -18, -13, -35,
    -- layer=1 filter=123 channel=105
    -6, -7, 1, 8, -6, -1, -4, 0, 10,
    -- layer=1 filter=123 channel=106
    9, 5, 18, 0, -11, 1, 1, 1, 8,
    -- layer=1 filter=123 channel=107
    7, -8, 7, 0, -7, -7, 14, 0, -2,
    -- layer=1 filter=123 channel=108
    -34, -91, -33, -53, -118, -62, -46, -106, -59,
    -- layer=1 filter=123 channel=109
    9, 4, 9, -5, -8, -7, 3, -5, 3,
    -- layer=1 filter=123 channel=110
    4, 4, 3, -7, 0, 6, 5, 0, -13,
    -- layer=1 filter=123 channel=111
    10, 23, 31, 23, 21, 23, 37, 18, 25,
    -- layer=1 filter=123 channel=112
    15, 40, 39, 8, 9, 9, 6, 16, 19,
    -- layer=1 filter=123 channel=113
    4, -6, 2, 39, 19, 35, 19, 29, 25,
    -- layer=1 filter=123 channel=114
    19, 8, -7, -30, -46, -34, 1, -29, -9,
    -- layer=1 filter=123 channel=115
    -1, -12, 6, -7, -14, 8, 0, -12, 0,
    -- layer=1 filter=123 channel=116
    -2, -9, 6, -6, -3, -3, -5, -10, 2,
    -- layer=1 filter=123 channel=117
    33, 38, 36, 38, 7, 1, 59, 36, 10,
    -- layer=1 filter=123 channel=118
    1, 35, 18, 19, 14, 24, 43, 17, 17,
    -- layer=1 filter=123 channel=119
    -53, -81, -32, -85, -127, -73, -64, -115, -47,
    -- layer=1 filter=123 channel=120
    4, -8, 1, 0, 0, 0, 1, 7, -1,
    -- layer=1 filter=123 channel=121
    10, 26, 8, 56, 26, 37, 32, 31, -6,
    -- layer=1 filter=123 channel=122
    -6, -9, 8, 4, 8, 6, 8, 8, -2,
    -- layer=1 filter=123 channel=123
    13, 6, 14, 26, 28, 32, 5, 18, 12,
    -- layer=1 filter=123 channel=124
    -21, -10, -3, 0, -11, -16, -25, -18, -13,
    -- layer=1 filter=123 channel=125
    29, 1, 22, 9, -14, -9, -16, -46, -58,
    -- layer=1 filter=123 channel=126
    7, -17, 0, 27, -13, 0, 20, 24, 3,
    -- layer=1 filter=123 channel=127
    9, 53, 43, 25, 32, 24, 41, 19, 35,
    -- layer=1 filter=124 channel=0
    -8, -8, -2, -4, 2, -10, -18, -15, 1,
    -- layer=1 filter=124 channel=1
    -15, -17, -6, -4, -6, -22, -16, 2, -6,
    -- layer=1 filter=124 channel=2
    -2, -1, -10, -3, 0, -7, 5, 7, 7,
    -- layer=1 filter=124 channel=3
    0, 3, -8, -6, -8, 1, -6, 5, -3,
    -- layer=1 filter=124 channel=4
    -4, 6, -1, 3, 5, -6, -3, -8, -6,
    -- layer=1 filter=124 channel=5
    -2, -13, -13, -2, -19, -18, -2, 1, -7,
    -- layer=1 filter=124 channel=6
    4, -5, -12, 0, -13, -6, -9, 2, -6,
    -- layer=1 filter=124 channel=7
    -12, 10, -12, -5, -3, 3, -18, -18, 10,
    -- layer=1 filter=124 channel=8
    -15, -13, -23, 0, -6, -19, 1, 0, -8,
    -- layer=1 filter=124 channel=9
    2, 5, -6, 0, -3, 0, -13, -5, 2,
    -- layer=1 filter=124 channel=10
    -9, 5, 4, -7, -3, -7, -2, -7, 2,
    -- layer=1 filter=124 channel=11
    -5, -2, 2, -7, -14, -14, -10, -12, -4,
    -- layer=1 filter=124 channel=12
    4, -1, -9, -9, 16, 9, 1, -6, -7,
    -- layer=1 filter=124 channel=13
    -8, -4, -2, -10, -11, -13, -3, -8, -12,
    -- layer=1 filter=124 channel=14
    1, 2, 9, 17, -4, 1, 0, 1, 8,
    -- layer=1 filter=124 channel=15
    -13, -22, 0, -12, -16, -3, -4, -11, -3,
    -- layer=1 filter=124 channel=16
    -18, -15, -20, -5, -2, -12, 0, -4, -14,
    -- layer=1 filter=124 channel=17
    -14, -11, -4, -5, -5, -2, -14, -9, -2,
    -- layer=1 filter=124 channel=18
    -12, 0, -19, -8, 0, 5, -1, -9, -2,
    -- layer=1 filter=124 channel=19
    -8, 0, -9, 10, -6, 2, 0, -10, -4,
    -- layer=1 filter=124 channel=20
    -7, -7, -14, -5, -7, 2, 0, -13, -4,
    -- layer=1 filter=124 channel=21
    -11, -2, -11, 1, 2, 0, -7, 6, -7,
    -- layer=1 filter=124 channel=22
    -7, -9, -12, -12, 0, -11, -16, -5, -13,
    -- layer=1 filter=124 channel=23
    -2, 10, 0, 0, -12, -15, -9, -8, 0,
    -- layer=1 filter=124 channel=24
    -12, -12, -8, 0, -3, -13, 6, -12, -1,
    -- layer=1 filter=124 channel=25
    -9, 3, -13, 0, -3, -11, -16, -10, -7,
    -- layer=1 filter=124 channel=26
    -3, -13, -2, 7, -18, -16, 1, -3, -21,
    -- layer=1 filter=124 channel=27
    -9, -2, -4, -11, -6, 6, -16, -8, -2,
    -- layer=1 filter=124 channel=28
    -14, 8, 3, -4, -3, -8, -9, -14, -12,
    -- layer=1 filter=124 channel=29
    -1, -6, 10, 0, 16, 19, -5, 13, 2,
    -- layer=1 filter=124 channel=30
    -4, 5, -7, -2, 2, 0, -4, -5, -2,
    -- layer=1 filter=124 channel=31
    -11, 0, -11, -5, -1, -7, 3, 1, 3,
    -- layer=1 filter=124 channel=32
    0, -8, -12, -4, -10, -4, -4, -5, -17,
    -- layer=1 filter=124 channel=33
    -7, -2, -7, -6, -6, 1, -9, -7, 2,
    -- layer=1 filter=124 channel=34
    -9, -14, 3, 5, -5, -11, -7, -10, -2,
    -- layer=1 filter=124 channel=35
    6, -6, -10, -6, -3, 0, -8, -10, 4,
    -- layer=1 filter=124 channel=36
    -4, -11, 0, -14, -15, -13, -17, -4, -9,
    -- layer=1 filter=124 channel=37
    -4, 0, -5, -18, -1, -10, 2, -9, -14,
    -- layer=1 filter=124 channel=38
    8, -9, 5, 9, 3, -5, 9, -8, -4,
    -- layer=1 filter=124 channel=39
    -17, -14, -4, -21, -8, -22, -6, -18, -11,
    -- layer=1 filter=124 channel=40
    -10, -5, 0, 7, -2, 2, 8, 4, 10,
    -- layer=1 filter=124 channel=41
    3, -13, 2, -9, -7, -11, -8, -3, 3,
    -- layer=1 filter=124 channel=42
    -6, 4, -3, -2, 6, 6, -2, 3, 1,
    -- layer=1 filter=124 channel=43
    -9, -13, -13, -5, -8, -7, -17, 0, 2,
    -- layer=1 filter=124 channel=44
    -14, -10, -23, -13, -13, -8, -8, -11, -8,
    -- layer=1 filter=124 channel=45
    -4, -5, -6, 8, -2, -2, -7, -10, -15,
    -- layer=1 filter=124 channel=46
    1, 6, 1, -8, 8, -14, -7, 3, -11,
    -- layer=1 filter=124 channel=47
    -5, -8, -9, -8, 1, 1, -7, -11, 1,
    -- layer=1 filter=124 channel=48
    -11, -4, -7, -14, 5, -11, -8, -14, -12,
    -- layer=1 filter=124 channel=49
    2, 0, -5, -11, 5, -8, 0, -5, -8,
    -- layer=1 filter=124 channel=50
    2, -3, 10, -4, 1, 6, 0, -6, 3,
    -- layer=1 filter=124 channel=51
    -13, 2, -14, -2, 1, -1, -10, 1, -9,
    -- layer=1 filter=124 channel=52
    -10, -1, 0, -7, 9, 2, -7, 2, -8,
    -- layer=1 filter=124 channel=53
    -1, -9, -11, -6, -6, 8, 4, 7, -4,
    -- layer=1 filter=124 channel=54
    -3, -1, -7, -19, -8, 0, -15, -15, 8,
    -- layer=1 filter=124 channel=55
    0, -10, -15, -16, 0, -10, -8, -17, -14,
    -- layer=1 filter=124 channel=56
    -8, -3, -1, 0, 6, 8, -7, -9, 8,
    -- layer=1 filter=124 channel=57
    -17, -10, -3, -6, -17, -5, -12, -22, -3,
    -- layer=1 filter=124 channel=58
    -11, 11, -13, -12, 0, -10, 3, -8, 3,
    -- layer=1 filter=124 channel=59
    5, -9, 2, 8, 9, -9, -4, 0, 5,
    -- layer=1 filter=124 channel=60
    3, 6, -5, 8, 4, 3, -7, 2, -4,
    -- layer=1 filter=124 channel=61
    -1, 5, 8, -8, -8, 8, -8, -5, 5,
    -- layer=1 filter=124 channel=62
    -6, -8, -16, -8, -1, -19, -6, -3, -16,
    -- layer=1 filter=124 channel=63
    -5, -3, -3, -10, -7, 0, -17, 0, 2,
    -- layer=1 filter=124 channel=64
    0, -7, -15, -12, -9, -14, -4, -15, -1,
    -- layer=1 filter=124 channel=65
    -2, 3, 2, -15, 2, 5, -4, -5, 0,
    -- layer=1 filter=124 channel=66
    -15, -1, -5, -3, -13, -5, -4, -10, -13,
    -- layer=1 filter=124 channel=67
    0, 1, 0, 3, -14, -7, 8, -2, -2,
    -- layer=1 filter=124 channel=68
    -5, -7, -17, -7, -5, -9, 1, 0, -21,
    -- layer=1 filter=124 channel=69
    -13, -12, -15, 5, 2, -16, 0, -9, -7,
    -- layer=1 filter=124 channel=70
    -10, -3, -6, -3, -3, 4, 3, -3, 2,
    -- layer=1 filter=124 channel=71
    -8, 4, -6, -17, 3, -8, -3, -12, 4,
    -- layer=1 filter=124 channel=72
    -6, 4, -9, 4, -7, 1, -16, -8, 1,
    -- layer=1 filter=124 channel=73
    1, -2, -6, 0, 9, -9, -11, -9, -9,
    -- layer=1 filter=124 channel=74
    0, 1, 0, 6, 2, -2, -2, 0, -9,
    -- layer=1 filter=124 channel=75
    3, -3, 0, 3, -4, 6, -5, 0, 0,
    -- layer=1 filter=124 channel=76
    4, 0, 0, 3, -10, -14, -2, -14, -10,
    -- layer=1 filter=124 channel=77
    0, -9, 3, -11, -7, -4, -2, -5, -14,
    -- layer=1 filter=124 channel=78
    -17, -7, -11, -17, -1, -10, 0, -8, -1,
    -- layer=1 filter=124 channel=79
    -12, -5, -19, -6, -1, -21, -9, 1, -8,
    -- layer=1 filter=124 channel=80
    7, -9, 6, 0, 3, 0, -3, -14, -9,
    -- layer=1 filter=124 channel=81
    -3, -8, -16, -3, -4, -15, -1, -10, -13,
    -- layer=1 filter=124 channel=82
    -12, -12, 1, -13, 2, -4, 4, -5, -12,
    -- layer=1 filter=124 channel=83
    -20, -2, -26, -7, -5, 2, -16, -6, -18,
    -- layer=1 filter=124 channel=84
    0, -11, -13, 2, 6, -1, -10, 0, 3,
    -- layer=1 filter=124 channel=85
    -9, 4, -10, 1, -5, -4, -14, -10, 8,
    -- layer=1 filter=124 channel=86
    -11, -7, -17, -2, -19, -4, -18, -11, -15,
    -- layer=1 filter=124 channel=87
    7, 0, -1, 8, 0, -4, -11, 7, -15,
    -- layer=1 filter=124 channel=88
    -2, -4, 0, 7, -4, 0, -2, 4, -4,
    -- layer=1 filter=124 channel=89
    -2, -5, -2, -11, 3, -8, -3, -8, -9,
    -- layer=1 filter=124 channel=90
    0, -18, -26, -9, -18, -22, -7, -2, -13,
    -- layer=1 filter=124 channel=91
    -1, 0, 3, 0, -11, -10, -11, 0, -6,
    -- layer=1 filter=124 channel=92
    1, -18, -4, 3, -15, -3, -5, -16, 1,
    -- layer=1 filter=124 channel=93
    -11, -5, -10, -15, -12, -11, -5, -1, 0,
    -- layer=1 filter=124 channel=94
    -12, -9, 0, -17, 0, -15, -10, -14, -14,
    -- layer=1 filter=124 channel=95
    -6, -7, -9, -10, -7, 0, 4, 9, -9,
    -- layer=1 filter=124 channel=96
    -5, 6, -7, -11, -6, -7, -9, 0, -8,
    -- layer=1 filter=124 channel=97
    -10, -15, -12, -13, -3, -2, -4, -18, -18,
    -- layer=1 filter=124 channel=98
    2, 0, -18, -12, -1, 0, -15, 8, -1,
    -- layer=1 filter=124 channel=99
    -6, 2, 8, -19, -2, -10, -13, -15, 0,
    -- layer=1 filter=124 channel=100
    -11, -9, -19, -12, -2, -6, -1, -6, -7,
    -- layer=1 filter=124 channel=101
    -5, 1, -8, 6, -5, -2, 5, -7, -1,
    -- layer=1 filter=124 channel=102
    -14, -1, 8, -7, -3, -1, 0, 0, 1,
    -- layer=1 filter=124 channel=103
    -17, -9, -10, 3, -4, -12, -11, -9, -3,
    -- layer=1 filter=124 channel=104
    -15, -8, 6, -4, -12, -6, 1, -1, -2,
    -- layer=1 filter=124 channel=105
    -16, 1, -2, -21, -9, -14, -11, -3, -10,
    -- layer=1 filter=124 channel=106
    2, -6, -14, 6, 0, 0, 5, -14, 0,
    -- layer=1 filter=124 channel=107
    4, 1, 3, 2, 4, -3, 6, -10, 6,
    -- layer=1 filter=124 channel=108
    3, -10, -9, -10, -23, -10, -8, -16, -25,
    -- layer=1 filter=124 channel=109
    0, -9, -8, 0, 4, 8, -3, 9, 7,
    -- layer=1 filter=124 channel=110
    -3, -4, -4, 0, 5, 8, -7, 6, -5,
    -- layer=1 filter=124 channel=111
    -7, 1, -14, -10, 0, -6, -5, 4, -8,
    -- layer=1 filter=124 channel=112
    4, -8, -15, 1, -3, -4, 0, -7, -10,
    -- layer=1 filter=124 channel=113
    -17, -19, -14, -12, -11, -11, -5, -9, -5,
    -- layer=1 filter=124 channel=114
    -12, -2, -15, 1, -15, -20, -12, -12, 0,
    -- layer=1 filter=124 channel=115
    -19, 2, -8, -5, -9, 1, -8, -23, 0,
    -- layer=1 filter=124 channel=116
    -2, -1, 7, -3, -8, -1, -8, -7, -10,
    -- layer=1 filter=124 channel=117
    9, 6, -8, -9, -5, 1, -1, -8, -11,
    -- layer=1 filter=124 channel=118
    3, -5, 0, 2, -9, -9, -10, -15, -4,
    -- layer=1 filter=124 channel=119
    -2, -16, -23, 1, -14, -3, -8, -3, -15,
    -- layer=1 filter=124 channel=120
    -1, -5, -2, -7, 0, -7, -9, -12, 6,
    -- layer=1 filter=124 channel=121
    -8, -8, -7, -11, -9, -5, -11, 0, 1,
    -- layer=1 filter=124 channel=122
    8, 0, 7, -3, 5, -2, 3, 8, 6,
    -- layer=1 filter=124 channel=123
    -4, -4, -12, -1, -8, -8, 3, -1, -9,
    -- layer=1 filter=124 channel=124
    3, -10, -8, 8, -3, -10, 5, 2, 0,
    -- layer=1 filter=124 channel=125
    -8, -5, -11, -11, -10, 2, 0, -18, 5,
    -- layer=1 filter=124 channel=126
    -2, -1, -8, -5, -5, 0, -6, 10, -4,
    -- layer=1 filter=124 channel=127
    -9, -4, -4, 8, -2, 0, -2, 2, 1,
    -- layer=1 filter=125 channel=0
    -2, -2, -13, 3, -7, 1, 0, -11, -3,
    -- layer=1 filter=125 channel=1
    -1, -2, -5, -14, -11, -18, -10, -4, -7,
    -- layer=1 filter=125 channel=2
    -17, -6, -11, -7, -6, -8, -10, -11, -10,
    -- layer=1 filter=125 channel=3
    9, -3, -8, 3, 2, 4, -1, -6, 1,
    -- layer=1 filter=125 channel=4
    0, -7, 6, 9, -2, -5, -5, 4, 2,
    -- layer=1 filter=125 channel=5
    -3, 8, 7, -15, -20, -9, -20, -7, -2,
    -- layer=1 filter=125 channel=6
    -6, -20, -17, -22, -2, -4, -4, -16, -18,
    -- layer=1 filter=125 channel=7
    -6, -7, 6, -3, -9, -1, 4, -20, -9,
    -- layer=1 filter=125 channel=8
    3, 13, -7, 4, -5, -21, -4, -8, -17,
    -- layer=1 filter=125 channel=9
    -16, -4, -3, -6, 7, 0, 0, 6, 5,
    -- layer=1 filter=125 channel=10
    -2, 4, -11, -13, -8, -16, -5, -20, 0,
    -- layer=1 filter=125 channel=11
    2, -8, -3, 5, -5, 9, 0, 2, 8,
    -- layer=1 filter=125 channel=12
    -1, 0, -2, 11, -8, 1, 1, 0, -15,
    -- layer=1 filter=125 channel=13
    -12, -7, -12, -8, -8, -18, -7, -15, -1,
    -- layer=1 filter=125 channel=14
    0, -9, -2, -4, -6, -5, -16, -11, 2,
    -- layer=1 filter=125 channel=15
    -11, -6, -11, 0, -18, -2, 0, -11, -13,
    -- layer=1 filter=125 channel=16
    -7, 11, 3, 2, -6, -2, -17, -12, -12,
    -- layer=1 filter=125 channel=17
    -5, -6, -2, -6, 0, -8, -3, -7, -7,
    -- layer=1 filter=125 channel=18
    -8, -13, -18, -4, -6, 4, -15, -15, -12,
    -- layer=1 filter=125 channel=19
    -12, 4, -10, -11, -13, -5, -14, -1, -5,
    -- layer=1 filter=125 channel=20
    -5, -2, -10, -6, -12, -6, -1, -9, -1,
    -- layer=1 filter=125 channel=21
    0, -15, 2, 0, -7, -16, -14, -3, -16,
    -- layer=1 filter=125 channel=22
    -9, 6, 4, 6, -15, -13, 0, 1, -18,
    -- layer=1 filter=125 channel=23
    0, 6, 5, -8, 1, -13, -2, 2, 4,
    -- layer=1 filter=125 channel=24
    -11, 5, -14, -7, -18, 1, -15, 3, 2,
    -- layer=1 filter=125 channel=25
    4, 3, 6, 0, 0, -11, -7, -4, -10,
    -- layer=1 filter=125 channel=26
    -5, 7, -8, 0, -7, -9, -15, 2, -3,
    -- layer=1 filter=125 channel=27
    -10, -17, -11, -11, -23, -9, -17, -11, -13,
    -- layer=1 filter=125 channel=28
    4, -9, 3, -1, -12, 0, -4, -21, 5,
    -- layer=1 filter=125 channel=29
    -3, 0, -14, 4, -4, -11, -4, -7, 1,
    -- layer=1 filter=125 channel=30
    -18, -10, -14, -17, -5, 3, -10, -8, -15,
    -- layer=1 filter=125 channel=31
    -13, -15, 2, 0, -3, 6, -16, -7, -12,
    -- layer=1 filter=125 channel=32
    -4, 2, -4, -3, -2, -11, 3, 0, -10,
    -- layer=1 filter=125 channel=33
    -2, 0, -8, 3, -6, -8, -6, 0, -5,
    -- layer=1 filter=125 channel=34
    -16, 0, -4, -14, 0, 1, 2, -15, 0,
    -- layer=1 filter=125 channel=35
    -11, -9, -7, 9, -18, -3, -9, -1, -6,
    -- layer=1 filter=125 channel=36
    4, 2, -14, -9, 1, -7, -8, 7, 8,
    -- layer=1 filter=125 channel=37
    -1, 9, 7, 1, -18, -18, -16, 2, 1,
    -- layer=1 filter=125 channel=38
    -15, -17, -9, 0, -17, -7, -9, -18, -10,
    -- layer=1 filter=125 channel=39
    6, -4, -2, -3, -8, 1, -9, -2, 4,
    -- layer=1 filter=125 channel=40
    -1, -5, -4, -8, 3, -8, -6, -11, -5,
    -- layer=1 filter=125 channel=41
    -3, 0, -1, 5, 0, 18, 0, 9, 0,
    -- layer=1 filter=125 channel=42
    1, -8, 3, -7, -15, -10, -12, 0, -10,
    -- layer=1 filter=125 channel=43
    -2, 3, 2, -6, -6, -6, -10, 3, -13,
    -- layer=1 filter=125 channel=44
    -1, 3, 0, -9, 5, 1, -1, -8, -6,
    -- layer=1 filter=125 channel=45
    -10, 4, 0, -14, -3, -8, 2, -10, -5,
    -- layer=1 filter=125 channel=46
    5, -6, -11, -13, -22, -8, -8, -9, 0,
    -- layer=1 filter=125 channel=47
    0, -1, -6, 2, -6, 10, -4, 5, -1,
    -- layer=1 filter=125 channel=48
    -12, 0, -18, 1, 0, -6, -4, -13, -8,
    -- layer=1 filter=125 channel=49
    -16, -3, -9, 0, -3, -15, -5, -11, -1,
    -- layer=1 filter=125 channel=50
    -8, 3, 3, 0, 4, -5, 7, 0, -5,
    -- layer=1 filter=125 channel=51
    0, 1, -10, -9, -14, -11, -4, -14, -13,
    -- layer=1 filter=125 channel=52
    4, -3, -10, 7, -5, 9, 1, -1, 7,
    -- layer=1 filter=125 channel=53
    0, 7, 5, 0, 4, 1, -10, -1, -8,
    -- layer=1 filter=125 channel=54
    0, 9, -8, 1, 1, -9, 1, -2, 3,
    -- layer=1 filter=125 channel=55
    1, 6, -4, -15, -8, 5, -6, -3, 4,
    -- layer=1 filter=125 channel=56
    -5, -9, 2, 0, -9, 2, 0, -11, 4,
    -- layer=1 filter=125 channel=57
    -5, 0, -3, -5, -2, -3, -13, -14, -11,
    -- layer=1 filter=125 channel=58
    -2, 4, -16, -6, -10, -8, -11, -11, 0,
    -- layer=1 filter=125 channel=59
    0, -9, 8, 8, -6, -9, -13, 0, 3,
    -- layer=1 filter=125 channel=60
    -4, 7, -3, 0, 6, 3, -5, 5, -1,
    -- layer=1 filter=125 channel=61
    5, -5, 6, 8, -4, -2, -9, -9, 4,
    -- layer=1 filter=125 channel=62
    -7, -1, -4, -12, -14, -2, -17, 0, -3,
    -- layer=1 filter=125 channel=63
    1, -3, 1, -6, 3, -5, 1, 3, -1,
    -- layer=1 filter=125 channel=64
    -8, -14, -10, -11, -4, -4, -1, 0, -14,
    -- layer=1 filter=125 channel=65
    -1, -11, -10, -2, -1, -12, -16, 0, -5,
    -- layer=1 filter=125 channel=66
    -14, -12, 4, 1, -6, 5, -8, -7, -6,
    -- layer=1 filter=125 channel=67
    6, 4, 3, 4, -3, -12, -3, -7, 0,
    -- layer=1 filter=125 channel=68
    -7, -12, -7, 1, 5, 2, 3, -2, -7,
    -- layer=1 filter=125 channel=69
    -10, -3, -1, -6, -8, -6, -11, -7, -7,
    -- layer=1 filter=125 channel=70
    0, -8, 6, -10, 3, -4, 2, -14, -13,
    -- layer=1 filter=125 channel=71
    0, -13, -9, -1, -12, -12, -6, -3, -15,
    -- layer=1 filter=125 channel=72
    -23, -17, -23, 4, -5, -5, -3, -2, -4,
    -- layer=1 filter=125 channel=73
    -7, 4, 5, 8, -12, 4, 1, -5, 9,
    -- layer=1 filter=125 channel=74
    0, -6, -12, -15, 1, 8, -8, -11, -11,
    -- layer=1 filter=125 channel=75
    -15, -5, -24, -9, 5, -11, -5, -21, -16,
    -- layer=1 filter=125 channel=76
    -10, -7, -13, -11, -12, 0, 0, -7, -13,
    -- layer=1 filter=125 channel=77
    -4, -12, -3, -10, -11, -1, 2, -18, -17,
    -- layer=1 filter=125 channel=78
    -10, -8, 2, 0, -18, -15, -11, -12, 2,
    -- layer=1 filter=125 channel=79
    -6, 10, -1, 0, 4, -13, -15, 1, -7,
    -- layer=1 filter=125 channel=80
    -8, -5, -2, 5, -13, -6, -12, -5, 0,
    -- layer=1 filter=125 channel=81
    -6, 6, -9, -11, -10, -15, -7, 4, -3,
    -- layer=1 filter=125 channel=82
    -10, -19, 1, -10, -4, -16, -1, -11, -11,
    -- layer=1 filter=125 channel=83
    8, 4, 6, -2, -9, -6, -10, 0, -11,
    -- layer=1 filter=125 channel=84
    -14, -18, -12, -15, -7, 5, -7, -11, -6,
    -- layer=1 filter=125 channel=85
    5, -3, -12, 2, -6, 11, 9, -2, -9,
    -- layer=1 filter=125 channel=86
    -2, -12, -2, 1, 3, -5, -2, 2, 4,
    -- layer=1 filter=125 channel=87
    -4, -10, 1, 10, -7, 8, -12, -3, 0,
    -- layer=1 filter=125 channel=88
    -8, -18, 0, -4, -10, 1, -9, -15, -17,
    -- layer=1 filter=125 channel=89
    -1, -7, -12, -2, -13, -15, 1, -8, -2,
    -- layer=1 filter=125 channel=90
    -7, 2, 7, -9, 0, 7, -5, -2, 0,
    -- layer=1 filter=125 channel=91
    -15, -8, 0, -16, -7, -5, 0, -9, -3,
    -- layer=1 filter=125 channel=92
    -1, -5, -4, 9, 8, 2, -7, 8, -2,
    -- layer=1 filter=125 channel=93
    0, -9, 0, -11, -9, -17, 2, -2, -5,
    -- layer=1 filter=125 channel=94
    -1, -7, -9, 0, -12, -9, -3, -14, -3,
    -- layer=1 filter=125 channel=95
    -22, -13, -14, -11, -12, 0, -5, 0, -16,
    -- layer=1 filter=125 channel=96
    -4, 8, -6, 2, 7, 16, -4, -6, 19,
    -- layer=1 filter=125 channel=97
    -9, -1, -10, -10, 3, -10, -13, 4, -13,
    -- layer=1 filter=125 channel=98
    -5, 9, 6, 5, -13, -20, -8, -20, -14,
    -- layer=1 filter=125 channel=99
    -17, -14, -5, -10, -13, -3, -8, -12, -9,
    -- layer=1 filter=125 channel=100
    -1, -6, -11, 7, -8, 1, -1, 7, -3,
    -- layer=1 filter=125 channel=101
    -14, -8, -17, -4, 0, -9, -6, -10, -18,
    -- layer=1 filter=125 channel=102
    -12, -19, -16, -12, -4, -12, -5, -11, -12,
    -- layer=1 filter=125 channel=103
    -7, -5, -5, -2, -6, -5, 0, 2, 3,
    -- layer=1 filter=125 channel=104
    -3, -5, 0, -9, 10, -4, -14, 9, -13,
    -- layer=1 filter=125 channel=105
    -2, -15, -3, -1, -13, -11, 2, -12, -6,
    -- layer=1 filter=125 channel=106
    -2, 0, -9, -14, -6, -1, -13, -13, -9,
    -- layer=1 filter=125 channel=107
    -9, 6, 9, 1, -6, -1, 4, -5, 7,
    -- layer=1 filter=125 channel=108
    -3, 0, 5, 0, 0, -2, -6, -14, 1,
    -- layer=1 filter=125 channel=109
    -7, 6, 0, -7, 1, 5, -10, 2, 4,
    -- layer=1 filter=125 channel=110
    -14, -6, -5, 2, 0, -2, 7, -17, -15,
    -- layer=1 filter=125 channel=111
    -22, -23, -17, -2, -10, -11, 4, -8, -11,
    -- layer=1 filter=125 channel=112
    -15, -19, -11, -4, 2, 3, -14, -17, -12,
    -- layer=1 filter=125 channel=113
    -11, 0, -10, -12, -1, -3, 6, -8, -14,
    -- layer=1 filter=125 channel=114
    -9, -2, -10, -16, -8, -3, -13, -9, -15,
    -- layer=1 filter=125 channel=115
    4, 6, -4, 2, -1, -2, -12, 0, 4,
    -- layer=1 filter=125 channel=116
    10, 4, 9, -1, 9, -9, 2, -1, -3,
    -- layer=1 filter=125 channel=117
    -12, -14, -8, -1, -4, -9, -7, -5, 0,
    -- layer=1 filter=125 channel=118
    -9, -4, -4, -3, 0, 6, -13, -13, 2,
    -- layer=1 filter=125 channel=119
    5, -2, -12, -13, 6, 6, 1, -12, 6,
    -- layer=1 filter=125 channel=120
    -4, -14, -3, 2, -16, -10, -13, -13, -4,
    -- layer=1 filter=125 channel=121
    -18, -12, -18, -10, -19, -2, -14, 6, 4,
    -- layer=1 filter=125 channel=122
    0, 0, -7, 4, 4, 7, 5, 7, 2,
    -- layer=1 filter=125 channel=123
    -24, -11, -4, -1, -10, -15, -3, 3, 4,
    -- layer=1 filter=125 channel=124
    -10, -5, -4, -1, 0, -8, 4, -2, -6,
    -- layer=1 filter=125 channel=125
    -5, -4, -13, -13, 3, 1, -15, -9, -15,
    -- layer=1 filter=125 channel=126
    12, 7, 0, -3, 6, -3, 8, -6, -11,
    -- layer=1 filter=125 channel=127
    -6, -12, -13, -3, -11, 8, -10, -15, -7,
    -- layer=1 filter=126 channel=0
    -5, 2, -10, 3, 3, -7, -1, -3, -7,
    -- layer=1 filter=126 channel=1
    -3, -3, 0, 0, -5, 2, 4, -7, 1,
    -- layer=1 filter=126 channel=2
    8, -3, 5, -6, -5, -10, -11, -11, -13,
    -- layer=1 filter=126 channel=3
    3, -6, 5, -8, -11, -8, -9, 8, 0,
    -- layer=1 filter=126 channel=4
    4, -5, 2, -9, 1, -8, 2, -5, -8,
    -- layer=1 filter=126 channel=5
    6, 10, -5, 0, 0, -3, -1, 10, -11,
    -- layer=1 filter=126 channel=6
    5, 7, 1, 4, 6, -10, -2, -9, 3,
    -- layer=1 filter=126 channel=7
    3, 4, -12, -2, -7, -12, 7, 6, -9,
    -- layer=1 filter=126 channel=8
    -4, 4, 7, -12, 4, -8, -8, 0, 5,
    -- layer=1 filter=126 channel=9
    7, -9, 1, 3, -3, -7, 5, -2, 5,
    -- layer=1 filter=126 channel=10
    9, -7, -6, 1, -7, -5, 8, -7, -12,
    -- layer=1 filter=126 channel=11
    6, -1, 7, 2, -9, -9, -11, 7, 0,
    -- layer=1 filter=126 channel=12
    -6, -4, 8, 4, -4, -6, -3, -10, 0,
    -- layer=1 filter=126 channel=13
    -9, 8, 6, 2, 3, 6, -12, -4, -1,
    -- layer=1 filter=126 channel=14
    1, 0, 5, -8, -8, -10, -3, -9, 0,
    -- layer=1 filter=126 channel=15
    -3, 7, -7, 1, 0, 0, 2, 9, -10,
    -- layer=1 filter=126 channel=16
    -1, -5, 10, -2, 5, -9, 6, 7, 4,
    -- layer=1 filter=126 channel=17
    0, -9, -6, 0, -9, -7, -9, -3, 3,
    -- layer=1 filter=126 channel=18
    -3, -9, 2, -2, 4, -10, 4, 5, 7,
    -- layer=1 filter=126 channel=19
    -2, 4, 0, 1, -11, 1, -7, 3, -6,
    -- layer=1 filter=126 channel=20
    -2, 2, -7, 4, 4, 9, -9, -8, 7,
    -- layer=1 filter=126 channel=21
    4, 6, -9, -9, 2, 4, -12, -7, 8,
    -- layer=1 filter=126 channel=22
    -5, 0, -3, -8, -5, -1, -7, -3, -4,
    -- layer=1 filter=126 channel=23
    6, 3, 5, -5, -11, 5, 6, 9, -10,
    -- layer=1 filter=126 channel=24
    -5, -1, 3, -3, -9, 2, 3, -9, 4,
    -- layer=1 filter=126 channel=25
    -7, 0, -10, 2, -13, -9, 8, 5, -4,
    -- layer=1 filter=126 channel=26
    4, 6, 1, -8, -10, 0, -8, -11, 7,
    -- layer=1 filter=126 channel=27
    4, 5, 6, 2, 10, -6, 1, 9, 1,
    -- layer=1 filter=126 channel=28
    -10, -11, -7, -5, -2, -11, -6, -8, 3,
    -- layer=1 filter=126 channel=29
    0, 0, 4, -2, 5, 9, -6, -4, -9,
    -- layer=1 filter=126 channel=30
    -10, 9, 0, 7, 0, -6, 3, -8, -4,
    -- layer=1 filter=126 channel=31
    -3, -12, -6, 0, -1, 2, 6, -4, -4,
    -- layer=1 filter=126 channel=32
    1, 0, 3, -8, 5, 5, 0, -3, -10,
    -- layer=1 filter=126 channel=33
    0, 2, -6, -4, 0, 6, 1, -4, 5,
    -- layer=1 filter=126 channel=34
    4, 3, -7, -10, -3, 1, 3, 4, 0,
    -- layer=1 filter=126 channel=35
    1, 0, -5, -7, -2, -4, -3, -1, 9,
    -- layer=1 filter=126 channel=36
    10, 11, -3, 9, 6, 8, -2, 2, 2,
    -- layer=1 filter=126 channel=37
    -7, 3, 5, -6, 1, -5, -8, -4, -11,
    -- layer=1 filter=126 channel=38
    1, 4, -7, 0, -2, -1, -2, -3, -10,
    -- layer=1 filter=126 channel=39
    9, -5, 10, -8, -8, 10, -3, 4, 2,
    -- layer=1 filter=126 channel=40
    -10, -4, 3, 5, 4, 4, -3, -4, 7,
    -- layer=1 filter=126 channel=41
    -6, -3, 0, -9, -2, -3, -7, 8, -3,
    -- layer=1 filter=126 channel=42
    -8, 8, 2, -1, -4, -1, 9, -2, -1,
    -- layer=1 filter=126 channel=43
    -4, 5, 5, -7, 6, -1, 10, -3, -1,
    -- layer=1 filter=126 channel=44
    -4, -10, -9, -11, -9, -3, -5, 0, 9,
    -- layer=1 filter=126 channel=45
    5, 7, 0, -3, -4, -6, 9, -1, -8,
    -- layer=1 filter=126 channel=46
    1, 5, -9, -8, 6, 7, 7, 3, -7,
    -- layer=1 filter=126 channel=47
    0, -2, 7, 2, -1, -9, 4, -8, -10,
    -- layer=1 filter=126 channel=48
    -4, -10, -6, -5, 0, 0, -3, -2, 5,
    -- layer=1 filter=126 channel=49
    -4, -6, -12, -10, 5, -7, 5, 3, 4,
    -- layer=1 filter=126 channel=50
    2, 5, -4, 7, -9, -2, 0, 7, 0,
    -- layer=1 filter=126 channel=51
    2, 0, -11, 9, 0, 8, 7, -6, -3,
    -- layer=1 filter=126 channel=52
    10, 4, -6, 1, -4, -8, -8, 6, 8,
    -- layer=1 filter=126 channel=53
    -6, -6, 8, 1, -7, -3, 1, -9, 8,
    -- layer=1 filter=126 channel=54
    2, -6, 5, -14, -1, -6, -3, 0, -5,
    -- layer=1 filter=126 channel=55
    4, 0, 0, -8, 3, 9, 8, -7, -10,
    -- layer=1 filter=126 channel=56
    2, -5, 6, 3, 0, -2, -6, -7, -3,
    -- layer=1 filter=126 channel=57
    7, -8, -9, 9, 8, -1, -2, -9, -1,
    -- layer=1 filter=126 channel=58
    2, 0, -2, 4, -2, 5, -7, -6, -6,
    -- layer=1 filter=126 channel=59
    2, -9, 0, -8, -8, -1, 3, 3, -7,
    -- layer=1 filter=126 channel=60
    3, -3, 0, 7, -8, 6, 2, -1, 0,
    -- layer=1 filter=126 channel=61
    0, 2, 6, 0, -3, 7, -4, -7, -4,
    -- layer=1 filter=126 channel=62
    8, 2, 0, -2, 6, -5, -5, -1, -2,
    -- layer=1 filter=126 channel=63
    -3, -6, 7, -7, -4, 3, -11, 3, 9,
    -- layer=1 filter=126 channel=64
    5, 3, -2, -10, 8, -9, -8, -10, 7,
    -- layer=1 filter=126 channel=65
    -5, -1, -1, 1, 1, -7, -6, -6, 8,
    -- layer=1 filter=126 channel=66
    8, -7, -5, -7, -6, -3, 4, 0, -8,
    -- layer=1 filter=126 channel=67
    4, -1, 5, -4, -5, 10, -1, 0, 0,
    -- layer=1 filter=126 channel=68
    8, -1, -9, -1, -8, -6, -7, -3, -5,
    -- layer=1 filter=126 channel=69
    4, -11, -8, -9, -5, -6, -5, 2, 5,
    -- layer=1 filter=126 channel=70
    -8, 8, 3, -2, 4, -10, 0, 2, -2,
    -- layer=1 filter=126 channel=71
    -3, 4, -9, 2, 0, -11, -9, 2, -8,
    -- layer=1 filter=126 channel=72
    4, 4, -6, -3, 7, 3, -10, -9, -6,
    -- layer=1 filter=126 channel=73
    0, -11, 0, -3, -5, 0, -8, 0, 1,
    -- layer=1 filter=126 channel=74
    10, -5, 0, 7, 4, 0, 7, -3, 6,
    -- layer=1 filter=126 channel=75
    7, -9, 3, 0, -9, 7, -2, -8, 1,
    -- layer=1 filter=126 channel=76
    -10, 6, 3, -5, -8, -10, -10, -1, -6,
    -- layer=1 filter=126 channel=77
    7, 0, 0, -3, -4, -9, 8, 4, -6,
    -- layer=1 filter=126 channel=78
    10, 5, 0, 9, -9, 10, 5, 0, -4,
    -- layer=1 filter=126 channel=79
    -11, 0, 7, 0, 6, -9, -10, -11, 4,
    -- layer=1 filter=126 channel=80
    9, -4, 11, -10, -1, -9, 5, 6, -9,
    -- layer=1 filter=126 channel=81
    9, 0, -2, 7, 2, -10, -10, 9, 0,
    -- layer=1 filter=126 channel=82
    0, 8, -5, -9, -10, 4, 3, -9, -3,
    -- layer=1 filter=126 channel=83
    6, 5, -3, 7, -11, 2, 0, -2, 8,
    -- layer=1 filter=126 channel=84
    6, -8, 6, -11, -5, -2, -6, 0, -1,
    -- layer=1 filter=126 channel=85
    0, 4, 7, 4, 0, -7, -1, -5, -9,
    -- layer=1 filter=126 channel=86
    5, 9, 2, 7, 0, -2, 4, -8, -4,
    -- layer=1 filter=126 channel=87
    3, 0, -8, 0, 0, -5, -5, -5, 7,
    -- layer=1 filter=126 channel=88
    -8, 3, -1, 5, -2, -3, -3, -2, -8,
    -- layer=1 filter=126 channel=89
    -4, -4, -7, -7, -3, 4, 0, -10, 3,
    -- layer=1 filter=126 channel=90
    -9, -8, 0, -11, -10, 5, 8, 9, 3,
    -- layer=1 filter=126 channel=91
    -2, 0, 5, 6, 0, 2, -7, -2, -3,
    -- layer=1 filter=126 channel=92
    0, 9, -9, -10, 5, -12, -5, -2, 6,
    -- layer=1 filter=126 channel=93
    -11, 3, -8, -5, 0, -2, -2, 6, -6,
    -- layer=1 filter=126 channel=94
    -8, -7, 4, -2, 3, 4, -9, -9, -6,
    -- layer=1 filter=126 channel=95
    -8, 6, -7, -2, 7, 3, 0, 8, -5,
    -- layer=1 filter=126 channel=96
    -1, -10, -7, -9, -2, 5, -3, -8, 10,
    -- layer=1 filter=126 channel=97
    6, -6, 5, -1, 0, 2, 6, -11, -7,
    -- layer=1 filter=126 channel=98
    -8, 5, -7, -3, -9, 3, 6, 6, 4,
    -- layer=1 filter=126 channel=99
    -5, 5, -4, -7, -7, 3, -8, -8, -11,
    -- layer=1 filter=126 channel=100
    7, -7, 2, -4, -9, -4, 9, 3, -4,
    -- layer=1 filter=126 channel=101
    7, -1, 8, -7, 6, 0, -6, -5, 3,
    -- layer=1 filter=126 channel=102
    0, -6, -1, -8, -10, 6, -2, -6, -4,
    -- layer=1 filter=126 channel=103
    -8, -10, -10, -6, 6, -6, 7, 6, -5,
    -- layer=1 filter=126 channel=104
    8, 3, -3, 3, 6, 0, 7, 7, 0,
    -- layer=1 filter=126 channel=105
    -6, -5, -9, -7, 9, -7, -11, 0, -8,
    -- layer=1 filter=126 channel=106
    -11, -8, -7, 7, 0, 4, -9, -1, 1,
    -- layer=1 filter=126 channel=107
    -6, 7, -5, 4, -6, -2, -5, 9, -2,
    -- layer=1 filter=126 channel=108
    -1, 0, 3, 5, -7, -6, -6, 6, -5,
    -- layer=1 filter=126 channel=109
    -5, 2, 3, -10, 7, -9, -7, 0, 3,
    -- layer=1 filter=126 channel=110
    -5, 3, -10, -9, -10, -1, -8, 0, 2,
    -- layer=1 filter=126 channel=111
    4, -8, -1, -7, -7, -8, 0, -6, -8,
    -- layer=1 filter=126 channel=112
    2, 0, -3, -5, 10, -5, 7, -2, 5,
    -- layer=1 filter=126 channel=113
    5, -9, -10, 0, -9, 2, -2, 7, -7,
    -- layer=1 filter=126 channel=114
    -11, 4, -1, 2, -4, 0, -5, -6, 1,
    -- layer=1 filter=126 channel=115
    4, -2, 1, 1, 6, -9, -7, -2, -11,
    -- layer=1 filter=126 channel=116
    5, 2, 7, -7, 7, -2, 4, 5, -1,
    -- layer=1 filter=126 channel=117
    -5, -6, -10, -7, 0, -1, 3, -7, -5,
    -- layer=1 filter=126 channel=118
    9, -8, -6, 5, 5, 2, -10, -4, 6,
    -- layer=1 filter=126 channel=119
    6, -13, 0, 1, 0, -12, 7, 6, 8,
    -- layer=1 filter=126 channel=120
    -3, 0, 0, -10, 5, 3, 4, 8, -1,
    -- layer=1 filter=126 channel=121
    6, -3, -5, -9, -8, -9, -6, -10, 2,
    -- layer=1 filter=126 channel=122
    9, -8, -5, 7, -7, -9, 4, -8, 0,
    -- layer=1 filter=126 channel=123
    1, -7, 7, -3, 0, 9, -8, -1, 11,
    -- layer=1 filter=126 channel=124
    -5, 0, -2, 11, 3, -1, 2, -1, -8,
    -- layer=1 filter=126 channel=125
    1, 7, 1, 4, -10, -8, 4, 1, -5,
    -- layer=1 filter=126 channel=126
    2, -4, -10, 4, -5, 4, 3, -11, 3,
    -- layer=1 filter=126 channel=127
    11, 6, 5, 2, -2, -9, 0, -3, -9,
    -- layer=1 filter=127 channel=0
    -13, -17, -6, -10, -9, -6, -12, -2, 4,
    -- layer=1 filter=127 channel=1
    -23, -12, -3, 0, -11, -9, -1, -2, -3,
    -- layer=1 filter=127 channel=2
    -7, -5, 4, 1, -10, -4, -1, 0, 6,
    -- layer=1 filter=127 channel=3
    1, 7, -9, -4, -2, -8, 8, -7, -6,
    -- layer=1 filter=127 channel=4
    6, -5, 1, -10, 7, 4, 7, -6, -6,
    -- layer=1 filter=127 channel=5
    -23, -24, -26, 4, 0, 2, 0, -21, -5,
    -- layer=1 filter=127 channel=6
    -15, -8, -6, 1, -4, 2, 1, -1, 0,
    -- layer=1 filter=127 channel=7
    -17, -21, 0, -16, -16, -4, -12, -8, -28,
    -- layer=1 filter=127 channel=8
    -25, -20, -22, -11, -3, 9, -17, -6, -20,
    -- layer=1 filter=127 channel=9
    -14, 5, 0, -14, 0, -2, -9, 13, -8,
    -- layer=1 filter=127 channel=10
    -26, -13, 7, -9, 0, 0, -8, -6, -22,
    -- layer=1 filter=127 channel=11
    -10, -12, 0, 3, -7, 3, 7, 5, 2,
    -- layer=1 filter=127 channel=12
    -8, -15, 11, -13, -11, -3, 18, 0, 4,
    -- layer=1 filter=127 channel=13
    -14, -5, -25, -17, 9, -18, -11, 8, -12,
    -- layer=1 filter=127 channel=14
    -1, -5, 4, -7, 15, 3, 10, 13, -16,
    -- layer=1 filter=127 channel=15
    -36, 0, -24, -12, 0, -7, -18, -6, -7,
    -- layer=1 filter=127 channel=16
    -14, -26, -16, 1, -19, 0, -17, -11, -11,
    -- layer=1 filter=127 channel=17
    -17, -14, -13, -6, -2, -10, -20, -12, -23,
    -- layer=1 filter=127 channel=18
    -9, 4, -3, -10, -1, 0, -5, 6, -14,
    -- layer=1 filter=127 channel=19
    -3, -16, 0, -17, 1, -14, -12, -4, -13,
    -- layer=1 filter=127 channel=20
    -19, -15, -16, -6, -15, -6, -24, -19, -19,
    -- layer=1 filter=127 channel=21
    -14, -7, -22, -13, -8, -8, -15, -17, -10,
    -- layer=1 filter=127 channel=22
    -31, -14, -10, -15, -17, -21, -26, -21, -11,
    -- layer=1 filter=127 channel=23
    -10, -9, 7, -15, -16, 4, 6, -21, 3,
    -- layer=1 filter=127 channel=24
    -6, -6, -18, -3, -11, -21, -12, -10, -3,
    -- layer=1 filter=127 channel=25
    -7, -3, -10, -3, -21, 4, -11, -19, -4,
    -- layer=1 filter=127 channel=26
    -10, 9, -12, -7, 12, -4, 1, 3, -14,
    -- layer=1 filter=127 channel=27
    10, 28, 18, 13, 14, 26, 20, 3, 10,
    -- layer=1 filter=127 channel=28
    -20, -13, -11, -2, -6, -9, -18, -11, -31,
    -- layer=1 filter=127 channel=29
    18, 24, 13, 14, 17, 27, 17, 25, 25,
    -- layer=1 filter=127 channel=30
    -16, -12, 0, 1, -14, -7, -6, -5, -8,
    -- layer=1 filter=127 channel=31
    -17, -17, -6, -8, -14, 2, 19, 12, -21,
    -- layer=1 filter=127 channel=32
    -21, 20, -11, 1, 0, -10, -12, 7, -21,
    -- layer=1 filter=127 channel=33
    -3, -6, 0, -8, -2, 3, 1, 9, 3,
    -- layer=1 filter=127 channel=34
    1, 0, 1, -12, -10, 3, 7, -11, 4,
    -- layer=1 filter=127 channel=35
    -3, -2, -2, -6, 4, 2, -11, 0, -6,
    -- layer=1 filter=127 channel=36
    -11, -4, -5, 0, 0, -6, 1, -13, -13,
    -- layer=1 filter=127 channel=37
    -23, -15, -19, -2, -13, -6, -18, -29, -15,
    -- layer=1 filter=127 channel=38
    -14, -19, -19, -23, -17, -19, -15, -12, -24,
    -- layer=1 filter=127 channel=39
    -10, -20, 0, -13, -12, -1, -19, -6, -14,
    -- layer=1 filter=127 channel=40
    -24, -13, -11, -5, -6, -11, -11, -20, -30,
    -- layer=1 filter=127 channel=41
    -3, -5, 10, 5, 6, -6, 9, 20, 6,
    -- layer=1 filter=127 channel=42
    -14, 0, -7, -7, 9, -6, 2, -7, -4,
    -- layer=1 filter=127 channel=43
    -9, -23, -18, -14, 0, 12, 0, -26, -15,
    -- layer=1 filter=127 channel=44
    -8, 11, -11, -9, 15, -6, -8, 1, -16,
    -- layer=1 filter=127 channel=45
    -20, -7, -17, -8, 5, -8, -17, -11, -5,
    -- layer=1 filter=127 channel=46
    -25, -6, -9, -8, -10, -9, -10, -2, -5,
    -- layer=1 filter=127 channel=47
    2, 0, -1, -1, -14, -10, 10, 2, 8,
    -- layer=1 filter=127 channel=48
    8, -1, -13, -1, 1, -2, -3, -21, -16,
    -- layer=1 filter=127 channel=49
    2, -11, -1, -5, 0, 2, 6, -3, -11,
    -- layer=1 filter=127 channel=50
    0, 4, -13, 1, -11, 2, 1, -2, -5,
    -- layer=1 filter=127 channel=51
    -8, -11, 6, 3, 8, -11, -11, -16, -25,
    -- layer=1 filter=127 channel=52
    -5, 9, 3, 7, -4, -9, -10, -8, 4,
    -- layer=1 filter=127 channel=53
    -6, 0, 3, -1, -2, -8, 4, -2, -1,
    -- layer=1 filter=127 channel=54
    -19, -4, -8, -10, -12, -4, -13, -11, -7,
    -- layer=1 filter=127 channel=55
    5, 6, -4, 2, -5, -10, 1, -9, 9,
    -- layer=1 filter=127 channel=56
    6, -2, 1, -5, 3, 4, 8, -6, 7,
    -- layer=1 filter=127 channel=57
    -9, -7, 2, -16, -9, -10, -14, -3, -22,
    -- layer=1 filter=127 channel=58
    -10, -19, 11, -9, -8, -3, 12, -16, 0,
    -- layer=1 filter=127 channel=59
    -9, 4, 4, -7, 8, -1, 2, 2, -2,
    -- layer=1 filter=127 channel=60
    6, 8, -11, -3, -7, -5, -2, 4, 0,
    -- layer=1 filter=127 channel=61
    8, 3, -4, 10, -4, 8, -4, 2, -4,
    -- layer=1 filter=127 channel=62
    -22, -22, -16, -16, -12, 0, -9, -13, -12,
    -- layer=1 filter=127 channel=63
    0, -10, 6, -10, 2, -9, -8, -13, -9,
    -- layer=1 filter=127 channel=64
    5, -2, 5, -12, -12, 1, -8, -3, 6,
    -- layer=1 filter=127 channel=65
    -10, -6, -6, -9, -1, -21, -10, -20, -10,
    -- layer=1 filter=127 channel=66
    2, 0, -6, -3, -7, -9, -15, -10, -9,
    -- layer=1 filter=127 channel=67
    4, 13, -2, -10, 14, -5, -2, -12, -8,
    -- layer=1 filter=127 channel=68
    -1, 9, -16, -11, 10, -16, -10, -7, -17,
    -- layer=1 filter=127 channel=69
    -19, -12, -4, 0, 11, -2, -20, -4, 1,
    -- layer=1 filter=127 channel=70
    6, -11, -4, 7, -14, 6, 3, -4, 2,
    -- layer=1 filter=127 channel=71
    -10, -12, -19, -21, -21, -12, -4, -4, -16,
    -- layer=1 filter=127 channel=72
    0, -7, -8, -4, -9, -14, 11, 1, 0,
    -- layer=1 filter=127 channel=73
    -5, -6, 0, 2, 5, -9, 1, 1, -10,
    -- layer=1 filter=127 channel=74
    4, 0, -4, -1, -7, -1, -3, -1, -11,
    -- layer=1 filter=127 channel=75
    0, 0, 8, 0, -8, 1, -7, -11, -4,
    -- layer=1 filter=127 channel=76
    0, 5, -5, -8, -2, -14, -12, -12, -18,
    -- layer=1 filter=127 channel=77
    2, -3, -9, 0, -1, -14, -6, -10, -7,
    -- layer=1 filter=127 channel=78
    -3, -1, 6, -10, -5, -4, -11, -4, 6,
    -- layer=1 filter=127 channel=79
    -32, -24, -20, -7, -1, -1, -11, -11, -16,
    -- layer=1 filter=127 channel=80
    7, 9, 4, 4, 0, 8, -2, 2, 6,
    -- layer=1 filter=127 channel=81
    -22, -5, 0, -10, -11, -13, -4, -6, -14,
    -- layer=1 filter=127 channel=82
    4, -11, -17, -16, -8, -3, -11, -1, -5,
    -- layer=1 filter=127 channel=83
    -22, -1, -11, -16, 4, 7, -6, 3, -1,
    -- layer=1 filter=127 channel=84
    -8, 0, 0, 2, -18, -2, 0, -8, -17,
    -- layer=1 filter=127 channel=85
    -15, -7, 14, -10, -17, 1, 6, -9, -2,
    -- layer=1 filter=127 channel=86
    -11, -9, -6, -8, -9, 1, -11, 0, -3,
    -- layer=1 filter=127 channel=87
    -9, -1, 3, 0, -15, -16, -2, -11, 0,
    -- layer=1 filter=127 channel=88
    7, -8, 0, 14, 7, -10, -11, 0, -5,
    -- layer=1 filter=127 channel=89
    1, -2, -13, -8, -7, -5, -21, -1, -22,
    -- layer=1 filter=127 channel=90
    -6, 18, -21, -18, 12, -5, -8, 5, -8,
    -- layer=1 filter=127 channel=91
    -10, -25, -17, -15, -16, -16, -20, -13, -30,
    -- layer=1 filter=127 channel=92
    -5, 12, -24, -10, 17, -5, -11, 12, -7,
    -- layer=1 filter=127 channel=93
    -19, -12, -8, -9, -6, -7, -8, -25, -10,
    -- layer=1 filter=127 channel=94
    -14, -17, -16, -10, -20, -16, -6, -10, -4,
    -- layer=1 filter=127 channel=95
    -7, -9, -8, 0, -2, 2, -4, -13, -24,
    -- layer=1 filter=127 channel=96
    -7, -8, 5, 5, 8, -6, 0, -7, -10,
    -- layer=1 filter=127 channel=97
    -3, -10, -7, -4, -9, -18, -4, -5, -10,
    -- layer=1 filter=127 channel=98
    -32, -30, -18, -15, -14, -12, -7, -5, -15,
    -- layer=1 filter=127 channel=99
    -18, -6, -8, -21, -3, -12, -2, -9, -19,
    -- layer=1 filter=127 channel=100
    -10, -6, 4, 0, -6, 7, 5, 3, -2,
    -- layer=1 filter=127 channel=101
    -18, -5, -14, -26, -24, -11, -27, -11, -17,
    -- layer=1 filter=127 channel=102
    -22, -26, -26, -13, -14, -19, -8, -9, -28,
    -- layer=1 filter=127 channel=103
    21, 21, 7, 14, 0, 2, 21, 5, 12,
    -- layer=1 filter=127 channel=104
    -2, 3, 3, -12, 0, -4, 2, 9, 5,
    -- layer=1 filter=127 channel=105
    -5, -13, -16, -2, -17, -17, -18, -11, -3,
    -- layer=1 filter=127 channel=106
    -3, 10, -18, -4, -5, -2, -12, -12, -25,
    -- layer=1 filter=127 channel=107
    2, -6, -1, 9, 0, -8, -10, -3, 5,
    -- layer=1 filter=127 channel=108
    -8, 3, -2, 5, 15, -10, 3, 8, -12,
    -- layer=1 filter=127 channel=109
    1, -5, -1, 2, 8, -3, -3, -1, 10,
    -- layer=1 filter=127 channel=110
    7, 1, 4, 3, -8, -13, 1, -6, -1,
    -- layer=1 filter=127 channel=111
    -24, -3, -9, -14, -7, -7, 0, -10, -22,
    -- layer=1 filter=127 channel=112
    0, 2, 0, -10, -7, -14, -12, -3, -18,
    -- layer=1 filter=127 channel=113
    -1, -3, -15, -9, 3, -8, -21, -19, -5,
    -- layer=1 filter=127 channel=114
    -13, 1, -15, 10, 8, 5, -8, -19, 1,
    -- layer=1 filter=127 channel=115
    -12, -9, -11, -5, -5, -17, -5, -4, -13,
    -- layer=1 filter=127 channel=116
    8, -8, 7, 7, -2, 9, -2, -5, 5,
    -- layer=1 filter=127 channel=117
    -22, -11, -11, -8, 4, -11, -1, -8, -20,
    -- layer=1 filter=127 channel=118
    -21, -12, -3, -10, -14, -12, 0, -13, -16,
    -- layer=1 filter=127 channel=119
    -2, 0, -1, -12, -3, -2, -4, -3, -11,
    -- layer=1 filter=127 channel=120
    -12, -7, 2, -15, -11, -19, -3, -18, -21,
    -- layer=1 filter=127 channel=121
    -13, 3, 0, -7, 5, -6, -11, -11, -10,
    -- layer=1 filter=127 channel=122
    10, 7, 5, 4, 7, -7, 5, 6, 0,
    -- layer=1 filter=127 channel=123
    1, 0, 13, 3, -4, 5, -5, 2, -9,
    -- layer=1 filter=127 channel=124
    -1, -6, -1, -10, 10, 7, -6, -8, -6,
    -- layer=1 filter=127 channel=125
    3, -4, 11, -5, -11, 0, -12, 2, 3,
    -- layer=1 filter=127 channel=126
    -13, -22, -17, -9, -8, 2, -11, 0, 11,
    -- layer=1 filter=127 channel=127
    -18, 4, -7, -7, -1, -6, 0, -5, -17,
    -- layer=1 filter=128 channel=0
    -6, 0, -1, 1, 5, 4, -3, -4, 0,
    -- layer=1 filter=128 channel=1
    -2, 1, 6, -4, -6, -11, -2, -8, 0,
    -- layer=1 filter=128 channel=2
    -8, -10, 0, 0, -4, 3, 1, -8, -7,
    -- layer=1 filter=128 channel=3
    5, -3, 5, -8, -10, 4, -11, -2, 5,
    -- layer=1 filter=128 channel=4
    0, 6, -2, -9, 8, 1, 0, -6, -11,
    -- layer=1 filter=128 channel=5
    -6, 1, 6, -9, -10, 9, 5, 1, -9,
    -- layer=1 filter=128 channel=6
    -1, 6, 0, -12, 3, -7, -11, -10, 3,
    -- layer=1 filter=128 channel=7
    -10, -8, 0, 1, 4, -5, -12, -14, -5,
    -- layer=1 filter=128 channel=8
    -10, -1, 2, -2, 6, 8, 3, -1, -6,
    -- layer=1 filter=128 channel=9
    -6, 0, 7, 0, 1, -6, -2, 1, 4,
    -- layer=1 filter=128 channel=10
    5, -3, 3, 0, 2, -7, -8, 6, -10,
    -- layer=1 filter=128 channel=11
    9, -3, -12, -5, 2, -5, 4, -3, 9,
    -- layer=1 filter=128 channel=12
    -9, -2, -8, -2, 1, 10, -8, -3, 6,
    -- layer=1 filter=128 channel=13
    1, -4, 1, -7, 0, -9, -5, -4, -9,
    -- layer=1 filter=128 channel=14
    -10, -6, -4, 5, -14, -8, 0, 2, 3,
    -- layer=1 filter=128 channel=15
    -6, 10, 9, 7, 2, -2, -7, -2, -5,
    -- layer=1 filter=128 channel=16
    0, -2, -4, 2, -2, -6, 4, -2, -1,
    -- layer=1 filter=128 channel=17
    0, -5, 0, -11, -10, 5, 7, 7, -4,
    -- layer=1 filter=128 channel=18
    -8, 10, 2, 8, -10, 0, 1, 6, -1,
    -- layer=1 filter=128 channel=19
    2, 2, 0, 8, 0, -11, 8, 7, -11,
    -- layer=1 filter=128 channel=20
    8, -10, 1, 7, -10, -11, 1, -5, -6,
    -- layer=1 filter=128 channel=21
    7, -2, 6, -7, -9, 0, 1, -3, 9,
    -- layer=1 filter=128 channel=22
    -8, 1, -1, 5, -3, -11, -2, 7, -11,
    -- layer=1 filter=128 channel=23
    -7, 0, 7, -10, 1, 4, -6, -2, -1,
    -- layer=1 filter=128 channel=24
    -6, -5, -7, 9, 6, 0, -4, 5, -4,
    -- layer=1 filter=128 channel=25
    9, 2, -3, 2, -8, -10, 6, 0, -7,
    -- layer=1 filter=128 channel=26
    1, -2, -1, 0, 5, 6, -7, 6, -1,
    -- layer=1 filter=128 channel=27
    0, -3, 2, -1, -6, 9, -7, -8, 8,
    -- layer=1 filter=128 channel=28
    5, 6, 0, -6, -1, 0, -8, 2, 5,
    -- layer=1 filter=128 channel=29
    -11, 3, -8, 5, -11, 0, -5, -3, 1,
    -- layer=1 filter=128 channel=30
    1, 5, -8, -9, 4, 0, 3, -8, -2,
    -- layer=1 filter=128 channel=31
    -9, -3, 5, 1, 5, 2, 5, -4, -9,
    -- layer=1 filter=128 channel=32
    -11, -6, 2, -11, 5, -4, -4, 2, 3,
    -- layer=1 filter=128 channel=33
    -8, -3, 0, 11, 7, -4, 11, -7, 4,
    -- layer=1 filter=128 channel=34
    5, -6, 0, 8, 7, 4, -8, 4, -7,
    -- layer=1 filter=128 channel=35
    10, -7, -6, 7, -5, 9, -1, -4, -8,
    -- layer=1 filter=128 channel=36
    -10, -4, -2, -3, -5, 1, 7, -1, 2,
    -- layer=1 filter=128 channel=37
    -6, 4, -12, -1, -6, -4, -9, -3, -1,
    -- layer=1 filter=128 channel=38
    5, -9, 3, -11, -2, -6, -8, 1, -4,
    -- layer=1 filter=128 channel=39
    -10, 0, -9, -9, 1, -1, 8, -5, 6,
    -- layer=1 filter=128 channel=40
    -5, 1, -7, 7, -11, -3, 0, 6, -10,
    -- layer=1 filter=128 channel=41
    -4, -3, -3, 8, 9, 7, -6, 8, -5,
    -- layer=1 filter=128 channel=42
    0, -8, 6, 5, 9, -6, -7, -7, -3,
    -- layer=1 filter=128 channel=43
    -5, -5, 0, 3, 5, 2, 9, -11, -4,
    -- layer=1 filter=128 channel=44
    -2, 1, 4, 5, 4, 9, -8, -7, 2,
    -- layer=1 filter=128 channel=45
    5, 6, -3, 5, -7, 3, 0, 4, -4,
    -- layer=1 filter=128 channel=46
    4, 3, -9, -9, -4, 9, -6, -6, -7,
    -- layer=1 filter=128 channel=47
    0, 9, -2, 0, -11, -4, -4, -3, -3,
    -- layer=1 filter=128 channel=48
    -9, -8, -1, 1, 3, 5, -10, -6, -1,
    -- layer=1 filter=128 channel=49
    -9, -7, 1, -4, 0, -12, 6, 2, -1,
    -- layer=1 filter=128 channel=50
    0, -7, 7, 0, 4, 0, -2, -2, 8,
    -- layer=1 filter=128 channel=51
    -5, 0, 3, 0, -7, -8, -7, 5, 6,
    -- layer=1 filter=128 channel=52
    7, -8, 5, 6, 11, 3, -9, 4, -10,
    -- layer=1 filter=128 channel=53
    -7, 7, 4, -2, -7, -1, -4, -9, 7,
    -- layer=1 filter=128 channel=54
    6, -4, -3, -1, 0, -4, 11, -6, -5,
    -- layer=1 filter=128 channel=55
    0, 6, -9, -11, 2, -2, 8, -5, 2,
    -- layer=1 filter=128 channel=56
    -6, 0, 9, 7, 6, 6, -2, 3, -3,
    -- layer=1 filter=128 channel=57
    -5, 0, 6, 3, -6, -6, 7, 7, -11,
    -- layer=1 filter=128 channel=58
    4, -2, 5, 1, 0, 0, -9, 2, -6,
    -- layer=1 filter=128 channel=59
    6, 2, 8, -8, -9, -1, 5, -9, -8,
    -- layer=1 filter=128 channel=60
    -1, -8, -9, 8, 4, -4, 0, 2, -8,
    -- layer=1 filter=128 channel=61
    7, 0, -3, 10, 1, 1, 8, 8, -4,
    -- layer=1 filter=128 channel=62
    10, -2, 1, -10, -10, -4, -7, 1, -3,
    -- layer=1 filter=128 channel=63
    7, 1, -4, 0, 9, 0, 5, 10, 0,
    -- layer=1 filter=128 channel=64
    -5, -10, -1, -5, -8, -7, 5, 8, 8,
    -- layer=1 filter=128 channel=65
    6, -11, 0, -7, 1, -8, -2, 6, -4,
    -- layer=1 filter=128 channel=66
    8, -10, -2, 6, -3, 1, 9, -4, -9,
    -- layer=1 filter=128 channel=67
    -6, 0, 0, 1, 0, 5, 6, -5, -1,
    -- layer=1 filter=128 channel=68
    1, 5, -3, -7, -3, 0, 10, 3, -6,
    -- layer=1 filter=128 channel=69
    5, 0, 0, -9, -5, -4, -8, -5, -3,
    -- layer=1 filter=128 channel=70
    1, -3, 3, -2, 0, -9, 5, 4, 3,
    -- layer=1 filter=128 channel=71
    4, -13, -8, -10, -6, 7, 6, 3, 1,
    -- layer=1 filter=128 channel=72
    8, -11, 4, -7, -7, 1, 0, -4, 8,
    -- layer=1 filter=128 channel=73
    -4, 0, -8, 0, -7, 6, 7, -1, -3,
    -- layer=1 filter=128 channel=74
    -4, -8, 1, -9, 2, 0, 5, 2, -3,
    -- layer=1 filter=128 channel=75
    5, -3, -6, -9, 4, -11, -5, 5, 5,
    -- layer=1 filter=128 channel=76
    0, -1, -3, -6, 0, 2, -6, -8, -2,
    -- layer=1 filter=128 channel=77
    -6, 0, 4, -1, 1, -1, -5, -5, 4,
    -- layer=1 filter=128 channel=78
    -10, -9, -8, 3, 7, 8, -5, 5, 5,
    -- layer=1 filter=128 channel=79
    3, -6, -8, 0, -2, -5, -2, -8, 7,
    -- layer=1 filter=128 channel=80
    3, 11, -7, 7, 8, -4, 5, 7, 8,
    -- layer=1 filter=128 channel=81
    0, -3, 0, 9, 7, -8, 6, -5, -3,
    -- layer=1 filter=128 channel=82
    -9, -8, 2, -7, 0, 4, -3, 2, 8,
    -- layer=1 filter=128 channel=83
    -4, -4, -10, 4, 5, -11, 5, -10, 0,
    -- layer=1 filter=128 channel=84
    4, 6, -4, -7, -3, -9, -1, -9, 8,
    -- layer=1 filter=128 channel=85
    -10, 0, -9, 8, -6, -6, -10, -8, 2,
    -- layer=1 filter=128 channel=86
    4, -8, -12, -5, -5, -9, -1, -5, 1,
    -- layer=1 filter=128 channel=87
    -9, 3, 2, 5, 1, 0, -2, -4, -8,
    -- layer=1 filter=128 channel=88
    2, -5, 11, -4, -3, 2, 0, -8, 2,
    -- layer=1 filter=128 channel=89
    0, -11, -3, 4, -3, -7, 8, -5, -5,
    -- layer=1 filter=128 channel=90
    -12, -9, 1, 5, -5, -5, -4, -8, -7,
    -- layer=1 filter=128 channel=91
    5, 4, 5, 6, -5, 5, 2, 5, -6,
    -- layer=1 filter=128 channel=92
    0, -12, 4, 2, 3, 4, 5, 2, -9,
    -- layer=1 filter=128 channel=93
    -6, 3, -3, 4, 0, -9, -3, -12, -4,
    -- layer=1 filter=128 channel=94
    -4, -4, -11, -12, -11, -7, -11, 0, 0,
    -- layer=1 filter=128 channel=95
    2, 2, -6, 5, 1, 5, -9, -10, 5,
    -- layer=1 filter=128 channel=96
    -3, -10, -10, -1, 8, -12, -11, -1, 0,
    -- layer=1 filter=128 channel=97
    1, 3, 1, 3, 0, 8, 4, -5, -3,
    -- layer=1 filter=128 channel=98
    -9, -1, 5, -10, -10, 2, -9, 10, -1,
    -- layer=1 filter=128 channel=99
    9, 6, 5, 3, 1, 2, -4, 2, -11,
    -- layer=1 filter=128 channel=100
    2, -8, -11, 4, 2, -9, 0, -9, -8,
    -- layer=1 filter=128 channel=101
    7, -8, -4, 5, 0, -11, 4, -3, -1,
    -- layer=1 filter=128 channel=102
    0, 7, -6, -2, -3, 6, -4, 0, 0,
    -- layer=1 filter=128 channel=103
    -1, 7, 4, 6, 6, -8, -2, -8, -3,
    -- layer=1 filter=128 channel=104
    -1, 7, 0, -5, -3, -10, -1, 1, 5,
    -- layer=1 filter=128 channel=105
    -7, -10, -3, -12, -1, -2, 2, -2, -9,
    -- layer=1 filter=128 channel=106
    4, 6, -1, -4, 8, 8, -3, -10, -10,
    -- layer=1 filter=128 channel=107
    -4, -7, 4, -7, -9, 0, 3, -11, 10,
    -- layer=1 filter=128 channel=108
    -5, -7, -11, -1, -9, -8, 6, -7, -1,
    -- layer=1 filter=128 channel=109
    -4, -1, 11, 0, 6, -1, 2, -2, -1,
    -- layer=1 filter=128 channel=110
    -10, 0, -6, 5, 1, 1, -7, -1, -2,
    -- layer=1 filter=128 channel=111
    8, -2, 5, -1, -8, 5, 2, 5, -1,
    -- layer=1 filter=128 channel=112
    0, 0, -12, 1, 6, 4, -5, 0, -3,
    -- layer=1 filter=128 channel=113
    -8, -2, 10, 7, 3, 9, 1, -3, 6,
    -- layer=1 filter=128 channel=114
    -8, -1, -1, -8, 2, 0, 8, -1, 0,
    -- layer=1 filter=128 channel=115
    -1, 7, -7, 4, 7, 4, 3, 2, 0,
    -- layer=1 filter=128 channel=116
    -6, -4, -3, -4, -1, 10, 5, 1, 3,
    -- layer=1 filter=128 channel=117
    4, -3, 3, -9, 1, 10, -5, 9, -2,
    -- layer=1 filter=128 channel=118
    -2, -1, 1, 5, 5, -2, -7, 6, 7,
    -- layer=1 filter=128 channel=119
    8, 5, -3, -1, -9, 8, -8, -9, -1,
    -- layer=1 filter=128 channel=120
    -4, -5, 0, 7, -11, 5, 1, 6, -1,
    -- layer=1 filter=128 channel=121
    5, -1, 8, -3, -2, -10, -11, -5, -4,
    -- layer=1 filter=128 channel=122
    -5, 3, -10, 8, 5, -4, -5, 5, 3,
    -- layer=1 filter=128 channel=123
    -11, 8, -3, 0, 4, 7, -6, 2, -2,
    -- layer=1 filter=128 channel=124
    0, 3, 2, -2, -2, -5, 9, 0, -4,
    -- layer=1 filter=128 channel=125
    4, 1, -3, 3, 5, -8, -6, 4, -7,
    -- layer=1 filter=128 channel=126
    7, 0, 7, 0, -2, -5, -9, -1, 5,
    -- layer=1 filter=128 channel=127
    -9, -8, 9, 2, 0, -8, 0, 8, -2,
    -- layer=1 filter=129 channel=0
    -12, -18, -3, 10, -3, 7, 8, -8, 1,
    -- layer=1 filter=129 channel=1
    -10, 1, -20, -7, -24, 9, 40, 16, 18,
    -- layer=1 filter=129 channel=2
    37, -20, -48, 31, -5, -21, 14, -33, -21,
    -- layer=1 filter=129 channel=3
    -4, 1, -15, -2, -4, -3, -17, 5, -12,
    -- layer=1 filter=129 channel=4
    3, 3, -3, 5, 0, -2, -1, 5, 0,
    -- layer=1 filter=129 channel=5
    -10, -14, -45, -29, -32, 3, 41, 10, 14,
    -- layer=1 filter=129 channel=6
    -4, -2, 5, -2, -16, -7, -23, -36, -6,
    -- layer=1 filter=129 channel=7
    -2, 36, 8, -7, 3, 29, -15, 0, -3,
    -- layer=1 filter=129 channel=8
    -11, -22, -49, -19, -32, 1, 18, 3, 11,
    -- layer=1 filter=129 channel=9
    -32, -51, -1, -46, -27, -9, 8, -18, 40,
    -- layer=1 filter=129 channel=10
    13, 29, 2, -6, 0, 14, -20, 12, -10,
    -- layer=1 filter=129 channel=11
    -10, -21, -7, -6, 3, -12, -8, 1, -17,
    -- layer=1 filter=129 channel=12
    -42, -51, -13, -30, -64, -13, -16, -36, -16,
    -- layer=1 filter=129 channel=13
    15, -6, 3, 0, 3, -11, 8, -17, 8,
    -- layer=1 filter=129 channel=14
    -7, 28, 13, 7, -24, -13, -12, -11, -4,
    -- layer=1 filter=129 channel=15
    -34, -60, -1, -42, -69, 14, 13, -52, -6,
    -- layer=1 filter=129 channel=16
    -18, -17, -39, -20, -21, 6, 20, -8, 24,
    -- layer=1 filter=129 channel=17
    8, -4, -14, 2, -2, 8, 12, 10, -5,
    -- layer=1 filter=129 channel=18
    -64, -58, -42, 27, -13, -14, 13, 8, 30,
    -- layer=1 filter=129 channel=19
    0, -45, 6, -13, 0, 6, 36, 5, 66,
    -- layer=1 filter=129 channel=20
    9, 20, 1, 8, 5, -5, 0, 8, -3,
    -- layer=1 filter=129 channel=21
    -10, 6, -7, -19, 1, -9, -12, 0, -4,
    -- layer=1 filter=129 channel=22
    0, 10, 5, -7, -13, -2, 16, 7, -8,
    -- layer=1 filter=129 channel=23
    -5, -30, 12, -21, -3, 20, 17, -38, 24,
    -- layer=1 filter=129 channel=24
    -28, -23, -11, -25, -7, 2, -15, -4, 14,
    -- layer=1 filter=129 channel=25
    20, 39, 8, -17, 8, 13, 19, 18, 17,
    -- layer=1 filter=129 channel=26
    -5, 0, 3, -16, -3, -3, 5, -12, -1,
    -- layer=1 filter=129 channel=27
    -7, -22, -35, -14, -4, -25, -33, -45, -38,
    -- layer=1 filter=129 channel=28
    15, 35, 4, -3, -2, 15, -16, 5, 7,
    -- layer=1 filter=129 channel=29
    12, 3, 3, 0, -1, -8, -26, -6, -4,
    -- layer=1 filter=129 channel=30
    -60, -64, -43, -13, -6, -19, 24, 14, 35,
    -- layer=1 filter=129 channel=31
    -3, -12, -9, -13, -18, -2, -9, -4, 6,
    -- layer=1 filter=129 channel=32
    -24, 19, 2, -28, 16, -8, 0, -3, 15,
    -- layer=1 filter=129 channel=33
    -4, -1, -4, 5, 8, -12, 0, 9, 0,
    -- layer=1 filter=129 channel=34
    -5, -25, 7, -7, -9, 12, 5, -4, 31,
    -- layer=1 filter=129 channel=35
    17, -2, 13, 17, 18, 8, -1, 10, 11,
    -- layer=1 filter=129 channel=36
    -9, -19, -16, -8, -15, -8, -16, -11, -22,
    -- layer=1 filter=129 channel=37
    -6, -31, -23, -23, -18, 0, 38, 6, 11,
    -- layer=1 filter=129 channel=38
    16, 5, -5, 1, 1, -10, 5, -4, 1,
    -- layer=1 filter=129 channel=39
    -15, -10, -16, -8, -27, -9, -17, -11, -1,
    -- layer=1 filter=129 channel=40
    11, 7, 2, -2, -14, 1, -6, -8, 15,
    -- layer=1 filter=129 channel=41
    -11, -16, 57, -7, -19, 10, -19, -30, 41,
    -- layer=1 filter=129 channel=42
    60, -29, -43, 36, -15, -17, 16, -5, -28,
    -- layer=1 filter=129 channel=43
    -13, -2, -48, -24, -28, 1, 15, -7, 23,
    -- layer=1 filter=129 channel=44
    0, 12, 2, -12, 1, 3, 6, 13, 2,
    -- layer=1 filter=129 channel=45
    3, -7, -17, -21, -18, -12, 7, -19, -4,
    -- layer=1 filter=129 channel=46
    8, -17, -8, 4, -27, -19, 34, 0, 19,
    -- layer=1 filter=129 channel=47
    -28, -35, 26, -33, -39, 0, 12, -56, 8,
    -- layer=1 filter=129 channel=48
    -8, 1, -10, 7, -2, -2, 2, 1, 2,
    -- layer=1 filter=129 channel=49
    17, -16, -8, 0, -27, 7, -8, -23, 6,
    -- layer=1 filter=129 channel=50
    -18, -6, -13, -4, -14, -7, -19, -2, 3,
    -- layer=1 filter=129 channel=51
    15, 24, 5, -3, -4, 0, 4, -3, -16,
    -- layer=1 filter=129 channel=52
    9, -3, 1, 4, 4, -3, 4, 1, 11,
    -- layer=1 filter=129 channel=53
    -2, 1, -1, 9, -5, 0, 7, 5, 5,
    -- layer=1 filter=129 channel=54
    28, 26, -11, -2, 11, 17, 16, 16, 5,
    -- layer=1 filter=129 channel=55
    3, -1, 6, -9, 0, -4, -22, -7, -17,
    -- layer=1 filter=129 channel=56
    10, 5, -11, 2, 8, -11, -2, 4, -7,
    -- layer=1 filter=129 channel=57
    26, 24, 9, 5, 6, 22, -14, 3, -28,
    -- layer=1 filter=129 channel=58
    -7, 3, 5, -24, -3, 23, -4, 4, -22,
    -- layer=1 filter=129 channel=59
    -2, 2, 7, 17, -1, 16, 7, 0, 0,
    -- layer=1 filter=129 channel=60
    -6, 3, -1, -1, -12, -6, -13, -3, -15,
    -- layer=1 filter=129 channel=61
    5, -5, -2, 1, 6, -13, -7, 0, -5,
    -- layer=1 filter=129 channel=62
    -9, -25, -37, 0, -12, 10, 34, -2, 17,
    -- layer=1 filter=129 channel=63
    -26, -10, -9, 2, -5, -12, 2, -7, 4,
    -- layer=1 filter=129 channel=64
    -6, 6, 0, -8, -15, 5, -8, -4, 7,
    -- layer=1 filter=129 channel=65
    0, 3, -2, -2, 3, -1, 6, 11, 3,
    -- layer=1 filter=129 channel=66
    -12, -6, -10, -5, 0, 14, -1, -7, 3,
    -- layer=1 filter=129 channel=67
    27, 13, 11, 0, -15, -8, -30, -33, -33,
    -- layer=1 filter=129 channel=68
    1, 25, -9, -34, 18, -16, -12, 17, 3,
    -- layer=1 filter=129 channel=69
    -4, -20, -6, -38, -15, -12, 33, -27, 2,
    -- layer=1 filter=129 channel=70
    -18, -28, -13, -25, -41, -16, -42, -60, -29,
    -- layer=1 filter=129 channel=71
    0, 2, -15, -19, 3, -3, -3, 15, 22,
    -- layer=1 filter=129 channel=72
    -51, -58, -22, -37, -29, 0, 21, -18, 42,
    -- layer=1 filter=129 channel=73
    -5, -13, 2, -5, 0, -6, -4, 8, 8,
    -- layer=1 filter=129 channel=74
    -3, -11, -20, -2, 24, -19, 11, 24, 30,
    -- layer=1 filter=129 channel=75
    -65, -55, -49, 2, -61, -47, 19, 0, 26,
    -- layer=1 filter=129 channel=76
    6, -10, -6, 13, 15, -21, 12, 6, 7,
    -- layer=1 filter=129 channel=77
    -16, -14, -6, -1, -5, 3, -4, 0, 5,
    -- layer=1 filter=129 channel=78
    9, -3, -2, 9, -5, 16, -13, 5, -9,
    -- layer=1 filter=129 channel=79
    -7, -33, -18, -23, -29, 7, 33, -6, 5,
    -- layer=1 filter=129 channel=80
    0, 0, -1, -10, 9, 8, -8, 8, -6,
    -- layer=1 filter=129 channel=81
    -22, -12, -12, -17, 2, -2, 0, 5, 5,
    -- layer=1 filter=129 channel=82
    2, 9, 0, -14, -15, 0, -1, -8, -6,
    -- layer=1 filter=129 channel=83
    -3, -19, -6, -21, -36, -11, 6, -14, 6,
    -- layer=1 filter=129 channel=84
    -38, -29, -11, 13, 3, -5, 24, 21, 58,
    -- layer=1 filter=129 channel=85
    -7, -13, 23, -20, -4, 23, 5, -29, 16,
    -- layer=1 filter=129 channel=86
    8, 1, -6, 13, 3, 8, 8, -5, 9,
    -- layer=1 filter=129 channel=87
    2, 4, 5, -56, -32, 24, 3, -57, 20,
    -- layer=1 filter=129 channel=88
    -10, 0, -16, -6, -16, -18, -1, -17, -5,
    -- layer=1 filter=129 channel=89
    -11, 4, 4, -3, -15, -3, 1, 0, 15,
    -- layer=1 filter=129 channel=90
    -3, 19, -2, -18, -6, -13, 7, -3, -23,
    -- layer=1 filter=129 channel=91
    20, 5, 1, 10, 1, -12, 2, 8, -8,
    -- layer=1 filter=129 channel=92
    -68, -59, 2, -107, -66, -25, -48, -38, -40,
    -- layer=1 filter=129 channel=93
    -1, 10, 2, 6, 2, 13, 1, 0, 2,
    -- layer=1 filter=129 channel=94
    -10, -21, -13, 3, -16, 10, -9, -11, -4,
    -- layer=1 filter=129 channel=95
    -56, -70, -26, 18, -13, -12, 24, 20, 46,
    -- layer=1 filter=129 channel=96
    -13, -12, 8, -10, 7, -4, -10, -5, -3,
    -- layer=1 filter=129 channel=97
    0, -11, 4, 3, -8, 5, 0, 0, -3,
    -- layer=1 filter=129 channel=98
    1, -4, -26, -7, -25, 2, 28, 3, 6,
    -- layer=1 filter=129 channel=99
    -6, 0, 3, 5, 10, 13, -19, 13, -24,
    -- layer=1 filter=129 channel=100
    2, -8, -14, -13, 0, -23, -9, 2, -4,
    -- layer=1 filter=129 channel=101
    16, 11, 8, 15, -2, 1, 8, 4, 8,
    -- layer=1 filter=129 channel=102
    -1, -7, -16, 6, 1, -14, -3, 4, 4,
    -- layer=1 filter=129 channel=103
    -11, -5, -12, -3, -21, -9, -29, -17, -1,
    -- layer=1 filter=129 channel=104
    -18, -10, 5, 2, -33, 25, 10, -52, -2,
    -- layer=1 filter=129 channel=105
    1, 0, 5, -4, 8, 3, -5, 7, 11,
    -- layer=1 filter=129 channel=106
    12, 11, 0, 0, -11, -14, -10, -11, 10,
    -- layer=1 filter=129 channel=107
    -17, -18, -9, -2, -3, -2, -3, -7, 0,
    -- layer=1 filter=129 channel=108
    1, 6, 12, -25, -10, 1, -20, -39, -9,
    -- layer=1 filter=129 channel=109
    3, 6, 1, -10, -2, 0, 9, -5, 2,
    -- layer=1 filter=129 channel=110
    4, 7, -1, 5, 1, 2, -1, -10, 4,
    -- layer=1 filter=129 channel=111
    -52, -56, -30, 28, 1, 4, 23, 19, 49,
    -- layer=1 filter=129 channel=112
    -23, -18, -13, 31, -2, -5, 23, 22, 33,
    -- layer=1 filter=129 channel=113
    10, -12, -26, -1, -21, -19, -8, -15, 0,
    -- layer=1 filter=129 channel=114
    -69, -61, -64, -64, -84, -63, -17, -48, -19,
    -- layer=1 filter=129 channel=115
    10, 1, 10, 3, -5, 17, -5, 1, -4,
    -- layer=1 filter=129 channel=116
    -10, 7, 4, 1, -9, 2, -2, -4, 3,
    -- layer=1 filter=129 channel=117
    0, -17, -13, 36, -3, -13, 5, 50, 3,
    -- layer=1 filter=129 channel=118
    -21, -30, -16, 16, 4, -4, 17, 18, 45,
    -- layer=1 filter=129 channel=119
    -24, 2, 16, -26, 2, 1, -17, -2, 3,
    -- layer=1 filter=129 channel=120
    12, 13, 1, -11, 0, -11, 0, -6, -12,
    -- layer=1 filter=129 channel=121
    -10, -25, -23, -22, -41, -34, 14, 4, -10,
    -- layer=1 filter=129 channel=122
    1, 2, 6, -1, 2, -3, 8, 3, 0,
    -- layer=1 filter=129 channel=123
    -22, -40, -35, -20, -23, -27, 1, -16, 7,
    -- layer=1 filter=129 channel=124
    -15, -2, -14, 0, 1, 0, -14, 0, -15,
    -- layer=1 filter=129 channel=125
    31, 22, 0, -6, -21, -21, -28, -16, -46,
    -- layer=1 filter=129 channel=126
    -6, -12, -14, -35, -18, -2, 7, -12, -2,
    -- layer=1 filter=129 channel=127
    -42, -54, -24, 23, 8, -5, 20, 15, 43,
    -- layer=1 filter=130 channel=0
    -4, -4, 7, -8, -10, 6, 2, -7, 5,
    -- layer=1 filter=130 channel=1
    -7, 2, -7, -11, -1, 7, 4, 3, -11,
    -- layer=1 filter=130 channel=2
    0, 9, 5, 1, 0, 7, 9, 8, -4,
    -- layer=1 filter=130 channel=3
    -9, 0, -8, 3, 2, -3, -7, 0, 4,
    -- layer=1 filter=130 channel=4
    -7, 2, -8, 0, 0, -3, -9, -3, -5,
    -- layer=1 filter=130 channel=5
    -7, -10, 8, 2, -7, 0, -2, 1, -8,
    -- layer=1 filter=130 channel=6
    3, -2, -3, -6, -1, -12, 4, 1, 0,
    -- layer=1 filter=130 channel=7
    0, 0, -2, 2, 10, 1, -4, -8, 7,
    -- layer=1 filter=130 channel=8
    0, 2, -11, 7, 1, -10, 3, -3, 8,
    -- layer=1 filter=130 channel=9
    4, 0, -2, -11, -4, 1, 2, -6, -1,
    -- layer=1 filter=130 channel=10
    6, -9, 1, -6, 10, 4, -7, -2, -1,
    -- layer=1 filter=130 channel=11
    7, -2, -3, -4, -7, 5, -3, 7, -4,
    -- layer=1 filter=130 channel=12
    -9, -9, 9, 7, -5, -7, -9, -9, 1,
    -- layer=1 filter=130 channel=13
    0, 3, -11, -6, 1, 2, 6, -7, 3,
    -- layer=1 filter=130 channel=14
    -5, 1, 9, -8, -5, -7, 9, 8, -10,
    -- layer=1 filter=130 channel=15
    3, -8, 4, -2, -2, -11, -12, 8, 3,
    -- layer=1 filter=130 channel=16
    -2, -4, -6, -9, 6, 0, -6, -4, 2,
    -- layer=1 filter=130 channel=17
    -6, 9, -11, 7, -7, 0, -12, 6, 6,
    -- layer=1 filter=130 channel=18
    -2, 4, 8, 1, 7, 0, 6, 5, -3,
    -- layer=1 filter=130 channel=19
    8, -1, 1, 3, -4, 2, 4, 7, 8,
    -- layer=1 filter=130 channel=20
    8, -5, -7, -9, -11, -11, 1, -3, -8,
    -- layer=1 filter=130 channel=21
    -9, 8, 3, 0, -5, 4, -9, -5, 6,
    -- layer=1 filter=130 channel=22
    -9, 6, -5, 4, 5, 3, 4, 7, -9,
    -- layer=1 filter=130 channel=23
    2, -5, -2, -7, -5, 7, 7, 4, -10,
    -- layer=1 filter=130 channel=24
    2, -1, 7, -8, 1, 3, -3, -8, 8,
    -- layer=1 filter=130 channel=25
    8, 10, 6, -1, 6, -4, 5, -10, 0,
    -- layer=1 filter=130 channel=26
    8, -6, 6, 8, -2, 8, -10, -3, 0,
    -- layer=1 filter=130 channel=27
    -8, 6, 6, 9, 8, -4, -3, 3, -8,
    -- layer=1 filter=130 channel=28
    -9, 7, -1, 5, 4, -6, -9, -2, -7,
    -- layer=1 filter=130 channel=29
    10, 1, -10, -6, -6, -11, -8, -1, -3,
    -- layer=1 filter=130 channel=30
    -9, -3, 10, -2, 0, 0, 6, -9, 7,
    -- layer=1 filter=130 channel=31
    -2, 10, 5, -1, 0, -10, 8, -3, 4,
    -- layer=1 filter=130 channel=32
    4, 8, -2, 1, -3, -9, 9, -9, -11,
    -- layer=1 filter=130 channel=33
    -2, 3, -9, -3, -7, 3, 3, 1, 7,
    -- layer=1 filter=130 channel=34
    -11, 4, 7, 0, 7, -12, -1, -5, -8,
    -- layer=1 filter=130 channel=35
    -3, -8, 5, -3, -9, -4, 7, 6, -10,
    -- layer=1 filter=130 channel=36
    5, 5, 0, 8, -12, -6, -7, -5, 7,
    -- layer=1 filter=130 channel=37
    10, 1, 0, 2, 3, 0, -5, -9, 3,
    -- layer=1 filter=130 channel=38
    0, 0, -8, -1, -4, -10, 2, -2, -3,
    -- layer=1 filter=130 channel=39
    1, -7, -2, -2, 3, 2, 0, -11, 3,
    -- layer=1 filter=130 channel=40
    0, -9, -9, -9, -4, -10, -10, -2, -5,
    -- layer=1 filter=130 channel=41
    -9, -9, 1, -12, 5, -6, -9, -4, 3,
    -- layer=1 filter=130 channel=42
    -5, 0, -5, 1, 1, -9, -7, 4, 6,
    -- layer=1 filter=130 channel=43
    -6, 3, -5, -2, -10, 2, -2, -8, 0,
    -- layer=1 filter=130 channel=44
    -10, -1, -4, -2, -10, -10, 3, -9, 1,
    -- layer=1 filter=130 channel=45
    1, -1, -10, -11, -3, 7, 0, 5, -5,
    -- layer=1 filter=130 channel=46
    -9, 0, -9, -1, -5, 3, 9, -9, -6,
    -- layer=1 filter=130 channel=47
    0, 0, 0, 6, 7, -2, 0, 4, -5,
    -- layer=1 filter=130 channel=48
    5, 4, -6, 2, 0, 3, 2, 8, 4,
    -- layer=1 filter=130 channel=49
    -3, -3, -9, 7, 0, 1, -2, -6, -6,
    -- layer=1 filter=130 channel=50
    -11, 0, 0, -4, -3, 2, 8, 7, 7,
    -- layer=1 filter=130 channel=51
    4, 7, 7, -8, -4, -1, -5, -10, 7,
    -- layer=1 filter=130 channel=52
    -7, -2, -3, 1, 1, 1, 0, 8, -8,
    -- layer=1 filter=130 channel=53
    -1, 9, 0, 4, -8, 0, -9, 3, 5,
    -- layer=1 filter=130 channel=54
    8, -8, 9, 2, -3, 6, 0, -8, -11,
    -- layer=1 filter=130 channel=55
    -5, -1, 5, 0, -10, -7, 8, 4, -9,
    -- layer=1 filter=130 channel=56
    7, -3, 5, -4, 9, 4, -6, -4, 8,
    -- layer=1 filter=130 channel=57
    6, -6, -6, 0, -3, 5, -1, 4, 8,
    -- layer=1 filter=130 channel=58
    9, 0, -6, -4, 0, 5, 2, -9, -11,
    -- layer=1 filter=130 channel=59
    -3, -9, -6, -6, 4, -11, 6, 5, 0,
    -- layer=1 filter=130 channel=60
    2, -9, -2, -8, -3, 2, -2, 0, 4,
    -- layer=1 filter=130 channel=61
    -4, 2, -9, 2, 5, 7, -6, 1, 0,
    -- layer=1 filter=130 channel=62
    6, -7, 0, -3, -1, -2, -7, 3, 1,
    -- layer=1 filter=130 channel=63
    -9, 0, -1, 7, -1, -7, -6, -11, 1,
    -- layer=1 filter=130 channel=64
    -7, -1, -9, 3, -2, -1, 0, 3, -7,
    -- layer=1 filter=130 channel=65
    -8, 3, 7, -8, -8, 2, 5, -6, 3,
    -- layer=1 filter=130 channel=66
    4, 2, -2, -2, 8, -4, -8, -9, -1,
    -- layer=1 filter=130 channel=67
    -1, -6, 5, -11, -4, 2, 0, 3, 10,
    -- layer=1 filter=130 channel=68
    -8, -9, 11, -2, -6, -4, 5, 5, -2,
    -- layer=1 filter=130 channel=69
    -8, 5, 0, 9, -1, 8, -1, -8, 10,
    -- layer=1 filter=130 channel=70
    -3, -5, -7, 2, -4, -5, -6, 0, -3,
    -- layer=1 filter=130 channel=71
    -2, -5, 1, -2, -10, -10, -3, -10, -4,
    -- layer=1 filter=130 channel=72
    -6, -1, 6, -2, -10, 5, -7, 2, -12,
    -- layer=1 filter=130 channel=73
    -9, -9, 2, -3, 5, 7, -3, -10, 5,
    -- layer=1 filter=130 channel=74
    3, 2, -7, -10, -4, -1, -1, 2, -11,
    -- layer=1 filter=130 channel=75
    -5, 1, -8, 6, -8, -4, 5, 1, -2,
    -- layer=1 filter=130 channel=76
    -2, -7, 5, 1, -6, 0, -2, -11, -7,
    -- layer=1 filter=130 channel=77
    8, -11, 8, 0, -4, -5, 8, -10, -8,
    -- layer=1 filter=130 channel=78
    -4, -8, 0, -3, -2, -10, -9, -11, -10,
    -- layer=1 filter=130 channel=79
    3, -2, -10, -7, -7, -5, -1, -12, -10,
    -- layer=1 filter=130 channel=80
    5, -9, 1, -4, 0, 4, 0, -5, -2,
    -- layer=1 filter=130 channel=81
    -3, -11, -8, -3, 7, 1, 6, 8, -6,
    -- layer=1 filter=130 channel=82
    -6, -4, -5, -4, -4, 1, 0, 6, 0,
    -- layer=1 filter=130 channel=83
    7, -9, -2, 4, -1, -9, 4, -4, 1,
    -- layer=1 filter=130 channel=84
    -11, -1, 6, -8, -2, -2, -9, 0, 6,
    -- layer=1 filter=130 channel=85
    -1, -2, 4, -9, -3, 6, -10, -8, 4,
    -- layer=1 filter=130 channel=86
    6, 6, 4, -5, -6, 3, -9, -3, -7,
    -- layer=1 filter=130 channel=87
    -8, 5, -4, -7, 5, 7, 5, 3, -9,
    -- layer=1 filter=130 channel=88
    -9, -5, -4, 2, 2, -7, 4, -2, -11,
    -- layer=1 filter=130 channel=89
    -5, 6, -6, 4, -7, 4, -2, 4, 8,
    -- layer=1 filter=130 channel=90
    -10, -7, -6, -4, -6, 0, 5, -3, -5,
    -- layer=1 filter=130 channel=91
    -3, -7, -2, 7, 2, -3, 1, -11, 0,
    -- layer=1 filter=130 channel=92
    0, -12, -12, -5, -7, 0, 3, 2, 0,
    -- layer=1 filter=130 channel=93
    5, 1, 7, 7, 6, -4, -4, -4, 0,
    -- layer=1 filter=130 channel=94
    8, -4, -8, 8, -12, 4, 2, 0, 0,
    -- layer=1 filter=130 channel=95
    -4, 6, -8, 8, 0, 2, -1, 2, -6,
    -- layer=1 filter=130 channel=96
    2, 0, 2, -2, 3, -6, 0, -12, -11,
    -- layer=1 filter=130 channel=97
    -7, -5, 0, -7, 0, -11, -12, 0, -6,
    -- layer=1 filter=130 channel=98
    -1, 5, 6, 9, -4, -5, 1, 3, 2,
    -- layer=1 filter=130 channel=99
    -2, -10, 2, 2, -10, -8, 7, -10, -2,
    -- layer=1 filter=130 channel=100
    2, -4, -9, 5, -9, -4, -7, 3, 6,
    -- layer=1 filter=130 channel=101
    -6, 6, -9, 7, -2, -10, -9, -4, 1,
    -- layer=1 filter=130 channel=102
    -9, 2, -11, -7, -4, -6, 7, 6, 0,
    -- layer=1 filter=130 channel=103
    -4, -8, -1, -7, 6, -10, -8, 1, -11,
    -- layer=1 filter=130 channel=104
    4, -6, -11, -1, -7, 3, -5, -6, 3,
    -- layer=1 filter=130 channel=105
    6, 0, 5, 7, -10, -10, -1, -8, -3,
    -- layer=1 filter=130 channel=106
    2, -1, -9, -3, -9, -10, -1, -2, 7,
    -- layer=1 filter=130 channel=107
    -6, 4, -9, -7, -10, -10, -1, 4, -6,
    -- layer=1 filter=130 channel=108
    4, 9, -3, -1, 7, 0, -1, -1, 4,
    -- layer=1 filter=130 channel=109
    -6, -6, -1, 0, -8, -5, 5, 0, -10,
    -- layer=1 filter=130 channel=110
    6, -11, -10, -1, -9, 6, -2, -10, -11,
    -- layer=1 filter=130 channel=111
    6, 6, -2, 3, -8, 5, 0, -7, 2,
    -- layer=1 filter=130 channel=112
    5, 3, -4, 3, -8, -8, 0, 1, 0,
    -- layer=1 filter=130 channel=113
    -5, -6, 1, -5, 6, 6, -10, 5, -10,
    -- layer=1 filter=130 channel=114
    7, 2, 2, 0, 5, 8, 0, -5, -9,
    -- layer=1 filter=130 channel=115
    -4, -10, 0, 2, -2, 4, 0, -11, -4,
    -- layer=1 filter=130 channel=116
    2, 2, 6, 5, 4, -5, -2, -2, -10,
    -- layer=1 filter=130 channel=117
    7, -7, 7, 3, -7, -5, 0, 5, 8,
    -- layer=1 filter=130 channel=118
    -7, -6, -9, -6, 0, -4, 0, -9, -9,
    -- layer=1 filter=130 channel=119
    0, -6, -5, -4, 7, 9, -6, -1, -7,
    -- layer=1 filter=130 channel=120
    8, -4, -6, 2, 0, -3, -7, 1, 6,
    -- layer=1 filter=130 channel=121
    0, 2, 9, 5, -2, 0, -6, -5, -6,
    -- layer=1 filter=130 channel=122
    0, 8, 4, -1, -5, -5, -9, 9, -10,
    -- layer=1 filter=130 channel=123
    -9, -7, -6, -2, 1, 4, -12, -10, -12,
    -- layer=1 filter=130 channel=124
    6, 3, -11, 0, 5, 1, -1, -4, 0,
    -- layer=1 filter=130 channel=125
    10, 7, 1, -3, 0, -1, 1, -7, -7,
    -- layer=1 filter=130 channel=126
    -5, -9, 7, -8, -12, 0, -12, -9, 5,
    -- layer=1 filter=130 channel=127
    7, -2, -2, 8, 8, -6, 6, 6, -3,
    -- layer=1 filter=131 channel=0
    -10, 6, -10, -6, -12, 3, -2, -9, 3,
    -- layer=1 filter=131 channel=1
    -1, -2, 0, -9, 1, -10, -2, 2, 7,
    -- layer=1 filter=131 channel=2
    4, 7, -1, -6, -7, 3, 0, -11, -1,
    -- layer=1 filter=131 channel=3
    9, -4, -7, -9, 7, 9, 0, 3, 3,
    -- layer=1 filter=131 channel=4
    6, 0, -11, -1, -6, -4, -3, -7, 7,
    -- layer=1 filter=131 channel=5
    -10, 10, -9, 5, 5, 0, -1, 6, 0,
    -- layer=1 filter=131 channel=6
    5, -7, -6, 6, 0, -10, -3, 0, 0,
    -- layer=1 filter=131 channel=7
    7, -9, 5, 9, -1, -6, -10, -6, 8,
    -- layer=1 filter=131 channel=8
    1, 7, -1, 0, -7, 4, -1, -1, -6,
    -- layer=1 filter=131 channel=9
    3, -3, -5, 0, 1, 5, -5, 2, 8,
    -- layer=1 filter=131 channel=10
    -2, -6, 4, -6, 6, 9, 4, 0, -2,
    -- layer=1 filter=131 channel=11
    -7, -9, -10, 1, -4, -8, 6, 5, -10,
    -- layer=1 filter=131 channel=12
    0, 9, 1, -10, 0, -4, 4, -2, -4,
    -- layer=1 filter=131 channel=13
    2, 2, 9, 5, 9, -2, -2, 5, 5,
    -- layer=1 filter=131 channel=14
    0, -2, 3, 8, 4, 4, -4, -4, 10,
    -- layer=1 filter=131 channel=15
    -10, 5, -10, 0, 6, -8, -8, 2, -5,
    -- layer=1 filter=131 channel=16
    -8, -3, 4, 2, 8, 5, 5, 3, 8,
    -- layer=1 filter=131 channel=17
    -11, -5, 0, 4, -3, -11, 0, 2, -2,
    -- layer=1 filter=131 channel=18
    -10, -10, -1, -10, 6, -3, 8, 0, -1,
    -- layer=1 filter=131 channel=19
    3, 8, -9, -8, 8, -1, 1, 8, 7,
    -- layer=1 filter=131 channel=20
    0, 7, 6, 5, 4, -7, -3, -4, -11,
    -- layer=1 filter=131 channel=21
    -7, -3, -5, -3, 6, -9, -9, 0, -1,
    -- layer=1 filter=131 channel=22
    0, 0, 5, 4, -10, 3, -1, -11, -9,
    -- layer=1 filter=131 channel=23
    4, -8, -11, -10, -6, 2, 7, 8, 7,
    -- layer=1 filter=131 channel=24
    7, 4, -5, -1, -10, 8, -7, -8, -5,
    -- layer=1 filter=131 channel=25
    1, 3, -5, -4, 3, -10, 1, -9, -9,
    -- layer=1 filter=131 channel=26
    -4, -8, 0, 1, 6, -1, 4, -11, 7,
    -- layer=1 filter=131 channel=27
    -10, -1, 5, -12, -3, -10, -1, -12, 0,
    -- layer=1 filter=131 channel=28
    -9, -11, 1, -10, 3, -6, 4, 4, 3,
    -- layer=1 filter=131 channel=29
    6, -6, -5, -7, -1, 1, -5, -10, 11,
    -- layer=1 filter=131 channel=30
    5, 8, -8, 1, -1, -11, -3, 1, 2,
    -- layer=1 filter=131 channel=31
    0, 4, -11, 0, -10, 5, -2, -7, -3,
    -- layer=1 filter=131 channel=32
    3, 0, -8, 7, 3, -9, -6, -8, -10,
    -- layer=1 filter=131 channel=33
    0, 0, -4, 8, -1, 7, 7, 10, 8,
    -- layer=1 filter=131 channel=34
    -11, -2, -4, 0, -1, -5, 1, -9, 0,
    -- layer=1 filter=131 channel=35
    3, 1, 0, 8, -6, -5, 2, -9, 8,
    -- layer=1 filter=131 channel=36
    7, -5, -4, 6, 7, 0, 5, -9, 0,
    -- layer=1 filter=131 channel=37
    -6, 9, 0, -6, 2, -6, 5, 1, -9,
    -- layer=1 filter=131 channel=38
    -5, 4, -9, -3, 1, 4, 7, -7, -5,
    -- layer=1 filter=131 channel=39
    -9, 5, -7, -4, -10, -7, -4, -7, -5,
    -- layer=1 filter=131 channel=40
    0, 3, 5, 3, 0, -7, 3, -2, -2,
    -- layer=1 filter=131 channel=41
    3, -4, -6, -9, 0, 6, -4, 9, -9,
    -- layer=1 filter=131 channel=42
    7, 7, 5, 0, 4, 5, 0, 2, 1,
    -- layer=1 filter=131 channel=43
    1, 0, 0, 0, 4, -11, -6, 3, -12,
    -- layer=1 filter=131 channel=44
    -6, 8, 4, 3, 0, -3, 8, 1, 7,
    -- layer=1 filter=131 channel=45
    -9, -2, 2, 0, 4, -6, 9, 6, 1,
    -- layer=1 filter=131 channel=46
    -2, -4, -3, 8, 3, -8, -1, -1, -6,
    -- layer=1 filter=131 channel=47
    1, 7, 5, 7, 0, 4, 4, 2, 5,
    -- layer=1 filter=131 channel=48
    4, -10, -1, -6, 4, -4, -9, -10, -2,
    -- layer=1 filter=131 channel=49
    1, 9, -6, 3, -9, 3, 8, 8, -6,
    -- layer=1 filter=131 channel=50
    -5, 2, -5, -12, 8, -1, -3, -6, -5,
    -- layer=1 filter=131 channel=51
    -4, 8, 7, -7, -10, 8, -5, -1, -4,
    -- layer=1 filter=131 channel=52
    -2, -1, -2, 0, -6, 9, -4, -6, 1,
    -- layer=1 filter=131 channel=53
    1, 5, -9, 5, 8, 7, 5, 5, 4,
    -- layer=1 filter=131 channel=54
    -2, -6, -7, 0, -8, -5, -9, -1, -5,
    -- layer=1 filter=131 channel=55
    -10, 5, 3, 2, 5, -11, -9, 3, 3,
    -- layer=1 filter=131 channel=56
    -8, 1, 7, -6, 0, 1, -8, -9, 2,
    -- layer=1 filter=131 channel=57
    7, 1, -8, -5, 8, -3, -10, 0, 1,
    -- layer=1 filter=131 channel=58
    -4, -9, 6, -7, 0, 0, 3, 0, -8,
    -- layer=1 filter=131 channel=59
    -8, -5, -2, -9, 5, -1, -3, 1, -11,
    -- layer=1 filter=131 channel=60
    6, -8, 2, 4, 4, 9, -9, 0, 0,
    -- layer=1 filter=131 channel=61
    2, -9, 7, 6, -2, -7, 0, -5, -10,
    -- layer=1 filter=131 channel=62
    -4, -1, 3, -3, 7, -4, -10, 6, 0,
    -- layer=1 filter=131 channel=63
    -7, 0, 0, -12, 4, 8, -10, 6, 4,
    -- layer=1 filter=131 channel=64
    7, 7, 1, -3, -7, -10, 0, -2, -11,
    -- layer=1 filter=131 channel=65
    -1, -10, 4, -5, -11, -2, -7, 7, 8,
    -- layer=1 filter=131 channel=66
    6, 7, 5, -1, 3, 1, -9, -5, -2,
    -- layer=1 filter=131 channel=67
    4, -9, -10, 0, 10, 0, 7, -1, -7,
    -- layer=1 filter=131 channel=68
    -8, -1, 1, 1, -2, 8, 4, 5, 4,
    -- layer=1 filter=131 channel=69
    4, -6, -5, -7, 1, -3, 8, 4, 6,
    -- layer=1 filter=131 channel=70
    0, -2, -10, 0, -4, 4, -7, 1, 0,
    -- layer=1 filter=131 channel=71
    1, 0, 7, -5, -8, -3, 6, -5, -8,
    -- layer=1 filter=131 channel=72
    -7, -1, -6, -1, -1, 5, -4, -7, 2,
    -- layer=1 filter=131 channel=73
    -6, -8, 0, -7, 0, -5, 4, -7, 0,
    -- layer=1 filter=131 channel=74
    6, -8, 8, 0, 0, 1, -4, -6, -1,
    -- layer=1 filter=131 channel=75
    -7, 8, 4, 0, -7, -9, -7, -4, -9,
    -- layer=1 filter=131 channel=76
    -2, -8, 0, 7, 5, -1, -2, 4, 0,
    -- layer=1 filter=131 channel=77
    -1, -12, -7, 4, 0, 7, 0, 8, -6,
    -- layer=1 filter=131 channel=78
    -7, -6, -9, -7, 5, 4, -6, 8, 6,
    -- layer=1 filter=131 channel=79
    1, -6, 0, -1, 1, -6, -1, -8, -3,
    -- layer=1 filter=131 channel=80
    -3, 0, -3, 9, -7, -5, -1, -5, -3,
    -- layer=1 filter=131 channel=81
    -10, 4, -2, 6, -5, 3, 0, 8, -5,
    -- layer=1 filter=131 channel=82
    2, -5, 8, -1, -4, 7, 6, 0, 1,
    -- layer=1 filter=131 channel=83
    2, 6, -5, -11, 0, 3, -1, -1, 8,
    -- layer=1 filter=131 channel=84
    6, -7, -10, -2, -2, 2, -5, -11, -4,
    -- layer=1 filter=131 channel=85
    0, 0, 3, 0, 1, 1, 8, 3, -3,
    -- layer=1 filter=131 channel=86
    -12, 1, -2, 5, 9, -10, -11, -11, 7,
    -- layer=1 filter=131 channel=87
    7, -10, 0, -8, 5, 0, -8, -1, -11,
    -- layer=1 filter=131 channel=88
    -2, -5, 1, 5, -7, -10, 4, -6, -9,
    -- layer=1 filter=131 channel=89
    3, 3, -6, -5, -9, 8, -9, -5, -9,
    -- layer=1 filter=131 channel=90
    -9, -9, 7, 6, 4, 9, -7, 5, -3,
    -- layer=1 filter=131 channel=91
    6, -10, -8, -9, 0, -4, 0, -6, -10,
    -- layer=1 filter=131 channel=92
    -10, 3, -1, -6, 0, -5, 9, -9, -7,
    -- layer=1 filter=131 channel=93
    -9, -2, 0, 1, -6, 3, -8, 7, -9,
    -- layer=1 filter=131 channel=94
    -4, -10, -9, -8, -1, 2, 6, -3, -1,
    -- layer=1 filter=131 channel=95
    -10, 0, -5, 9, -6, -2, 6, 5, -7,
    -- layer=1 filter=131 channel=96
    -4, 9, -8, 0, -4, -10, -10, 2, -8,
    -- layer=1 filter=131 channel=97
    6, -6, -11, 3, -9, -2, -7, -4, 3,
    -- layer=1 filter=131 channel=98
    -7, 0, 8, 0, 1, -3, 7, -10, 5,
    -- layer=1 filter=131 channel=99
    0, -10, -9, 5, 8, 2, -8, -1, 4,
    -- layer=1 filter=131 channel=100
    7, -2, 1, 1, 3, 5, 8, 0, 1,
    -- layer=1 filter=131 channel=101
    6, 4, -1, -11, -9, -12, -5, 0, -3,
    -- layer=1 filter=131 channel=102
    2, 0, 3, 3, -11, -3, -8, -11, -11,
    -- layer=1 filter=131 channel=103
    8, 1, 2, -8, 6, -3, 0, 5, -10,
    -- layer=1 filter=131 channel=104
    -4, 0, 7, -9, 0, 2, 6, -4, 3,
    -- layer=1 filter=131 channel=105
    2, -1, 6, 1, -5, -1, -10, 0, 4,
    -- layer=1 filter=131 channel=106
    -4, 1, 0, -1, -9, 1, -3, -5, 3,
    -- layer=1 filter=131 channel=107
    7, 4, -6, -10, 8, -1, 0, 8, 8,
    -- layer=1 filter=131 channel=108
    5, 8, 1, 4, -4, -2, -2, -8, -3,
    -- layer=1 filter=131 channel=109
    0, 4, -5, -10, -4, -9, 2, 3, 4,
    -- layer=1 filter=131 channel=110
    -3, -11, 1, 8, 7, 0, 5, 4, -2,
    -- layer=1 filter=131 channel=111
    0, -2, -8, 4, -6, 0, 2, 8, 8,
    -- layer=1 filter=131 channel=112
    -6, -3, -2, -2, 6, -1, -4, 0, 7,
    -- layer=1 filter=131 channel=113
    4, 9, -3, 5, -4, -5, 5, 3, 0,
    -- layer=1 filter=131 channel=114
    -6, -5, 7, -4, -7, 0, -4, -2, 7,
    -- layer=1 filter=131 channel=115
    0, 8, 5, 0, 0, -8, -1, -10, 0,
    -- layer=1 filter=131 channel=116
    3, 9, 9, -9, 7, 7, 1, -2, -3,
    -- layer=1 filter=131 channel=117
    -8, -1, 1, -1, 8, 5, -6, -8, -9,
    -- layer=1 filter=131 channel=118
    -10, -6, -4, -7, 3, -6, -9, -7, 2,
    -- layer=1 filter=131 channel=119
    -6, -5, 0, -3, 1, 3, -4, 6, 7,
    -- layer=1 filter=131 channel=120
    -2, 6, -4, -9, 5, -10, -10, -10, -7,
    -- layer=1 filter=131 channel=121
    2, 0, 6, 2, 4, -12, 4, -7, 5,
    -- layer=1 filter=131 channel=122
    2, -2, 9, -1, -4, 2, 6, 8, -10,
    -- layer=1 filter=131 channel=123
    5, -11, 8, 0, -2, -9, 7, -8, 6,
    -- layer=1 filter=131 channel=124
    -7, 5, -7, -1, 5, 5, 0, -7, 0,
    -- layer=1 filter=131 channel=125
    -3, 8, 0, 8, 10, -7, -10, -5, -5,
    -- layer=1 filter=131 channel=126
    6, 0, 7, 7, -3, -10, -7, 0, -3,
    -- layer=1 filter=131 channel=127
    6, -3, -6, 9, -6, 0, -10, -7, -2,
    -- layer=1 filter=132 channel=0
    6, 1, -3, 14, -8, -8, -15, -30, -11,
    -- layer=1 filter=132 channel=1
    -3, 15, 5, 18, 19, 29, -46, -24, -43,
    -- layer=1 filter=132 channel=2
    25, 4, 23, 12, 32, 35, 27, 38, 12,
    -- layer=1 filter=132 channel=3
    -6, 1, 6, 4, 6, -8, 8, 1, -2,
    -- layer=1 filter=132 channel=4
    2, -5, 6, -3, 8, -14, 21, 21, 17,
    -- layer=1 filter=132 channel=5
    4, 11, -22, 37, 25, 26, -37, -8, -23,
    -- layer=1 filter=132 channel=6
    37, 44, 8, 18, 18, -20, 9, -18, -37,
    -- layer=1 filter=132 channel=7
    8, -16, -36, -7, -68, -44, -77, -37, -30,
    -- layer=1 filter=132 channel=8
    4, 3, -2, 35, 30, 31, -27, 22, -5,
    -- layer=1 filter=132 channel=9
    -26, 7, 83, 10, 18, 59, 28, 58, -27,
    -- layer=1 filter=132 channel=10
    15, -18, -26, -11, -37, -41, -56, -43, -19,
    -- layer=1 filter=132 channel=11
    -17, 0, 9, 0, 8, 2, -16, -26, -13,
    -- layer=1 filter=132 channel=12
    7, 38, 0, 18, 42, 6, 45, 2, -19,
    -- layer=1 filter=132 channel=13
    18, 29, 17, 0, 8, -7, -12, -27, -29,
    -- layer=1 filter=132 channel=14
    3, -12, -33, 32, -5, -31, -1, -22, -32,
    -- layer=1 filter=132 channel=15
    19, 20, -36, 33, 10, -18, -22, -26, -8,
    -- layer=1 filter=132 channel=16
    0, 19, 1, 33, 48, 26, -13, 19, 18,
    -- layer=1 filter=132 channel=17
    8, 16, 11, -11, -7, -15, -46, -31, -27,
    -- layer=1 filter=132 channel=18
    0, -10, 14, 32, 47, 31, 29, -3, -20,
    -- layer=1 filter=132 channel=19
    24, 25, 45, 116, 73, 83, 49, 32, 23,
    -- layer=1 filter=132 channel=20
    21, 27, 7, 20, 1, -2, -15, 0, -13,
    -- layer=1 filter=132 channel=21
    6, 12, 11, -3, -10, -34, -34, -40, -29,
    -- layer=1 filter=132 channel=22
    27, 51, 20, 24, 37, 22, -23, -13, -29,
    -- layer=1 filter=132 channel=23
    35, 37, -19, -9, -57, -52, -70, -68, -75,
    -- layer=1 filter=132 channel=24
    3, -2, 0, 8, -6, 28, -6, -12, -11,
    -- layer=1 filter=132 channel=25
    42, 48, 22, 7, 35, 16, -43, 31, 8,
    -- layer=1 filter=132 channel=26
    0, 22, 24, 0, 10, 5, 1, -34, -27,
    -- layer=1 filter=132 channel=27
    -23, -22, -15, -16, -18, -3, 6, 18, 20,
    -- layer=1 filter=132 channel=28
    43, 8, 8, -19, -20, -27, -75, -8, -16,
    -- layer=1 filter=132 channel=29
    -24, -11, 25, -7, 0, 4, 1, 0, -6,
    -- layer=1 filter=132 channel=30
    -22, -35, -7, 28, 45, 29, 43, 32, -26,
    -- layer=1 filter=132 channel=31
    24, 25, 24, 24, 36, 37, 3, -12, -24,
    -- layer=1 filter=132 channel=32
    -13, 7, 36, -18, 31, 13, -6, -28, -87,
    -- layer=1 filter=132 channel=33
    23, 26, 4, 4, 34, 19, -5, -7, -13,
    -- layer=1 filter=132 channel=34
    23, 7, 0, -1, -2, -29, -10, -30, -47,
    -- layer=1 filter=132 channel=35
    -15, -22, -19, -15, -10, -28, -12, -12, -31,
    -- layer=1 filter=132 channel=36
    -9, -16, 1, 0, 6, 5, 0, -3, -16,
    -- layer=1 filter=132 channel=37
    4, 24, 0, 43, 63, 53, -17, 0, 1,
    -- layer=1 filter=132 channel=38
    28, 24, 6, 6, 7, -14, -10, -20, -31,
    -- layer=1 filter=132 channel=39
    14, 14, 9, -14, -16, -18, -19, -7, -4,
    -- layer=1 filter=132 channel=40
    36, 27, 18, 25, 30, 0, -5, -29, -51,
    -- layer=1 filter=132 channel=41
    -33, -15, 50, 23, 51, 66, 5, 19, -64,
    -- layer=1 filter=132 channel=42
    21, 32, 16, 28, 31, 33, 40, 13, 30,
    -- layer=1 filter=132 channel=43
    10, 29, -11, 11, 35, 24, -22, 6, 0,
    -- layer=1 filter=132 channel=44
    -20, 13, 18, -18, -10, -33, -19, -76, -121,
    -- layer=1 filter=132 channel=45
    11, 16, -26, 14, 6, -7, -19, -24, -18,
    -- layer=1 filter=132 channel=46
    32, 19, -25, 102, 79, 40, 15, -7, -32,
    -- layer=1 filter=132 channel=47
    6, 28, 19, -7, 18, -8, -38, -17, -62,
    -- layer=1 filter=132 channel=48
    10, 7, -11, -8, -20, -58, -15, -47, -47,
    -- layer=1 filter=132 channel=49
    36, 36, 39, 17, 25, 7, -5, -3, -50,
    -- layer=1 filter=132 channel=50
    25, -5, 12, -9, -1, 26, -7, 7, -6,
    -- layer=1 filter=132 channel=51
    32, 16, -6, 14, -30, -38, -33, -32, -26,
    -- layer=1 filter=132 channel=52
    18, 23, 15, 8, 15, 16, 16, 25, 16,
    -- layer=1 filter=132 channel=53
    -2, 10, -3, 12, 5, -1, 18, 11, 21,
    -- layer=1 filter=132 channel=54
    30, 36, 36, 11, 40, 46, -24, 12, 20,
    -- layer=1 filter=132 channel=55
    3, 0, 0, -3, 15, 17, 0, 0, 21,
    -- layer=1 filter=132 channel=56
    -11, 9, -11, 8, -6, 1, -9, -16, 3,
    -- layer=1 filter=132 channel=57
    48, 29, 1, -1, -5, -15, -30, -19, 0,
    -- layer=1 filter=132 channel=58
    27, -2, 9, -31, -45, -24, -100, -71, -42,
    -- layer=1 filter=132 channel=59
    4, -3, -32, -17, -44, -36, 6, -5, 0,
    -- layer=1 filter=132 channel=60
    0, 8, 1, 24, 14, -2, 16, -2, -9,
    -- layer=1 filter=132 channel=61
    -5, 1, 5, -5, -4, 5, -7, 2, -9,
    -- layer=1 filter=132 channel=62
    16, 13, -13, 13, 38, 17, -14, -7, 5,
    -- layer=1 filter=132 channel=63
    -21, 0, -6, -1, 35, 10, 2, -15, 0,
    -- layer=1 filter=132 channel=64
    0, 18, -4, 5, 7, -9, -43, -32, -51,
    -- layer=1 filter=132 channel=65
    15, 5, -26, 9, -50, -67, -35, -27, -36,
    -- layer=1 filter=132 channel=66
    -1, 4, -10, 5, -2, -4, -8, -16, -4,
    -- layer=1 filter=132 channel=67
    61, 64, 42, -1, -27, -56, 12, -53, -65,
    -- layer=1 filter=132 channel=68
    -15, 12, 22, -39, 18, -26, -30, -98, -119,
    -- layer=1 filter=132 channel=69
    6, 15, -36, 38, 12, 11, -4, -3, -13,
    -- layer=1 filter=132 channel=70
    35, 34, 11, 24, 35, 6, 11, -12, -45,
    -- layer=1 filter=132 channel=71
    5, 0, -23, -2, -6, -6, -11, -15, -11,
    -- layer=1 filter=132 channel=72
    -16, -32, 3, 54, 56, 45, 60, 42, 12,
    -- layer=1 filter=132 channel=73
    -7, 0, -3, 2, -16, 5, 0, -2, -16,
    -- layer=1 filter=132 channel=74
    1, 15, 41, 7, 57, 16, 5, -30, -61,
    -- layer=1 filter=132 channel=75
    -13, -15, -28, 42, 33, 0, 42, 9, 2,
    -- layer=1 filter=132 channel=76
    -35, -1, 21, -14, 41, 28, 15, -22, -40,
    -- layer=1 filter=132 channel=77
    4, 11, -17, -26, -46, -53, -45, -41, -31,
    -- layer=1 filter=132 channel=78
    -2, 21, 0, -13, 8, 2, -13, -11, -1,
    -- layer=1 filter=132 channel=79
    29, 27, 5, 30, 46, 32, -4, 2, -5,
    -- layer=1 filter=132 channel=80
    -2, -13, -12, 6, 2, -22, 7, 4, 14,
    -- layer=1 filter=132 channel=81
    3, -19, -24, -11, 2, -13, -17, -16, 21,
    -- layer=1 filter=132 channel=82
    17, 24, -4, -6, -20, -51, -12, -35, -53,
    -- layer=1 filter=132 channel=83
    -2, 12, -19, -4, -22, -22, -42, -59, -45,
    -- layer=1 filter=132 channel=84
    12, 15, 40, 13, 72, 41, 33, -12, -35,
    -- layer=1 filter=132 channel=85
    11, 29, 21, 5, 4, 7, -50, -26, -26,
    -- layer=1 filter=132 channel=86
    -5, -13, 0, 0, -1, 2, -7, 1, 4,
    -- layer=1 filter=132 channel=87
    -20, -4, 24, 86, 69, 91, 22, 60, 4,
    -- layer=1 filter=132 channel=88
    13, 9, -7, -4, -11, -32, -4, -35, -60,
    -- layer=1 filter=132 channel=89
    -3, 13, 6, -2, -27, -71, -21, -49, -79,
    -- layer=1 filter=132 channel=90
    -27, -5, -8, -30, -32, -43, -19, -60, -100,
    -- layer=1 filter=132 channel=91
    11, 24, 0, 3, 9, -5, 0, -14, -18,
    -- layer=1 filter=132 channel=92
    4, 0, -6, -7, 15, 17, -15, -16, -87,
    -- layer=1 filter=132 channel=93
    0, -8, -10, -14, -17, -23, -22, -22, -21,
    -- layer=1 filter=132 channel=94
    -24, -14, -20, -1, -2, -17, -34, -17, -25,
    -- layer=1 filter=132 channel=95
    0, 6, 32, 33, 62, 10, 36, 3, -28,
    -- layer=1 filter=132 channel=96
    -1, 5, 18, -25, 4, -10, -21, -44, -52,
    -- layer=1 filter=132 channel=97
    -14, 10, -3, -17, -30, -25, -18, -18, -2,
    -- layer=1 filter=132 channel=98
    30, 30, 14, 20, 30, 21, -15, 9, 20,
    -- layer=1 filter=132 channel=99
    47, 0, 21, -18, -38, -73, -86, -114, -84,
    -- layer=1 filter=132 channel=100
    -33, -22, -10, 7, 27, 6, 1, -7, -5,
    -- layer=1 filter=132 channel=101
    21, 31, 14, 16, 2, -28, -9, -29, -53,
    -- layer=1 filter=132 channel=102
    -12, -26, -15, -2, 19, 3, -32, -34, -28,
    -- layer=1 filter=132 channel=103
    -6, 1, 12, 4, 12, 23, -12, 5, -8,
    -- layer=1 filter=132 channel=104
    -2, -10, 17, 25, 11, 24, 0, 8, -27,
    -- layer=1 filter=132 channel=105
    -10, -9, -8, -4, -15, -20, -33, -26, -4,
    -- layer=1 filter=132 channel=106
    17, 30, 39, 0, 22, -19, -20, -46, -68,
    -- layer=1 filter=132 channel=107
    -29, -15, -21, 14, -4, 2, -16, 1, 7,
    -- layer=1 filter=132 channel=108
    -3, -10, -3, -12, -15, -26, 1, -37, -80,
    -- layer=1 filter=132 channel=109
    -10, -10, -5, -6, -8, -2, -8, -7, -9,
    -- layer=1 filter=132 channel=110
    -5, -3, -9, -7, -8, -14, -17, -24, -31,
    -- layer=1 filter=132 channel=111
    -21, -13, -6, 22, 50, -1, 35, -21, -60,
    -- layer=1 filter=132 channel=112
    14, 30, 61, 23, 72, 4, 12, -24, -39,
    -- layer=1 filter=132 channel=113
    67, 62, 33, 43, 33, 11, 7, -1, 0,
    -- layer=1 filter=132 channel=114
    -4, -7, -42, 18, 22, 25, -5, 5, 14,
    -- layer=1 filter=132 channel=115
    -2, -9, -11, -4, -30, -21, -34, -20, -8,
    -- layer=1 filter=132 channel=116
    -4, -2, -4, 8, -5, -3, 7, 6, 4,
    -- layer=1 filter=132 channel=117
    57, 47, 62, 61, 56, -2, 22, -38, -41,
    -- layer=1 filter=132 channel=118
    -15, -2, 25, 10, 56, 15, 26, 12, -22,
    -- layer=1 filter=132 channel=119
    -24, -2, 23, -21, 12, -14, -21, -55, -106,
    -- layer=1 filter=132 channel=120
    21, 32, -1, 16, 17, -13, -15, 7, 0,
    -- layer=1 filter=132 channel=121
    5, -23, -26, 62, 35, 56, 33, 41, -10,
    -- layer=1 filter=132 channel=122
    -8, -9, 4, 1, -3, -3, -6, 7, 0,
    -- layer=1 filter=132 channel=123
    3, -27, -24, 40, 32, 39, 8, 14, 4,
    -- layer=1 filter=132 channel=124
    -16, -23, -27, -20, -10, -15, -14, -5, -29,
    -- layer=1 filter=132 channel=125
    40, 52, 35, 40, 39, 11, -10, -15, -50,
    -- layer=1 filter=132 channel=126
    9, 32, -3, 19, 20, 7, -37, -12, -33,
    -- layer=1 filter=132 channel=127
    -22, 3, 3, 17, 63, 26, 51, 26, -22,
    -- layer=1 filter=133 channel=0
    -2, 5, -3, -6, 1, -17, 1, -22, -17,
    -- layer=1 filter=133 channel=1
    20, 8, -7, 16, -18, -6, -33, -40, 0,
    -- layer=1 filter=133 channel=2
    22, -29, 18, 25, 8, 48, 6, 6, 22,
    -- layer=1 filter=133 channel=3
    9, -10, 7, -8, 0, -9, 0, -10, 4,
    -- layer=1 filter=133 channel=4
    0, -6, 12, 0, 0, 2, -6, 7, 4,
    -- layer=1 filter=133 channel=5
    25, 0, -19, 15, -61, -35, -42, -33, 14,
    -- layer=1 filter=133 channel=6
    -2, 19, 13, -13, 12, -5, 31, 18, -24,
    -- layer=1 filter=133 channel=7
    11, 21, -28, 26, -20, -41, 10, -9, 26,
    -- layer=1 filter=133 channel=8
    30, 12, -8, 11, -65, -51, -37, -16, 39,
    -- layer=1 filter=133 channel=9
    3, 5, 4, -8, 22, 36, 9, 38, -14,
    -- layer=1 filter=133 channel=10
    -4, 14, -35, 18, -29, -35, -16, -18, 25,
    -- layer=1 filter=133 channel=11
    -25, -29, -8, -10, 2, 15, 14, 21, 8,
    -- layer=1 filter=133 channel=12
    9, 4, 16, -67, -29, 1, -24, -21, 3,
    -- layer=1 filter=133 channel=13
    4, 12, 0, -7, 27, 4, 23, 16, -21,
    -- layer=1 filter=133 channel=14
    -6, -10, -11, -9, -27, -37, 8, -24, -7,
    -- layer=1 filter=133 channel=15
    10, -7, -27, -24, -76, -31, -20, -21, 2,
    -- layer=1 filter=133 channel=16
    11, 2, -35, 10, -52, -66, -40, 5, 52,
    -- layer=1 filter=133 channel=17
    -7, 11, 13, 0, -3, -17, -33, -25, -29,
    -- layer=1 filter=133 channel=18
    -16, -32, 22, -54, 15, 34, 30, 30, 10,
    -- layer=1 filter=133 channel=19
    64, 68, 15, 64, 29, 68, 41, 110, 73,
    -- layer=1 filter=133 channel=20
    17, 17, -2, 16, 16, -19, 7, -2, -9,
    -- layer=1 filter=133 channel=21
    18, 21, 0, 3, -7, -15, -13, -26, 15,
    -- layer=1 filter=133 channel=22
    19, 34, 10, 24, 8, -21, -12, -11, -12,
    -- layer=1 filter=133 channel=23
    65, 3, -25, 3, -58, 0, 0, 8, 1,
    -- layer=1 filter=133 channel=24
    16, -22, -10, -27, -17, -13, -9, 5, -13,
    -- layer=1 filter=133 channel=25
    30, 36, -12, 54, 9, -35, -9, 25, 61,
    -- layer=1 filter=133 channel=26
    -11, -12, -1, -20, 1, 11, 32, 46, -20,
    -- layer=1 filter=133 channel=27
    47, 28, 24, 15, 18, 12, -9, -24, -15,
    -- layer=1 filter=133 channel=28
    22, 49, -12, 12, -2, -54, -30, -54, 6,
    -- layer=1 filter=133 channel=29
    32, 16, 9, 4, -8, -15, -12, -42, -29,
    -- layer=1 filter=133 channel=30
    0, -4, 41, -37, -14, 52, 36, 55, 3,
    -- layer=1 filter=133 channel=31
    7, 7, 41, -23, 14, 21, 9, 13, 14,
    -- layer=1 filter=133 channel=32
    -18, -20, -15, -10, 21, 27, 35, 36, 6,
    -- layer=1 filter=133 channel=33
    1, 25, 7, -10, 13, 8, -15, 2, -26,
    -- layer=1 filter=133 channel=34
    2, 7, 11, -6, 6, -16, -2, 7, -3,
    -- layer=1 filter=133 channel=35
    -1, -13, -14, -13, -20, -14, -11, -17, -15,
    -- layer=1 filter=133 channel=36
    -30, -13, -6, -17, 6, 11, 1, 10, 2,
    -- layer=1 filter=133 channel=37
    28, 0, -13, 15, -17, -26, -50, 4, 50,
    -- layer=1 filter=133 channel=38
    15, 9, 0, -4, 14, -1, 3, 13, -9,
    -- layer=1 filter=133 channel=39
    -1, 3, -3, 8, -11, -14, -27, -15, -2,
    -- layer=1 filter=133 channel=40
    -4, -1, 15, -7, -9, 7, 15, 23, -8,
    -- layer=1 filter=133 channel=41
    9, -30, -21, 5, 45, 48, 55, 98, 0,
    -- layer=1 filter=133 channel=42
    21, -7, -4, 12, -13, 12, 8, -3, 21,
    -- layer=1 filter=133 channel=43
    25, 39, -21, 18, -23, -63, -23, 13, 57,
    -- layer=1 filter=133 channel=44
    -24, -8, -2, -7, 19, 4, 25, 28, -21,
    -- layer=1 filter=133 channel=45
    3, -4, -11, -21, -19, -16, -1, -11, -1,
    -- layer=1 filter=133 channel=46
    32, 37, 4, -19, -43, 9, -4, 32, 15,
    -- layer=1 filter=133 channel=47
    32, -20, -7, 27, -6, 38, 10, 32, 11,
    -- layer=1 filter=133 channel=48
    30, 16, 23, -1, -14, -1, 0, -14, -25,
    -- layer=1 filter=133 channel=49
    0, -1, -9, -15, 1, 2, -8, 5, -14,
    -- layer=1 filter=133 channel=50
    0, -15, -11, -6, -5, 14, -23, -9, -22,
    -- layer=1 filter=133 channel=51
    22, 14, 7, 8, -26, -19, -15, -36, 0,
    -- layer=1 filter=133 channel=52
    9, -11, -12, -15, -6, -6, 6, 15, 20,
    -- layer=1 filter=133 channel=53
    -13, -4, -12, -5, -19, -12, -5, 0, -4,
    -- layer=1 filter=133 channel=54
    35, 29, -10, 59, 7, -21, 1, 41, 89,
    -- layer=1 filter=133 channel=55
    2, -6, 12, 7, 1, 25, 7, 16, 9,
    -- layer=1 filter=133 channel=56
    -8, -2, -6, 12, 6, 11, -3, 5, 5,
    -- layer=1 filter=133 channel=57
    11, 11, -14, 25, -20, -25, -25, -11, 20,
    -- layer=1 filter=133 channel=58
    48, 12, -8, 45, -24, 26, 25, 46, 63,
    -- layer=1 filter=133 channel=59
    10, 0, 4, 3, 3, 4, -11, 6, -9,
    -- layer=1 filter=133 channel=60
    9, 15, 15, 2, 26, 17, 17, 9, 11,
    -- layer=1 filter=133 channel=61
    4, 6, -2, 1, -14, 0, 2, -2, 1,
    -- layer=1 filter=133 channel=62
    30, 5, -16, 16, -43, -65, -56, 3, 38,
    -- layer=1 filter=133 channel=63
    -9, -3, 1, -29, 15, 21, 3, 14, -18,
    -- layer=1 filter=133 channel=64
    23, 16, 5, 9, 5, -12, -7, -18, -10,
    -- layer=1 filter=133 channel=65
    9, 24, 8, 1, 2, -5, -14, -20, -10,
    -- layer=1 filter=133 channel=66
    -6, 5, 0, 5, -4, -8, -17, -26, -17,
    -- layer=1 filter=133 channel=67
    28, 15, 12, -2, -23, -38, -17, -32, -23,
    -- layer=1 filter=133 channel=68
    -25, -2, 11, -7, 41, 29, 51, 47, 3,
    -- layer=1 filter=133 channel=69
    -2, -30, -58, -25, -78, -28, -28, -10, 32,
    -- layer=1 filter=133 channel=70
    -17, -10, 5, -49, -29, -9, -16, -17, -33,
    -- layer=1 filter=133 channel=71
    38, 21, 0, 0, -37, -23, -40, -42, 13,
    -- layer=1 filter=133 channel=72
    18, 4, 15, 2, 26, 71, 30, 86, 37,
    -- layer=1 filter=133 channel=73
    -1, 9, -2, 3, -4, 9, -2, -10, 0,
    -- layer=1 filter=133 channel=74
    -16, -6, 27, -21, 51, 21, 48, 58, -4,
    -- layer=1 filter=133 channel=75
    -41, -14, 44, -76, -34, 5, 0, -17, 23,
    -- layer=1 filter=133 channel=76
    -34, -26, 5, -20, 28, 0, 35, 31, -20,
    -- layer=1 filter=133 channel=77
    18, 15, 10, 6, -18, -30, -23, -34, -5,
    -- layer=1 filter=133 channel=78
    6, 20, 5, 20, 12, -4, -17, 4, -9,
    -- layer=1 filter=133 channel=79
    27, 8, -35, 18, -54, -75, -39, 0, 29,
    -- layer=1 filter=133 channel=80
    12, 15, 3, 7, 0, 5, -5, 15, 19,
    -- layer=1 filter=133 channel=81
    30, 9, -2, -11, -50, -53, -43, -41, -2,
    -- layer=1 filter=133 channel=82
    25, 15, 7, 6, -16, -7, -17, -29, -21,
    -- layer=1 filter=133 channel=83
    14, 7, -11, -25, -18, -34, -34, -21, -26,
    -- layer=1 filter=133 channel=84
    -4, -11, 46, -28, 53, 55, 83, 58, 0,
    -- layer=1 filter=133 channel=85
    33, 6, -26, 28, -29, 11, 13, 45, 7,
    -- layer=1 filter=133 channel=86
    12, 20, 11, 6, 10, 9, -13, -5, 9,
    -- layer=1 filter=133 channel=87
    51, 48, -7, 35, 26, 68, 23, 98, 43,
    -- layer=1 filter=133 channel=88
    10, -12, 0, -9, -14, 1, -15, -1, -9,
    -- layer=1 filter=133 channel=89
    11, 8, 23, -2, 6, -12, 16, -20, -22,
    -- layer=1 filter=133 channel=90
    -36, -14, -3, -34, 2, 5, 7, 33, 0,
    -- layer=1 filter=133 channel=91
    15, 16, 23, 16, 10, 0, 7, -1, -3,
    -- layer=1 filter=133 channel=92
    -39, -11, -29, -60, 1, 7, 7, 7, 30,
    -- layer=1 filter=133 channel=93
    25, 8, 6, 14, -8, -22, -19, -40, -20,
    -- layer=1 filter=133 channel=94
    -18, 8, -6, -6, 9, -5, -11, -22, -27,
    -- layer=1 filter=133 channel=95
    -19, -14, 56, -30, 38, 35, 49, 43, 0,
    -- layer=1 filter=133 channel=96
    15, 22, 7, 3, 5, 1, 10, 17, -2,
    -- layer=1 filter=133 channel=97
    12, 21, 0, 7, 7, -22, -9, -25, -22,
    -- layer=1 filter=133 channel=98
    37, 11, -15, -5, -24, -69, -52, -23, 49,
    -- layer=1 filter=133 channel=99
    -14, 14, -4, -4, -19, -33, -41, -41, 5,
    -- layer=1 filter=133 channel=100
    -25, -12, 9, -36, 12, 3, 7, 27, -8,
    -- layer=1 filter=133 channel=101
    17, 16, 18, 1, 15, -10, 19, -6, -15,
    -- layer=1 filter=133 channel=102
    -6, 2, 14, 2, -3, -15, -5, -23, -54,
    -- layer=1 filter=133 channel=103
    -6, -3, 18, -22, 0, 21, 5, 11, 3,
    -- layer=1 filter=133 channel=104
    19, -10, -35, 5, -22, 13, 18, 29, 21,
    -- layer=1 filter=133 channel=105
    -9, 0, 9, 10, -4, -10, -18, -28, -24,
    -- layer=1 filter=133 channel=106
    -5, 11, 16, -7, 37, 14, 35, 15, -19,
    -- layer=1 filter=133 channel=107
    -13, -1, -18, -14, -19, -13, -6, -2, -4,
    -- layer=1 filter=133 channel=108
    -6, -35, -28, -11, -7, -11, 23, 22, -13,
    -- layer=1 filter=133 channel=109
    0, -4, 0, 1, 5, -5, 9, 7, 1,
    -- layer=1 filter=133 channel=110
    0, -4, -1, 11, 0, 0, -8, -15, -11,
    -- layer=1 filter=133 channel=111
    -17, -56, 48, -58, -3, 29, 25, 16, -26,
    -- layer=1 filter=133 channel=112
    -14, -19, 28, -29, 42, -3, 47, 5, 4,
    -- layer=1 filter=133 channel=113
    13, 7, 0, -15, -22, -2, -5, -18, -7,
    -- layer=1 filter=133 channel=114
    -21, -26, -38, -33, -68, -18, -26, -12, -3,
    -- layer=1 filter=133 channel=115
    15, 16, -4, 22, -19, -7, -7, -22, 8,
    -- layer=1 filter=133 channel=116
    4, 3, -3, -9, 1, 0, -9, 10, 0,
    -- layer=1 filter=133 channel=117
    -31, -56, 21, -17, 4, 13, 26, -34, -18,
    -- layer=1 filter=133 channel=118
    -17, -22, 45, -40, 17, 27, 42, 57, -7,
    -- layer=1 filter=133 channel=119
    -2, -13, 0, -19, 14, 33, 38, 48, 1,
    -- layer=1 filter=133 channel=120
    27, 1, -17, 8, -18, -36, -21, -14, 24,
    -- layer=1 filter=133 channel=121
    8, 8, 13, -24, -28, 37, -40, 6, 25,
    -- layer=1 filter=133 channel=122
    2, -2, -2, 8, -8, 9, 1, 10, 5,
    -- layer=1 filter=133 channel=123
    1, -9, -23, -25, -21, 13, -22, -7, 22,
    -- layer=1 filter=133 channel=124
    6, 11, 7, -10, -9, 0, -9, 5, -6,
    -- layer=1 filter=133 channel=125
    -11, -26, -16, -5, -39, -15, -32, -19, -14,
    -- layer=1 filter=133 channel=126
    36, 16, 3, -34, -30, -61, -84, -56, -3,
    -- layer=1 filter=133 channel=127
    -12, -10, 41, -43, 35, 42, 66, 45, 15,
    -- layer=1 filter=134 channel=0
    6, -31, -31, 2, -44, -25, 15, -39, -18,
    -- layer=1 filter=134 channel=1
    50, 46, -61, -20, -58, 15, -52, -36, 23,
    -- layer=1 filter=134 channel=2
    -62, -62, 16, 12, 28, 34, 24, 27, -19,
    -- layer=1 filter=134 channel=3
    5, 3, -1, 1, -1, 0, 4, -4, -2,
    -- layer=1 filter=134 channel=4
    -14, -7, -15, -7, 4, -13, 0, -7, -14,
    -- layer=1 filter=134 channel=5
    39, -10, -52, -58, -56, 5, -45, -12, 31,
    -- layer=1 filter=134 channel=6
    12, 44, 39, 33, -11, -30, -11, -42, -14,
    -- layer=1 filter=134 channel=7
    -45, -85, -60, -125, -42, 37, -100, 40, 54,
    -- layer=1 filter=134 channel=8
    102, 19, -43, -46, -26, 25, -51, -11, 37,
    -- layer=1 filter=134 channel=9
    33, 45, 101, 21, 114, 5, 40, 8, -16,
    -- layer=1 filter=134 channel=10
    -69, -94, -32, -144, -43, 45, -86, 43, 56,
    -- layer=1 filter=134 channel=11
    13, -14, -36, 13, -21, -30, -3, -36, -18,
    -- layer=1 filter=134 channel=12
    76, 69, 53, 33, -30, -42, 24, 23, -39,
    -- layer=1 filter=134 channel=13
    -5, 16, 28, 20, 23, -11, 17, -31, -40,
    -- layer=1 filter=134 channel=14
    -25, -38, -57, -52, -61, -24, -58, -6, 2,
    -- layer=1 filter=134 channel=15
    -65, -51, -62, -74, -26, -28, -33, -16, -35,
    -- layer=1 filter=134 channel=16
    69, -14, -34, -79, -32, 28, -42, -24, 48,
    -- layer=1 filter=134 channel=17
    16, -19, -32, -5, -30, -3, -23, -30, -25,
    -- layer=1 filter=134 channel=18
    22, 29, 31, 19, -2, -71, -28, -27, -12,
    -- layer=1 filter=134 channel=19
    48, 31, 85, -8, 98, 41, 19, 24, 11,
    -- layer=1 filter=134 channel=20
    25, -12, 0, -9, -12, 35, -16, -19, 11,
    -- layer=1 filter=134 channel=21
    15, 0, -22, -26, -39, 16, -32, 7, 34,
    -- layer=1 filter=134 channel=22
    32, 5, -29, -6, -60, 15, -35, -18, 16,
    -- layer=1 filter=134 channel=23
    8, -62, -53, -117, 1, -39, -48, -8, -60,
    -- layer=1 filter=134 channel=24
    -9, -18, 16, -19, 36, 22, 12, 16, -41,
    -- layer=1 filter=134 channel=25
    65, -4, -36, -86, -2, 65, -54, 39, 66,
    -- layer=1 filter=134 channel=26
    -42, 8, 16, 5, 30, -37, 40, -43, -94,
    -- layer=1 filter=134 channel=27
    -4, -58, -72, -12, -62, -2, -42, -3, 7,
    -- layer=1 filter=134 channel=28
    -17, -58, -56, -88, -79, 26, -93, 27, 51,
    -- layer=1 filter=134 channel=29
    44, -19, 26, -7, -37, 22, -6, 38, 90,
    -- layer=1 filter=134 channel=30
    20, 26, 64, 41, 52, -29, 15, -18, -24,
    -- layer=1 filter=134 channel=31
    40, 43, 30, 36, -15, -71, 6, -43, -18,
    -- layer=1 filter=134 channel=32
    -41, 46, 22, 23, 45, -51, 44, -27, -90,
    -- layer=1 filter=134 channel=33
    -13, -24, 21, 8, 2, 37, -1, -10, -26,
    -- layer=1 filter=134 channel=34
    -11, -2, -2, -19, -30, -22, -14, -27, -32,
    -- layer=1 filter=134 channel=35
    -1, -5, -16, -24, -9, -14, 0, 0, -12,
    -- layer=1 filter=134 channel=36
    -1, -25, -49, -8, -40, -45, -14, -35, -13,
    -- layer=1 filter=134 channel=37
    38, -32, -37, -77, -33, 40, -41, -8, 28,
    -- layer=1 filter=134 channel=38
    -4, -6, 20, 0, -11, 3, -1, 5, 8,
    -- layer=1 filter=134 channel=39
    7, 3, -22, 6, -25, -39, -9, -11, -4,
    -- layer=1 filter=134 channel=40
    6, 28, 39, 13, -24, -50, -55, -29, -5,
    -- layer=1 filter=134 channel=41
    -36, 53, 64, 9, 99, 15, 19, 31, -118,
    -- layer=1 filter=134 channel=42
    -62, -93, 1, -26, 19, 47, 14, 54, 10,
    -- layer=1 filter=134 channel=43
    79, 10, -52, -55, -62, 59, -56, 3, 35,
    -- layer=1 filter=134 channel=44
    -17, 43, -7, 28, 6, -78, 29, -35, -111,
    -- layer=1 filter=134 channel=45
    8, 1, -26, -26, -18, 2, 9, -23, -26,
    -- layer=1 filter=134 channel=46
    7, -39, 2, -12, 6, 6, -22, -4, -38,
    -- layer=1 filter=134 channel=47
    -18, -10, -8, -20, 48, -24, 27, -20, -89,
    -- layer=1 filter=134 channel=48
    11, -8, 11, -18, 4, 4, -29, 27, 15,
    -- layer=1 filter=134 channel=49
    -31, -28, 38, -3, -4, -6, 13, -9, -17,
    -- layer=1 filter=134 channel=50
    25, 12, 30, 3, 12, -6, 15, 16, 23,
    -- layer=1 filter=134 channel=51
    8, -28, -10, -26, -38, 26, -37, 27, 50,
    -- layer=1 filter=134 channel=52
    15, 14, 9, 22, 47, -30, 49, 36, 38,
    -- layer=1 filter=134 channel=53
    4, 12, -15, -3, 11, -2, -11, -8, 9,
    -- layer=1 filter=134 channel=54
    68, -30, -2, -88, 38, 86, -26, 49, 69,
    -- layer=1 filter=134 channel=55
    4, -22, -48, -10, -13, -2, -25, -19, -19,
    -- layer=1 filter=134 channel=56
    6, 7, 1, -5, 1, -11, -11, -3, 5,
    -- layer=1 filter=134 channel=57
    -57, -105, -32, -97, -47, 18, -68, 26, 40,
    -- layer=1 filter=134 channel=58
    24, -74, -4, -135, 19, 30, -51, 46, -3,
    -- layer=1 filter=134 channel=59
    18, 5, -13, -2, -4, 0, -5, -5, -10,
    -- layer=1 filter=134 channel=60
    -15, -16, -2, -1, 24, -2, -23, 17, 5,
    -- layer=1 filter=134 channel=61
    2, -11, -7, -8, 6, 5, 0, 13, -8,
    -- layer=1 filter=134 channel=62
    72, -12, -28, -69, -29, 54, -28, 0, 38,
    -- layer=1 filter=134 channel=63
    4, 9, -14, 21, -22, -75, 5, -45, 0,
    -- layer=1 filter=134 channel=64
    37, 23, -8, 13, -28, 18, -35, 5, 24,
    -- layer=1 filter=134 channel=65
    -4, -4, -7, -2, 4, 18, -3, 27, 44,
    -- layer=1 filter=134 channel=66
    0, -17, -32, 6, -34, -12, 3, -12, 5,
    -- layer=1 filter=134 channel=67
    64, 30, 28, 15, 2, 4, 28, 4, 13,
    -- layer=1 filter=134 channel=68
    -22, 49, -11, 33, 0, -62, 32, -53, -75,
    -- layer=1 filter=134 channel=69
    -4, -20, -55, -75, -6, 5, -10, -8, -16,
    -- layer=1 filter=134 channel=70
    20, 20, 48, 0, -29, -53, -37, -93, -20,
    -- layer=1 filter=134 channel=71
    -15, -28, -17, -45, -26, 29, -13, 26, 24,
    -- layer=1 filter=134 channel=72
    48, 25, 56, 26, 54, 7, 0, 6, -17,
    -- layer=1 filter=134 channel=73
    4, -9, 9, 5, 1, -11, -10, 7, -2,
    -- layer=1 filter=134 channel=74
    23, 80, 39, 78, -7, -85, 0, -63, -18,
    -- layer=1 filter=134 channel=75
    47, 39, 24, 1, -23, -60, 1, -16, -24,
    -- layer=1 filter=134 channel=76
    -4, 32, 0, 48, 13, -42, 11, -41, -11,
    -- layer=1 filter=134 channel=77
    8, 5, -28, -32, -40, 10, 1, 27, 39,
    -- layer=1 filter=134 channel=78
    -35, -20, -9, -11, -14, 9, -2, -18, 20,
    -- layer=1 filter=134 channel=79
    68, -6, -23, -68, -12, 32, -35, 1, 29,
    -- layer=1 filter=134 channel=80
    15, -13, -17, -9, 21, 6, 3, 0, 9,
    -- layer=1 filter=134 channel=81
    6, -14, -19, -40, -49, 15, -29, 18, 27,
    -- layer=1 filter=134 channel=82
    0, 6, -1, -7, -23, 14, -7, 7, 10,
    -- layer=1 filter=134 channel=83
    4, 6, -58, -19, -21, -23, -36, -16, -31,
    -- layer=1 filter=134 channel=84
    13, 75, 41, 61, 14, -110, 12, -60, -42,
    -- layer=1 filter=134 channel=85
    24, -28, 36, -56, 39, 17, -17, 30, -20,
    -- layer=1 filter=134 channel=86
    5, -29, -39, -5, -31, -13, -15, -18, 10,
    -- layer=1 filter=134 channel=87
    41, 23, 82, 14, 117, 43, 6, 10, -19,
    -- layer=1 filter=134 channel=88
    -13, -15, 32, 2, 3, 29, 26, 43, 17,
    -- layer=1 filter=134 channel=89
    8, 49, 24, 35, -12, -35, 11, -11, 12,
    -- layer=1 filter=134 channel=90
    -11, 20, -30, 14, 18, -59, 24, -41, -104,
    -- layer=1 filter=134 channel=91
    8, 1, 15, 7, 6, 3, -22, -1, 10,
    -- layer=1 filter=134 channel=92
    -52, 35, -39, -14, 71, -49, 33, 5, -46,
    -- layer=1 filter=134 channel=93
    27, 2, -11, -16, -23, 18, -15, 0, 13,
    -- layer=1 filter=134 channel=94
    -7, -31, -45, 0, -61, -24, -8, -50, -1,
    -- layer=1 filter=134 channel=95
    7, 61, 30, 44, 9, -109, 31, -77, -7,
    -- layer=1 filter=134 channel=96
    16, 16, 2, 6, 2, 1, 22, 4, -18,
    -- layer=1 filter=134 channel=97
    34, 5, -39, -2, -14, 6, -12, -13, 33,
    -- layer=1 filter=134 channel=98
    52, 16, -51, -27, -30, 70, -53, -17, 38,
    -- layer=1 filter=134 channel=99
    -58, -42, -49, -81, -79, -39, -96, -13, 16,
    -- layer=1 filter=134 channel=100
    -5, 22, -15, 11, -27, -51, 7, -26, -11,
    -- layer=1 filter=134 channel=101
    5, 31, 25, 26, -19, -10, -3, -18, 26,
    -- layer=1 filter=134 channel=102
    14, 1, -6, 32, -19, -9, -8, -20, 17,
    -- layer=1 filter=134 channel=103
    10, 3, -17, 6, 0, -41, 0, 11, 9,
    -- layer=1 filter=134 channel=104
    20, -1, 33, -35, 53, -44, -5, 9, -49,
    -- layer=1 filter=134 channel=105
    4, -8, -29, 1, -34, -14, -32, -14, 31,
    -- layer=1 filter=134 channel=106
    -3, 48, 28, 44, 9, -58, 14, -37, -57,
    -- layer=1 filter=134 channel=107
    5, 4, 5, -16, 3, 7, 5, 10, 10,
    -- layer=1 filter=134 channel=108
    -54, 27, 17, 8, 41, -62, 24, -20, -105,
    -- layer=1 filter=134 channel=109
    -3, 7, 0, 5, 1, 6, -2, -3, 0,
    -- layer=1 filter=134 channel=110
    2, 5, -10, -1, -14, 1, -10, -2, 0,
    -- layer=1 filter=134 channel=111
    12, 56, 42, 41, 5, -122, -24, -77, -41,
    -- layer=1 filter=134 channel=112
    43, 70, 36, 51, -8, -112, -17, -57, -22,
    -- layer=1 filter=134 channel=113
    -18, -72, -18, -18, -52, 23, 7, -9, -16,
    -- layer=1 filter=134 channel=114
    16, 1, -54, -43, -52, -48, -24, -14, 14,
    -- layer=1 filter=134 channel=115
    -25, -35, -31, -31, -32, 11, -63, -3, 12,
    -- layer=1 filter=134 channel=116
    8, -8, 1, 6, 4, 9, 2, -8, 9,
    -- layer=1 filter=134 channel=117
    6, 30, 13, 36, -29, -136, -95, -95, -65,
    -- layer=1 filter=134 channel=118
    20, 56, 37, 64, 41, -89, 24, -53, -35,
    -- layer=1 filter=134 channel=119
    -32, 29, 14, 31, 56, -43, 40, -14, -90,
    -- layer=1 filter=134 channel=120
    31, -36, -19, -67, -35, 43, -47, 27, 40,
    -- layer=1 filter=134 channel=121
    2, -16, 31, -33, -15, -26, -36, -23, -66,
    -- layer=1 filter=134 channel=122
    7, 6, 2, 1, 3, -9, -9, -2, 1,
    -- layer=1 filter=134 channel=123
    -5, -29, -13, -31, -14, -32, -33, 2, -20,
    -- layer=1 filter=134 channel=124
    2, -18, 15, 3, 13, 11, 16, 22, 1,
    -- layer=1 filter=134 channel=125
    7, -13, 35, 22, -25, -40, -13, -54, 15,
    -- layer=1 filter=134 channel=126
    50, 0, -143, -14, -46, 35, -71, -44, -12,
    -- layer=1 filter=134 channel=127
    12, 51, 41, 63, 13, -92, 22, -80, -13,
    -- layer=1 filter=135 channel=0
    -25, -43, -40, -20, -20, -33, 7, 0, 9,
    -- layer=1 filter=135 channel=1
    -30, -8, -17, 12, -32, -53, 63, 55, 36,
    -- layer=1 filter=135 channel=2
    -32, -48, -39, -50, -45, -30, -85, -31, -46,
    -- layer=1 filter=135 channel=3
    -1, 5, -9, 1, -1, 5, 5, 8, 0,
    -- layer=1 filter=135 channel=4
    -11, -2, -16, -4, -22, -13, 3, -4, 12,
    -- layer=1 filter=135 channel=5
    -43, 4, -9, 2, -30, -32, 71, 88, 65,
    -- layer=1 filter=135 channel=6
    -17, -21, -45, -36, -13, -57, -58, -96, -112,
    -- layer=1 filter=135 channel=7
    -27, -54, -62, -29, -101, -29, -38, -62, -57,
    -- layer=1 filter=135 channel=8
    -31, -1, -20, -12, -37, -49, 65, 61, 33,
    -- layer=1 filter=135 channel=9
    -6, -34, 1, -47, -2, 0, -11, 5, 16,
    -- layer=1 filter=135 channel=10
    2, -65, -33, 6, -93, -41, 0, -49, -37,
    -- layer=1 filter=135 channel=11
    -81, -73, -107, -36, -80, -75, 6, -21, -36,
    -- layer=1 filter=135 channel=12
    -38, 0, -8, -24, 22, -11, 11, 22, -24,
    -- layer=1 filter=135 channel=13
    2, -14, 0, -20, -29, -21, 13, -5, 5,
    -- layer=1 filter=135 channel=14
    -18, -20, -29, -9, -51, 4, -2, -42, -16,
    -- layer=1 filter=135 channel=15
    12, 31, 52, -36, -27, 29, -18, 12, 5,
    -- layer=1 filter=135 channel=16
    -23, -18, -11, 16, -9, -44, 75, 75, 47,
    -- layer=1 filter=135 channel=17
    -15, -18, -33, -26, -11, -10, 43, 25, 20,
    -- layer=1 filter=135 channel=18
    -68, -42, -65, -41, -29, -85, 13, -1, -9,
    -- layer=1 filter=135 channel=19
    19, -21, 2, 21, -36, 4, 105, 67, 71,
    -- layer=1 filter=135 channel=20
    -4, -16, -24, -32, -34, -36, 13, 28, 6,
    -- layer=1 filter=135 channel=21
    6, 9, 24, 7, 22, 1, 26, 13, 4,
    -- layer=1 filter=135 channel=22
    2, -15, -30, -40, -43, -37, 25, 3, 10,
    -- layer=1 filter=135 channel=23
    -52, -42, 11, -41, -53, 11, -42, -15, -12,
    -- layer=1 filter=135 channel=24
    0, 6, 40, 1, 23, 9, 36, 27, 34,
    -- layer=1 filter=135 channel=25
    -26, -54, -42, -3, -78, -35, 31, 28, 12,
    -- layer=1 filter=135 channel=26
    -27, -20, 0, -51, -62, 3, -13, -12, -3,
    -- layer=1 filter=135 channel=27
    -29, -29, -34, -23, -13, -35, -20, -10, -22,
    -- layer=1 filter=135 channel=28
    7, -28, -35, -9, -57, -35, 26, -15, -11,
    -- layer=1 filter=135 channel=29
    3, 33, 0, 10, 7, 13, -3, 22, 13,
    -- layer=1 filter=135 channel=30
    -4, -10, 22, -23, -22, -35, 25, -1, 6,
    -- layer=1 filter=135 channel=31
    -69, -35, -60, -21, 8, -15, 20, 40, -21,
    -- layer=1 filter=135 channel=32
    -18, -57, 42, -24, -66, 32, -26, -17, -15,
    -- layer=1 filter=135 channel=33
    30, 30, 5, 69, 43, 12, 0, 23, -1,
    -- layer=1 filter=135 channel=34
    12, 17, 14, 58, 51, 41, 40, 15, 6,
    -- layer=1 filter=135 channel=35
    9, -1, -1, -4, -15, 5, 16, 4, 24,
    -- layer=1 filter=135 channel=36
    -73, -91, -106, -48, -86, -104, 12, -31, -19,
    -- layer=1 filter=135 channel=37
    -11, -4, -7, 20, -29, -28, 76, 71, 60,
    -- layer=1 filter=135 channel=38
    16, 7, 2, -9, 8, -18, -1, -9, 0,
    -- layer=1 filter=135 channel=39
    -38, -55, -70, -9, -53, -17, 37, 30, -9,
    -- layer=1 filter=135 channel=40
    -23, -21, -53, 17, 12, -11, -45, -41, -40,
    -- layer=1 filter=135 channel=41
    -23, -48, 56, -24, -19, 17, -15, -6, 27,
    -- layer=1 filter=135 channel=42
    -27, -56, -49, -29, -68, -33, -47, -48, -12,
    -- layer=1 filter=135 channel=43
    -17, 1, -24, 2, -43, -54, 65, 42, 24,
    -- layer=1 filter=135 channel=44
    -34, -38, 29, -17, -77, 21, -14, -4, 18,
    -- layer=1 filter=135 channel=45
    -10, -18, 3, -15, -25, 3, 29, 17, 24,
    -- layer=1 filter=135 channel=46
    -1, -15, 15, -2, -46, -16, 65, 77, 48,
    -- layer=1 filter=135 channel=47
    -50, -100, 51, -60, -44, 2, -69, -2, 10,
    -- layer=1 filter=135 channel=48
    3, 25, 6, -9, 7, -7, -9, -6, -19,
    -- layer=1 filter=135 channel=49
    -16, -18, 13, 0, 17, 0, -34, -24, -14,
    -- layer=1 filter=135 channel=50
    -13, -11, 10, -9, -1, -5, -1, 3, 6,
    -- layer=1 filter=135 channel=51
    12, 19, -15, 12, -5, 0, -20, -39, -29,
    -- layer=1 filter=135 channel=52
    34, 38, -4, 54, 24, 18, -4, -23, 1,
    -- layer=1 filter=135 channel=53
    16, 3, 12, 19, 1, 0, 14, 4, 17,
    -- layer=1 filter=135 channel=54
    -9, -35, -30, 4, -97, -49, 35, 34, 13,
    -- layer=1 filter=135 channel=55
    -62, -50, -42, -17, -36, -39, 15, -1, 0,
    -- layer=1 filter=135 channel=56
    -7, -11, 8, -5, 2, 6, 3, 4, 5,
    -- layer=1 filter=135 channel=57
    -17, -62, -37, 1, -65, -35, 8, -67, -31,
    -- layer=1 filter=135 channel=58
    -66, -66, -4, -37, -96, -14, -17, -42, 11,
    -- layer=1 filter=135 channel=59
    -14, 0, -5, -17, 1, -4, -6, -8, -14,
    -- layer=1 filter=135 channel=60
    4, 18, -25, -3, 14, -7, 0, -13, -4,
    -- layer=1 filter=135 channel=61
    5, -2, 0, 1, 2, -1, 1, -6, -4,
    -- layer=1 filter=135 channel=62
    -32, -13, -14, 16, -19, -41, 82, 64, 61,
    -- layer=1 filter=135 channel=63
    -44, -42, -62, -25, -36, -53, -3, -32, -53,
    -- layer=1 filter=135 channel=64
    -6, -16, -21, -12, -11, -27, 6, 0, -11,
    -- layer=1 filter=135 channel=65
    8, -2, 11, -10, 8, 2, -11, 2, -1,
    -- layer=1 filter=135 channel=66
    -20, -39, -41, -10, -5, -11, 24, 31, 5,
    -- layer=1 filter=135 channel=67
    -31, -17, -34, -42, -20, -25, -52, -42, -65,
    -- layer=1 filter=135 channel=68
    -39, -29, 6, -35, -50, 32, -30, -32, 13,
    -- layer=1 filter=135 channel=69
    -29, -14, 16, -19, -31, -3, 51, 67, 33,
    -- layer=1 filter=135 channel=70
    -20, 12, -32, 63, 79, 15, -27, -21, 1,
    -- layer=1 filter=135 channel=71
    15, 40, 11, 24, 16, 16, 26, 34, 21,
    -- layer=1 filter=135 channel=72
    5, -39, 1, -60, -71, -73, 87, -48, 15,
    -- layer=1 filter=135 channel=73
    34, -9, 0, 5, -1, -3, -17, -4, -11,
    -- layer=1 filter=135 channel=74
    -3, 18, -7, 13, 22, 11, -33, -2, -7,
    -- layer=1 filter=135 channel=75
    -32, -10, -22, -61, -57, -42, -18, 17, -47,
    -- layer=1 filter=135 channel=76
    -40, -32, -17, -44, -63, -23, -11, -43, -17,
    -- layer=1 filter=135 channel=77
    3, 16, 24, 10, 3, 7, -1, 12, 3,
    -- layer=1 filter=135 channel=78
    0, -26, -14, -19, -20, -12, 10, 6, 0,
    -- layer=1 filter=135 channel=79
    -17, -3, -1, -8, -22, -46, 60, 53, 37,
    -- layer=1 filter=135 channel=80
    -7, 15, 24, -2, -19, -31, 39, 10, -7,
    -- layer=1 filter=135 channel=81
    1, 11, 9, -2, 13, 2, 20, 30, 17,
    -- layer=1 filter=135 channel=82
    28, 30, 11, 17, 24, 10, -10, -4, -6,
    -- layer=1 filter=135 channel=83
    14, -16, 0, -27, -21, 18, 38, 51, 45,
    -- layer=1 filter=135 channel=84
    -64, -31, -17, -15, -19, -55, -37, -52, -29,
    -- layer=1 filter=135 channel=85
    -69, -71, 16, -29, -83, -17, -12, -38, 2,
    -- layer=1 filter=135 channel=86
    -39, -53, -77, 11, -27, -22, 54, 49, 25,
    -- layer=1 filter=135 channel=87
    -3, -47, -12, 1, -4, -47, 73, 40, 77,
    -- layer=1 filter=135 channel=88
    -4, 13, 6, -11, 21, 4, -24, -10, -16,
    -- layer=1 filter=135 channel=89
    19, 27, 15, 3, 28, 19, -14, 1, -17,
    -- layer=1 filter=135 channel=90
    -48, -23, 16, -35, -69, 15, 10, 25, 30,
    -- layer=1 filter=135 channel=91
    3, 3, -4, -25, -1, -18, -45, -37, -36,
    -- layer=1 filter=135 channel=92
    -23, 6, 49, -29, -9, 55, -24, 15, 17,
    -- layer=1 filter=135 channel=93
    15, 28, 7, 14, 20, 3, 17, 23, 17,
    -- layer=1 filter=135 channel=94
    -18, -40, -61, -14, -10, -36, 14, -2, 1,
    -- layer=1 filter=135 channel=95
    -19, -11, 6, -14, -12, -41, -16, -21, -22,
    -- layer=1 filter=135 channel=96
    1, 0, -5, 5, -2, 8, 6, 3, -18,
    -- layer=1 filter=135 channel=97
    -5, 12, -2, 14, 9, 8, 32, 24, 7,
    -- layer=1 filter=135 channel=98
    -23, 0, -16, -8, -40, -73, 66, 33, 33,
    -- layer=1 filter=135 channel=99
    16, -8, 12, 33, -3, -11, 16, -32, -11,
    -- layer=1 filter=135 channel=100
    -50, -64, -78, -27, -85, -91, 41, 29, -21,
    -- layer=1 filter=135 channel=101
    7, 15, 2, -7, 1, -10, -11, -7, -12,
    -- layer=1 filter=135 channel=102
    -5, -8, -32, -16, -16, -28, -27, -11, -27,
    -- layer=1 filter=135 channel=103
    -66, -80, -70, -42, -32, -91, 21, 13, 4,
    -- layer=1 filter=135 channel=104
    -39, -59, 11, -16, -42, -55, -33, -7, -24,
    -- layer=1 filter=135 channel=105
    10, 0, -19, 5, 4, 5, 27, 1, 0,
    -- layer=1 filter=135 channel=106
    -1, -5, 18, -4, -3, -10, -35, -35, -30,
    -- layer=1 filter=135 channel=107
    11, -9, 12, -1, 13, 0, 0, -4, -9,
    -- layer=1 filter=135 channel=108
    -46, -43, 43, -28, -48, 37, 1, 33, 40,
    -- layer=1 filter=135 channel=109
    -6, -9, 7, -9, 0, -9, -4, 8, 9,
    -- layer=1 filter=135 channel=110
    -19, -5, -7, -20, 0, 1, -15, -18, -6,
    -- layer=1 filter=135 channel=111
    -15, -12, -12, 2, 27, -50, -7, -29, -7,
    -- layer=1 filter=135 channel=112
    -27, -7, -5, 29, 23, -10, -55, -15, -38,
    -- layer=1 filter=135 channel=113
    -28, -34, -44, -17, -32, -22, -19, -36, -3,
    -- layer=1 filter=135 channel=114
    -10, 0, 0, 15, 8, -32, 39, 60, 20,
    -- layer=1 filter=135 channel=115
    -13, -62, -45, 9, -34, -29, 40, -2, -1,
    -- layer=1 filter=135 channel=116
    0, 5, -2, -4, 2, -1, -8, -10, 7,
    -- layer=1 filter=135 channel=117
    -19, -7, -28, 38, 46, -4, -64, -16, -29,
    -- layer=1 filter=135 channel=118
    -22, -6, 15, -6, 12, -21, -40, -44, -27,
    -- layer=1 filter=135 channel=119
    -37, -36, 36, -34, -53, 25, -15, -28, -7,
    -- layer=1 filter=135 channel=120
    15, 5, 0, 3, 20, 5, 13, 14, 14,
    -- layer=1 filter=135 channel=121
    12, -19, -17, -35, -35, -21, 86, 78, 55,
    -- layer=1 filter=135 channel=122
    4, -4, 0, -2, 9, 5, 4, 7, 6,
    -- layer=1 filter=135 channel=123
    -9, -23, -37, -25, -53, -49, 11, 20, 18,
    -- layer=1 filter=135 channel=124
    -3, 2, -1, 5, 29, 0, 20, 20, 8,
    -- layer=1 filter=135 channel=125
    -37, -7, -29, 0, 28, 8, -55, -9, -19,
    -- layer=1 filter=135 channel=126
    -25, -13, -15, -4, -39, -16, 50, 47, 26,
    -- layer=1 filter=135 channel=127
    -38, -22, -3, -15, -16, -49, -7, -20, -25,
    -- layer=1 filter=136 channel=0
    -46, 1, -25, -30, -13, -28, -21, -1, 0,
    -- layer=1 filter=136 channel=1
    34, -61, -40, -27, 11, -27, 20, -1, -12,
    -- layer=1 filter=136 channel=2
    -39, 25, 27, -62, 39, 42, -104, -51, 5,
    -- layer=1 filter=136 channel=3
    9, -2, 2, -8, 4, -4, -10, 6, -10,
    -- layer=1 filter=136 channel=4
    -9, 8, 5, 0, -1, 8, -11, 2, -10,
    -- layer=1 filter=136 channel=5
    28, -49, -37, -25, 26, -11, -8, -12, -21,
    -- layer=1 filter=136 channel=6
    -37, -34, -74, -12, -66, -44, 27, -63, -60,
    -- layer=1 filter=136 channel=7
    -3, -54, -47, -72, -14, -35, -49, 32, -22,
    -- layer=1 filter=136 channel=8
    10, -83, -39, -12, 17, -28, -16, -21, 2,
    -- layer=1 filter=136 channel=9
    -33, 1, 17, -52, -37, -45, -25, -39, -22,
    -- layer=1 filter=136 channel=10
    -42, -36, -42, -75, -1, -49, -41, 26, -39,
    -- layer=1 filter=136 channel=11
    -10, -21, -12, -47, -52, 17, -26, -23, 31,
    -- layer=1 filter=136 channel=12
    0, 38, -60, -104, -56, 62, -65, -95, -84,
    -- layer=1 filter=136 channel=13
    42, -71, -53, 73, -33, -11, 76, 34, -19,
    -- layer=1 filter=136 channel=14
    26, -16, -65, -66, -3, 37, -70, -33, -50,
    -- layer=1 filter=136 channel=15
    85, -82, -21, 54, 45, 32, 99, 64, -42,
    -- layer=1 filter=136 channel=16
    23, -28, -35, 10, 14, -5, -17, -12, 9,
    -- layer=1 filter=136 channel=17
    -58, -60, -52, 18, -56, -7, -12, -58, 6,
    -- layer=1 filter=136 channel=18
    29, 31, -16, -90, -25, 23, -63, -73, -30,
    -- layer=1 filter=136 channel=19
    -61, -24, -49, -40, -7, -51, -46, -38, -67,
    -- layer=1 filter=136 channel=20
    12, -67, -58, 44, -29, -52, 62, -11, -23,
    -- layer=1 filter=136 channel=21
    0, 27, -13, -17, 30, 2, 5, 20, -2,
    -- layer=1 filter=136 channel=22
    -22, -86, -71, 33, -4, -22, 38, 0, 15,
    -- layer=1 filter=136 channel=23
    53, -123, -16, 29, -39, 2, 51, 4, -52,
    -- layer=1 filter=136 channel=24
    25, 6, 8, 40, 8, 4, 22, 15, 12,
    -- layer=1 filter=136 channel=25
    -58, -48, -46, -74, 23, -40, -54, 25, 9,
    -- layer=1 filter=136 channel=26
    48, -98, -42, 79, -31, 22, 72, 38, -42,
    -- layer=1 filter=136 channel=27
    -40, -39, -24, -61, -32, -51, -78, -66, -73,
    -- layer=1 filter=136 channel=28
    9, -15, -30, -95, 19, -55, 7, 3, -36,
    -- layer=1 filter=136 channel=29
    -29, -51, -73, -30, -41, -61, -22, -47, -62,
    -- layer=1 filter=136 channel=30
    -2, 30, -12, -103, -12, -7, -86, -114, -74,
    -- layer=1 filter=136 channel=31
    8, 29, -34, -28, -1, 42, -11, -53, -20,
    -- layer=1 filter=136 channel=32
    68, -89, -8, 73, -30, -47, 51, 47, -59,
    -- layer=1 filter=136 channel=33
    1, 12, 13, 18, -7, 26, -19, -31, -21,
    -- layer=1 filter=136 channel=34
    31, -22, -11, 19, -20, 14, 25, 17, 5,
    -- layer=1 filter=136 channel=35
    16, -24, -16, -4, 0, 7, 0, 9, 7,
    -- layer=1 filter=136 channel=36
    -33, -24, -1, -65, -54, 28, -55, -49, 24,
    -- layer=1 filter=136 channel=37
    -3, -38, -48, 2, 19, -12, -24, -20, -6,
    -- layer=1 filter=136 channel=38
    5, -13, -13, 38, -13, -30, 58, 11, -18,
    -- layer=1 filter=136 channel=39
    -38, -26, -26, -48, 5, -18, -65, -91, -2,
    -- layer=1 filter=136 channel=40
    -20, 7, -28, -40, -44, -11, 25, -61, -32,
    -- layer=1 filter=136 channel=41
    22, -63, -5, 75, -91, -78, 53, -16, -96,
    -- layer=1 filter=136 channel=42
    -41, 18, 15, -24, 31, 52, -99, -48, 10,
    -- layer=1 filter=136 channel=43
    -28, -61, -67, -26, 16, -32, -24, -20, 11,
    -- layer=1 filter=136 channel=44
    51, -114, -47, 54, -36, -10, 49, 44, -36,
    -- layer=1 filter=136 channel=45
    29, -51, -45, 56, 4, 16, 41, 19, -17,
    -- layer=1 filter=136 channel=46
    -47, -57, -42, -36, 20, 31, -34, -20, -26,
    -- layer=1 filter=136 channel=47
    65, -49, 14, 86, 33, -49, 78, 57, -11,
    -- layer=1 filter=136 channel=48
    -8, 16, -7, -12, -17, -28, 2, 3, -32,
    -- layer=1 filter=136 channel=49
    -5, 5, -5, 19, 11, 19, -2, 5, 18,
    -- layer=1 filter=136 channel=50
    12, 27, 38, -12, 5, 10, -15, 7, -3,
    -- layer=1 filter=136 channel=51
    -21, 9, -17, -36, -10, -27, 13, -11, -17,
    -- layer=1 filter=136 channel=52
    -1, 5, 24, -20, -24, -35, -11, 6, 3,
    -- layer=1 filter=136 channel=53
    -1, -13, 11, 2, -9, 19, -12, -7, -4,
    -- layer=1 filter=136 channel=54
    -38, -38, -48, -74, 27, -51, -36, 27, 16,
    -- layer=1 filter=136 channel=55
    18, -22, 15, 13, -3, 25, 0, -4, 44,
    -- layer=1 filter=136 channel=56
    1, 8, 6, 0, 6, -7, -2, 0, 3,
    -- layer=1 filter=136 channel=57
    -33, -10, -45, -37, -17, -48, -29, 14, -6,
    -- layer=1 filter=136 channel=58
    -43, -98, -15, -39, -11, -27, 1, -6, -1,
    -- layer=1 filter=136 channel=59
    7, 0, -1, 6, 7, -4, 14, -4, -9,
    -- layer=1 filter=136 channel=60
    -6, 6, 30, -20, 8, 10, -9, 3, -12,
    -- layer=1 filter=136 channel=61
    -10, -11, -3, -4, -8, -9, 8, 5, -7,
    -- layer=1 filter=136 channel=62
    0, -74, -62, 23, -5, -23, -11, -39, 3,
    -- layer=1 filter=136 channel=63
    10, -9, -5, -20, -28, 4, -23, -69, 0,
    -- layer=1 filter=136 channel=64
    -29, -25, -52, -48, -34, -85, 3, -35, -31,
    -- layer=1 filter=136 channel=65
    -7, -4, -14, 4, 12, -27, 26, 3, -7,
    -- layer=1 filter=136 channel=66
    -43, -30, -13, -72, -39, -7, -43, -35, -10,
    -- layer=1 filter=136 channel=67
    27, 43, -3, -1, 26, 0, 3, 23, -3,
    -- layer=1 filter=136 channel=68
    40, -88, -56, 53, -59, -4, 51, 44, -24,
    -- layer=1 filter=136 channel=69
    51, -78, -35, 61, 27, 20, 64, 0, -38,
    -- layer=1 filter=136 channel=70
    -22, -3, -43, -74, -59, -22, 13, -54, -44,
    -- layer=1 filter=136 channel=71
    5, 12, 13, -12, 19, 5, -8, 0, 4,
    -- layer=1 filter=136 channel=72
    -25, -21, -10, -79, -9, -9, -62, -71, -71,
    -- layer=1 filter=136 channel=73
    -14, -10, 3, -1, -2, -22, -12, -6, 2,
    -- layer=1 filter=136 channel=74
    -8, 27, -36, -28, -57, -56, -27, -40, -70,
    -- layer=1 filter=136 channel=75
    0, 8, -25, -65, -14, 60, -89, -124, -34,
    -- layer=1 filter=136 channel=76
    6, -39, -26, 37, -69, -28, 0, -21, -25,
    -- layer=1 filter=136 channel=77
    -7, 29, 7, 12, 20, -21, 30, 1, -15,
    -- layer=1 filter=136 channel=78
    8, -12, -23, -4, 15, -10, 11, 11, -18,
    -- layer=1 filter=136 channel=79
    21, -37, -54, 27, 21, -11, -1, -16, 6,
    -- layer=1 filter=136 channel=80
    -4, -50, -17, 15, 31, -21, -27, -1, -37,
    -- layer=1 filter=136 channel=81
    -16, 22, 7, -2, 29, -9, -3, 9, 6,
    -- layer=1 filter=136 channel=82
    23, 12, -2, 40, 8, -20, 20, 25, 3,
    -- layer=1 filter=136 channel=83
    33, -127, -66, 62, -3, 2, 47, -10, -55,
    -- layer=1 filter=136 channel=84
    37, 20, -11, 30, -100, -68, 3, -77, -28,
    -- layer=1 filter=136 channel=85
    -40, -31, -11, -22, -29, -21, 35, -11, -5,
    -- layer=1 filter=136 channel=86
    -36, -47, -11, -69, -17, 6, -35, -49, 9,
    -- layer=1 filter=136 channel=87
    -65, -20, -23, -90, 1, -73, -66, -59, -61,
    -- layer=1 filter=136 channel=88
    -39, 11, 23, -15, 5, -2, -25, -17, 0,
    -- layer=1 filter=136 channel=89
    25, 17, -7, 33, 37, -18, 25, 20, -3,
    -- layer=1 filter=136 channel=90
    49, -116, -51, 80, -46, 3, 63, 52, -26,
    -- layer=1 filter=136 channel=91
    -18, -5, -27, 1, -1, -43, 43, -6, -33,
    -- layer=1 filter=136 channel=92
    68, -114, -16, 81, -12, -29, 61, 73, -63,
    -- layer=1 filter=136 channel=93
    1, 0, 5, 10, 9, -11, 18, -2, -11,
    -- layer=1 filter=136 channel=94
    -24, -8, -27, -63, 1, -2, -12, -17, -24,
    -- layer=1 filter=136 channel=95
    38, 11, -16, -24, -58, -32, -65, -160, -63,
    -- layer=1 filter=136 channel=96
    11, 9, 7, 12, 5, -8, 10, -6, -14,
    -- layer=1 filter=136 channel=97
    -14, -28, -21, -16, -17, -24, 2, -21, -17,
    -- layer=1 filter=136 channel=98
    -31, -77, -64, 18, 7, -32, -10, -17, 23,
    -- layer=1 filter=136 channel=99
    1, 21, 9, -75, -44, -41, 52, -47, -61,
    -- layer=1 filter=136 channel=100
    12, -23, -6, 4, -32, 5, 1, -46, 0,
    -- layer=1 filter=136 channel=101
    8, -11, -33, 28, -8, -29, 33, 5, -27,
    -- layer=1 filter=136 channel=102
    -52, -29, -11, -39, -30, -27, -4, -28, -21,
    -- layer=1 filter=136 channel=103
    -5, -5, 4, -52, -92, -34, -1, -59, -22,
    -- layer=1 filter=136 channel=104
    11, -72, 1, 1, -26, -50, 40, -21, -60,
    -- layer=1 filter=136 channel=105
    -56, -3, -14, -71, -11, -37, -24, -15, -25,
    -- layer=1 filter=136 channel=106
    36, -40, -29, 61, -20, -30, 69, 46, -27,
    -- layer=1 filter=136 channel=107
    -9, -3, 9, -12, -14, 7, 5, -12, -6,
    -- layer=1 filter=136 channel=108
    74, -115, -33, 82, -19, -2, 55, 47, -42,
    -- layer=1 filter=136 channel=109
    -6, 8, 9, 4, 7, 2, 1, -8, -7,
    -- layer=1 filter=136 channel=110
    -6, -2, -13, 1, -7, 6, 5, 12, -11,
    -- layer=1 filter=136 channel=111
    25, 53, -4, -67, -60, -35, -70, -97, -64,
    -- layer=1 filter=136 channel=112
    37, 37, -22, -10, -20, -63, -18, -37, 25,
    -- layer=1 filter=136 channel=113
    -41, -36, -38, 14, -11, 5, -4, -48, -14,
    -- layer=1 filter=136 channel=114
    20, -70, -27, -23, 23, 18, -17, -31, -26,
    -- layer=1 filter=136 channel=115
    2, -24, -12, -60, -5, -25, -52, -2, 7,
    -- layer=1 filter=136 channel=116
    5, -2, 7, 2, 2, -6, 9, -6, -2,
    -- layer=1 filter=136 channel=117
    73, 41, 26, -4, -76, -39, -33, 1, 8,
    -- layer=1 filter=136 channel=118
    18, 33, 3, -13, -76, -36, -14, -95, -71,
    -- layer=1 filter=136 channel=119
    50, -85, -22, 74, -59, -34, 48, 50, -34,
    -- layer=1 filter=136 channel=120
    -48, 4, -19, -30, 25, -27, -2, 18, 12,
    -- layer=1 filter=136 channel=121
    14, 7, 6, -43, 41, 38, -77, -29, -12,
    -- layer=1 filter=136 channel=122
    -8, -2, 4, -7, -2, 0, -1, -3, 0,
    -- layer=1 filter=136 channel=123
    -8, -1, 7, -48, 24, 46, -97, -51, 10,
    -- layer=1 filter=136 channel=124
    22, 22, 11, -11, 28, 18, -2, 11, 8,
    -- layer=1 filter=136 channel=125
    -26, -8, -31, -14, -62, -33, 0, -56, -52,
    -- layer=1 filter=136 channel=126
    -17, -57, -51, 42, -39, -42, 17, -10, 23,
    -- layer=1 filter=136 channel=127
    29, 25, -18, -59, -48, 13, -67, -123, -65,
    -- layer=1 filter=137 channel=0
    -34, -35, -31, 8, 4, -46, 29, -4, -20,
    -- layer=1 filter=137 channel=1
    40, 10, -28, 51, -21, -41, 14, -19, -34,
    -- layer=1 filter=137 channel=2
    39, 68, 59, 28, 66, 69, 12, 66, 69,
    -- layer=1 filter=137 channel=3
    7, 8, 7, 5, 2, 12, -6, 0, -5,
    -- layer=1 filter=137 channel=4
    -10, 8, -3, 0, 7, 7, -11, 9, 7,
    -- layer=1 filter=137 channel=5
    63, 16, -19, 46, -8, -52, 2, -1, -13,
    -- layer=1 filter=137 channel=6
    27, -52, -53, 25, -25, -42, -3, -35, -41,
    -- layer=1 filter=137 channel=7
    11, -81, -41, 8, -92, -42, -76, -47, -61,
    -- layer=1 filter=137 channel=8
    54, 0, -41, 29, -39, -35, 6, -27, -19,
    -- layer=1 filter=137 channel=9
    6, -5, 25, -14, 47, 18, 32, 28, 46,
    -- layer=1 filter=137 channel=10
    40, -71, -44, 13, -72, -60, -59, -47, -46,
    -- layer=1 filter=137 channel=11
    -17, -20, -23, -8, -36, -12, 29, -7, -8,
    -- layer=1 filter=137 channel=12
    -17, 56, 0, 38, -12, 54, -13, 19, 23,
    -- layer=1 filter=137 channel=13
    11, -44, -55, 34, -7, -36, 38, 10, -29,
    -- layer=1 filter=137 channel=14
    14, 9, 22, 31, -19, 21, -32, -23, -36,
    -- layer=1 filter=137 channel=15
    120, 40, 39, 141, 42, 45, 102, 68, -13,
    -- layer=1 filter=137 channel=16
    58, -2, -38, 12, -55, -50, -1, -41, -28,
    -- layer=1 filter=137 channel=17
    -35, -39, -72, 6, -5, -52, 33, -34, -23,
    -- layer=1 filter=137 channel=18
    -47, -47, 1, -81, -33, -30, -41, 10, -18,
    -- layer=1 filter=137 channel=19
    -25, -43, -35, -21, -27, -55, -28, 14, 20,
    -- layer=1 filter=137 channel=20
    11, -35, -45, 28, -29, -38, 20, -15, -48,
    -- layer=1 filter=137 channel=21
    23, 10, -23, 2, -6, -22, -14, -20, -18,
    -- layer=1 filter=137 channel=22
    23, 9, -32, 47, -21, -18, 8, -16, -28,
    -- layer=1 filter=137 channel=23
    55, -61, 9, 73, -20, 26, 32, 60, -69,
    -- layer=1 filter=137 channel=24
    14, -7, -2, 25, -14, -23, 21, 1, -12,
    -- layer=1 filter=137 channel=25
    46, -54, -35, 23, -69, -56, -39, -15, -34,
    -- layer=1 filter=137 channel=26
    20, -59, -67, 59, -18, -37, 60, 29, -55,
    -- layer=1 filter=137 channel=27
    39, 38, 24, 29, 24, 21, 3, 17, 28,
    -- layer=1 filter=137 channel=28
    21, -57, -48, 3, -66, -58, -54, -40, -56,
    -- layer=1 filter=137 channel=29
    -30, -63, -46, -32, -57, -55, 9, -44, -67,
    -- layer=1 filter=137 channel=30
    -79, -97, -27, -99, -62, -69, -62, -51, -71,
    -- layer=1 filter=137 channel=31
    5, 32, 8, 28, 35, 47, 25, 33, 26,
    -- layer=1 filter=137 channel=32
    24, -67, -80, 41, -8, -33, 44, 74, -69,
    -- layer=1 filter=137 channel=33
    15, -11, 3, -6, -20, -19, -9, -3, -5,
    -- layer=1 filter=137 channel=34
    42, -5, -14, 20, 6, -2, 23, -2, -7,
    -- layer=1 filter=137 channel=35
    5, -7, 5, 12, 11, 3, 3, 4, 3,
    -- layer=1 filter=137 channel=36
    -42, -40, -22, -34, -29, -27, 16, -27, -5,
    -- layer=1 filter=137 channel=37
    49, 6, -16, -5, -27, -54, -12, -28, 7,
    -- layer=1 filter=137 channel=38
    -8, -39, -46, -15, -35, -48, 11, -54, -10,
    -- layer=1 filter=137 channel=39
    5, -7, -22, 13, 9, -38, -12, -30, -8,
    -- layer=1 filter=137 channel=40
    -10, -21, -2, -6, -6, -7, -47, -30, 3,
    -- layer=1 filter=137 channel=41
    14, -61, -36, 47, 12, -28, 63, 66, -26,
    -- layer=1 filter=137 channel=42
    36, 69, 63, 18, 61, 63, 18, 62, 66,
    -- layer=1 filter=137 channel=43
    12, -49, -76, 19, -80, -74, -36, -45, -28,
    -- layer=1 filter=137 channel=44
    14, -65, -96, 56, -14, -59, 59, 43, -72,
    -- layer=1 filter=137 channel=45
    46, 0, -30, 67, -14, -26, 43, 0, -29,
    -- layer=1 filter=137 channel=46
    43, 42, 38, 4, 39, 27, 25, 59, 66,
    -- layer=1 filter=137 channel=47
    69, -28, 29, 68, 35, -4, 37, 72, -15,
    -- layer=1 filter=137 channel=48
    -27, -80, -53, -16, -54, -60, -1, -63, -53,
    -- layer=1 filter=137 channel=49
    19, 6, 30, 14, 25, 25, 20, 49, 32,
    -- layer=1 filter=137 channel=50
    10, -1, 8, 17, 0, -16, 11, 3, 12,
    -- layer=1 filter=137 channel=51
    -18, -50, -28, -15, -61, -26, -65, -57, -48,
    -- layer=1 filter=137 channel=52
    3, 2, -25, -21, -33, -48, -13, -30, -38,
    -- layer=1 filter=137 channel=53
    -5, -3, -14, -9, 6, -5, 5, -7, -4,
    -- layer=1 filter=137 channel=54
    46, -14, -7, 2, -11, -37, -9, -3, 16,
    -- layer=1 filter=137 channel=55
    29, 4, 17, 12, -2, 0, 9, 18, -7,
    -- layer=1 filter=137 channel=56
    -8, 4, -3, 0, 8, -3, 0, -9, -11,
    -- layer=1 filter=137 channel=57
    22, -56, -23, 27, -35, -19, -47, -15, -19,
    -- layer=1 filter=137 channel=58
    57, -72, 2, 20, -49, -32, -22, -54, -36,
    -- layer=1 filter=137 channel=59
    8, -2, -5, -9, -6, -2, -13, 1, 9,
    -- layer=1 filter=137 channel=60
    5, -38, -31, -26, -5, -34, 0, 11, -29,
    -- layer=1 filter=137 channel=61
    -10, -8, 4, -2, -3, 6, 2, 3, -7,
    -- layer=1 filter=137 channel=62
    44, -34, -57, 25, -79, -68, -28, -50, -30,
    -- layer=1 filter=137 channel=63
    -29, -58, -23, -17, -29, -33, -7, 24, -32,
    -- layer=1 filter=137 channel=64
    -13, -7, -45, 10, -4, -27, 23, -1, -14,
    -- layer=1 filter=137 channel=65
    -15, -47, -50, -17, -38, -54, 1, -69, -71,
    -- layer=1 filter=137 channel=66
    -37, -57, -33, -10, -24, -31, -2, -33, -31,
    -- layer=1 filter=137 channel=67
    -62, -43, -44, -11, -39, -74, -79, -23, -61,
    -- layer=1 filter=137 channel=68
    18, -68, -107, 59, -10, -63, 72, 26, -76,
    -- layer=1 filter=137 channel=69
    72, 19, 2, 83, -16, 2, 43, 26, -26,
    -- layer=1 filter=137 channel=70
    -35, -57, -43, -9, -20, -44, 3, 19, -18,
    -- layer=1 filter=137 channel=71
    11, 10, -16, -1, -13, -28, -19, -23, -7,
    -- layer=1 filter=137 channel=72
    -40, -61, -25, -18, -5, -44, -29, -7, -12,
    -- layer=1 filter=137 channel=73
    -4, 3, 5, -5, -7, -9, -9, 12, -9,
    -- layer=1 filter=137 channel=74
    -1, -44, -18, 13, -24, -79, 39, 21, -53,
    -- layer=1 filter=137 channel=75
    7, 15, 25, 10, -17, 51, -22, 10, -26,
    -- layer=1 filter=137 channel=76
    -23, -105, -63, 14, -42, -48, 35, 49, -14,
    -- layer=1 filter=137 channel=77
    12, -27, -44, 30, -23, -56, 27, -57, -38,
    -- layer=1 filter=137 channel=78
    5, -2, -18, 10, -6, -20, -14, -11, -21,
    -- layer=1 filter=137 channel=79
    57, -24, -34, 9, -44, -56, -29, -11, -23,
    -- layer=1 filter=137 channel=80
    -6, 15, 6, -12, 6, 8, 5, -13, 13,
    -- layer=1 filter=137 channel=81
    -2, -19, -45, 0, -27, -46, -28, -18, -40,
    -- layer=1 filter=137 channel=82
    -25, -30, -55, 13, -32, -36, -18, -21, -45,
    -- layer=1 filter=137 channel=83
    43, -8, -11, 98, 22, -38, 56, 20, -34,
    -- layer=1 filter=137 channel=84
    -41, -110, -70, -12, -44, -92, 39, 36, -35,
    -- layer=1 filter=137 channel=85
    65, -40, 2, 49, -44, 3, 48, 17, 15,
    -- layer=1 filter=137 channel=86
    -29, -42, -13, -7, -34, -30, -13, -35, -35,
    -- layer=1 filter=137 channel=87
    -6, 9, 23, -22, 45, -18, -27, 19, 50,
    -- layer=1 filter=137 channel=88
    -7, -1, 0, -9, 15, 10, -33, -1, -2,
    -- layer=1 filter=137 channel=89
    -1, -30, -60, 37, -7, -37, 11, 12, -46,
    -- layer=1 filter=137 channel=90
    27, -79, -97, 54, -36, -64, 67, 29, -60,
    -- layer=1 filter=137 channel=91
    -20, -43, -48, -18, -48, -50, -8, -62, -52,
    -- layer=1 filter=137 channel=92
    75, -25, 2, 103, 40, 45, 81, 90, -12,
    -- layer=1 filter=137 channel=93
    -24, -32, -70, 5, -50, -52, -2, -47, -66,
    -- layer=1 filter=137 channel=94
    -47, -52, -15, -12, -33, -61, 14, -16, -57,
    -- layer=1 filter=137 channel=95
    -50, -110, -48, -72, -55, -62, -4, -23, -86,
    -- layer=1 filter=137 channel=96
    5, 19, 2, 27, 13, 28, -14, 9, 9,
    -- layer=1 filter=137 channel=97
    -30, -54, -63, 2, -39, -60, 6, -55, -72,
    -- layer=1 filter=137 channel=98
    16, -39, -79, 4, -101, -67, -50, -69, -56,
    -- layer=1 filter=137 channel=99
    12, -52, -30, 10, -49, -51, 21, -52, -36,
    -- layer=1 filter=137 channel=100
    -21, -44, -9, -17, -20, -27, 12, 13, -32,
    -- layer=1 filter=137 channel=101
    -34, -47, -52, -11, -35, -48, 9, -25, -48,
    -- layer=1 filter=137 channel=102
    -92, -59, -22, -27, -31, -62, 13, -27, -71,
    -- layer=1 filter=137 channel=103
    -27, -24, -19, -44, -33, -6, 8, -2, 18,
    -- layer=1 filter=137 channel=104
    21, -46, 10, 45, 0, 14, 49, 24, -23,
    -- layer=1 filter=137 channel=105
    -65, -73, -57, 0, -48, -69, 30, -67, -49,
    -- layer=1 filter=137 channel=106
    19, -57, -58, 39, -1, -32, 60, 42, -49,
    -- layer=1 filter=137 channel=107
    0, -5, 2, 7, -7, -2, 6, 8, -5,
    -- layer=1 filter=137 channel=108
    38, -60, -69, 50, 2, -34, 59, 64, -49,
    -- layer=1 filter=137 channel=109
    -3, 3, 11, -9, -2, -8, 5, -1, -7,
    -- layer=1 filter=137 channel=110
    -1, 0, 11, -7, -2, -2, 5, 4, -20,
    -- layer=1 filter=137 channel=111
    -85, -99, -39, -116, -54, -75, -33, -15, -42,
    -- layer=1 filter=137 channel=112
    -22, -51, -53, -26, 0, -5, 19, 6, -13,
    -- layer=1 filter=137 channel=113
    32, 52, 30, 29, 34, 61, 10, 52, 63,
    -- layer=1 filter=137 channel=114
    60, 25, 10, 48, -10, -15, 24, -9, -3,
    -- layer=1 filter=137 channel=115
    -20, -49, -25, 5, -60, -50, -11, -48, -18,
    -- layer=1 filter=137 channel=116
    9, -6, 0, -4, -4, 7, -8, 0, 1,
    -- layer=1 filter=137 channel=117
    8, -69, -58, -21, -60, -34, 0, -6, -13,
    -- layer=1 filter=137 channel=118
    -62, -90, -61, -23, -66, -99, 31, -22, -31,
    -- layer=1 filter=137 channel=119
    26, -87, -88, 43, -5, -62, 49, 62, -50,
    -- layer=1 filter=137 channel=120
    27, -20, -14, -18, -20, -22, -60, -29, -34,
    -- layer=1 filter=137 channel=121
    -14, -13, 28, -36, 9, 14, -45, 8, 12,
    -- layer=1 filter=137 channel=122
    -9, 6, -3, 2, 0, 6, 7, -6, -1,
    -- layer=1 filter=137 channel=123
    7, 6, 16, -17, 20, 0, -48, -8, 9,
    -- layer=1 filter=137 channel=124
    25, 31, 42, 30, 16, 17, 28, 20, 33,
    -- layer=1 filter=137 channel=125
    -4, -11, 19, 16, 10, -23, 22, -33, 27,
    -- layer=1 filter=137 channel=126
    -3, 31, -76, 59, -59, -37, 14, -25, -33,
    -- layer=1 filter=137 channel=127
    -88, -94, -34, -84, -84, -71, -27, -7, -64,
    -- layer=1 filter=138 channel=0
    -27, -54, -52, 34, 11, -3, -10, -27, -40,
    -- layer=1 filter=138 channel=1
    37, 49, 27, -14, -91, -78, -35, 37, 54,
    -- layer=1 filter=138 channel=2
    40, 38, 60, 44, 69, 86, 42, -33, -45,
    -- layer=1 filter=138 channel=3
    -11, -3, -2, 3, -4, -6, -7, 7, -7,
    -- layer=1 filter=138 channel=4
    14, 0, 15, 7, 17, 6, 0, -1, -7,
    -- layer=1 filter=138 channel=5
    77, 58, 40, -44, -95, -64, -14, 60, 73,
    -- layer=1 filter=138 channel=6
    -95, -36, -48, -83, -66, -46, -37, -45, -11,
    -- layer=1 filter=138 channel=7
    -23, 30, -54, -39, -45, -48, 14, 14, -23,
    -- layer=1 filter=138 channel=8
    68, 62, 23, -68, -126, -82, -11, 47, 63,
    -- layer=1 filter=138 channel=9
    78, 11, 17, 69, 57, 37, -12, -29, -75,
    -- layer=1 filter=138 channel=10
    -37, 13, -53, -28, -56, -66, 15, 34, -18,
    -- layer=1 filter=138 channel=11
    -7, -57, -32, 30, -12, 11, -3, -44, -42,
    -- layer=1 filter=138 channel=12
    -21, 10, 8, 12, 29, 39, 1, -60, -55,
    -- layer=1 filter=138 channel=13
    19, -23, -44, -14, -35, -52, 0, -14, 15,
    -- layer=1 filter=138 channel=14
    -13, 29, -19, 7, -12, 14, -6, -116, -63,
    -- layer=1 filter=138 channel=15
    60, 39, 34, 5, -12, -12, 11, 49, 102,
    -- layer=1 filter=138 channel=16
    53, 52, 25, -97, -101, -76, 8, 45, 76,
    -- layer=1 filter=138 channel=17
    -3, -27, -29, -12, -33, -33, 16, -9, -10,
    -- layer=1 filter=138 channel=18
    -82, -76, -36, 2, 1, 25, -33, -92, -57,
    -- layer=1 filter=138 channel=19
    0, -22, -38, -14, -46, -41, 45, 73, 23,
    -- layer=1 filter=138 channel=20
    -48, -31, -52, -65, -122, -136, -27, -2, 10,
    -- layer=1 filter=138 channel=21
    7, 13, -26, -14, -18, -56, -45, -24, -13,
    -- layer=1 filter=138 channel=22
    31, 22, 0, -39, -91, -109, -33, 20, 49,
    -- layer=1 filter=138 channel=23
    27, 33, 15, -8, 57, -16, -53, -9, 4,
    -- layer=1 filter=138 channel=24
    54, 4, 0, 10, -15, -5, 16, 39, 52,
    -- layer=1 filter=138 channel=25
    0, 32, 0, -66, -55, -53, 14, 57, 37,
    -- layer=1 filter=138 channel=26
    53, -19, 6, 8, 11, 2, 16, -26, 32,
    -- layer=1 filter=138 channel=27
    -49, -29, -24, -58, -45, -26, -46, -49, -56,
    -- layer=1 filter=138 channel=28
    -6, 35, -25, 5, -26, -51, -12, 36, 2,
    -- layer=1 filter=138 channel=29
    -27, -27, -25, -26, -40, -7, -10, 11, 10,
    -- layer=1 filter=138 channel=30
    -31, -75, -57, -16, -25, -28, -2, -36, -56,
    -- layer=1 filter=138 channel=31
    -84, -16, 13, -18, -1, 40, -12, -78, -48,
    -- layer=1 filter=138 channel=32
    34, -10, 9, 31, 25, -5, -23, -13, -35,
    -- layer=1 filter=138 channel=33
    32, 23, 24, 58, 57, 35, 19, 8, 9,
    -- layer=1 filter=138 channel=34
    -19, 8, -10, 1, 24, 24, 10, 23, 5,
    -- layer=1 filter=138 channel=35
    -7, -8, -17, -6, 3, -4, 18, 1, 19,
    -- layer=1 filter=138 channel=36
    -22, -70, -43, 19, -29, -18, 7, -35, -51,
    -- layer=1 filter=138 channel=37
    79, 47, 35, -79, -95, -54, 2, 53, 72,
    -- layer=1 filter=138 channel=38
    -51, -39, -55, -27, -51, -57, -37, -10, -16,
    -- layer=1 filter=138 channel=39
    37, 12, 16, -34, -16, -7, 5, 48, 59,
    -- layer=1 filter=138 channel=40
    -106, -26, -47, -42, -14, 3, 8, -74, -45,
    -- layer=1 filter=138 channel=41
    59, -12, 7, 21, 62, 32, 0, -23, -12,
    -- layer=1 filter=138 channel=42
    27, 33, 54, 31, 59, 81, 55, -11, -36,
    -- layer=1 filter=138 channel=43
    49, 42, 1, -72, -113, -51, -19, 48, 51,
    -- layer=1 filter=138 channel=44
    51, -9, -13, 48, -12, 15, -24, -26, 35,
    -- layer=1 filter=138 channel=45
    45, -1, -5, -13, -65, -30, -23, 6, 51,
    -- layer=1 filter=138 channel=46
    13, -12, -25, -55, -30, -19, -11, 54, 35,
    -- layer=1 filter=138 channel=47
    70, 46, 75, 27, 61, 26, -28, -62, -6,
    -- layer=1 filter=138 channel=48
    -49, -64, -85, -55, -63, -102, -59, -58, -67,
    -- layer=1 filter=138 channel=49
    26, 10, 15, 9, 50, 25, 24, 1, -43,
    -- layer=1 filter=138 channel=50
    4, -3, -20, 38, -33, 10, -13, 2, -6,
    -- layer=1 filter=138 channel=51
    -33, -25, -69, -32, -38, -65, -20, -37, -59,
    -- layer=1 filter=138 channel=52
    6, 22, 38, 17, 41, 28, -5, 10, 3,
    -- layer=1 filter=138 channel=53
    -1, 1, 22, 14, 1, 6, -1, 11, 12,
    -- layer=1 filter=138 channel=54
    35, 30, 4, -27, -63, -39, 22, 75, 62,
    -- layer=1 filter=138 channel=55
    32, 28, 24, 0, 7, 13, 4, 5, 39,
    -- layer=1 filter=138 channel=56
    -9, -4, 6, -11, 3, 0, -3, -2, 3,
    -- layer=1 filter=138 channel=57
    -22, 1, -29, -51, -71, -57, 0, 27, -8,
    -- layer=1 filter=138 channel=58
    15, -8, -8, -40, -9, -37, -6, 24, 5,
    -- layer=1 filter=138 channel=59
    -7, 2, 3, 0, -1, 4, -5, 9, 12,
    -- layer=1 filter=138 channel=60
    14, -36, -16, -14, -3, -8, 4, -9, -18,
    -- layer=1 filter=138 channel=61
    -6, -4, -7, 9, 7, -3, 8, -10, 8,
    -- layer=1 filter=138 channel=62
    55, 39, 0, -73, -115, -57, 14, 56, 56,
    -- layer=1 filter=138 channel=63
    -48, -58, -42, 9, -10, 2, -35, -39, -37,
    -- layer=1 filter=138 channel=64
    -66, -33, -33, 2, -47, -53, -28, -7, -42,
    -- layer=1 filter=138 channel=65
    -64, -37, -77, -43, -61, -86, -74, -57, -53,
    -- layer=1 filter=138 channel=66
    -33, -43, -41, -1, -40, -37, -34, -32, -47,
    -- layer=1 filter=138 channel=67
    -9, -20, -23, 4, -12, 17, 0, 8, 31,
    -- layer=1 filter=138 channel=68
    49, -10, -25, 41, -3, 36, -12, -42, 35,
    -- layer=1 filter=138 channel=69
    82, 42, 38, -11, -30, -35, 0, 63, 95,
    -- layer=1 filter=138 channel=70
    -47, -13, -17, -34, -1, 7, 51, 24, 16,
    -- layer=1 filter=138 channel=71
    -22, 2, -14, -53, -37, -46, -24, 30, 11,
    -- layer=1 filter=138 channel=72
    -14, -31, -29, 0, -17, -27, 23, 21, -70,
    -- layer=1 filter=138 channel=73
    9, 7, -10, -8, -11, 1, 0, 1, -1,
    -- layer=1 filter=138 channel=74
    -41, -63, -30, 7, -27, 22, 16, -15, -8,
    -- layer=1 filter=138 channel=75
    -57, -33, -10, -17, -10, 25, -11, -99, -73,
    -- layer=1 filter=138 channel=76
    16, -63, -57, 12, -9, -16, -2, -20, -5,
    -- layer=1 filter=138 channel=77
    -10, -24, -25, -27, -34, -48, -51, 11, -1,
    -- layer=1 filter=138 channel=78
    -16, -13, -11, 20, -21, -10, 14, 0, -4,
    -- layer=1 filter=138 channel=79
    56, 36, 14, -97, -98, -74, 13, 59, 69,
    -- layer=1 filter=138 channel=80
    -55, 9, 2, 6, 1, -4, -37, -2, -26,
    -- layer=1 filter=138 channel=81
    37, 19, 3, -37, -48, -54, -13, 33, 48,
    -- layer=1 filter=138 channel=82
    -11, -23, -41, -15, -36, -45, -60, -22, -36,
    -- layer=1 filter=138 channel=83
    52, 44, 5, 3, -66, -28, -19, 25, 63,
    -- layer=1 filter=138 channel=84
    -7, -71, -30, 7, 27, 11, -75, -32, -18,
    -- layer=1 filter=138 channel=85
    10, 2, 3, 3, 28, 16, -9, 44, -16,
    -- layer=1 filter=138 channel=86
    -33, -13, -24, -42, -66, -65, -15, 7, 10,
    -- layer=1 filter=138 channel=87
    34, 19, 9, 38, 6, -10, 46, 83, -22,
    -- layer=1 filter=138 channel=88
    15, 10, -19, 3, 9, -4, 3, -5, -39,
    -- layer=1 filter=138 channel=89
    -29, -43, -58, -1, -9, -25, -70, -47, -47,
    -- layer=1 filter=138 channel=90
    40, -3, -14, 19, -7, 11, 4, -22, 27,
    -- layer=1 filter=138 channel=91
    -100, -71, -64, -81, -52, -91, -57, -90, -111,
    -- layer=1 filter=138 channel=92
    65, 60, 26, 51, 48, 12, -37, 16, -20,
    -- layer=1 filter=138 channel=93
    -14, -28, -66, -34, -86, -87, -50, -9, -10,
    -- layer=1 filter=138 channel=94
    -64, -51, -52, -2, -6, -17, -10, -23, -56,
    -- layer=1 filter=138 channel=95
    -51, -63, -47, 6, -12, 1, -32, -55, -29,
    -- layer=1 filter=138 channel=96
    -1, 6, -11, 35, 28, 11, -11, -6, -34,
    -- layer=1 filter=138 channel=97
    -34, -62, -72, -28, -76, -80, -31, -9, -16,
    -- layer=1 filter=138 channel=98
    65, 36, 12, -64, -112, -70, -2, 67, 65,
    -- layer=1 filter=138 channel=99
    -1, 5, -8, 72, 0, -5, 36, 0, 7,
    -- layer=1 filter=138 channel=100
    -16, -49, -38, 0, -15, -24, -30, -29, -37,
    -- layer=1 filter=138 channel=101
    -93, -80, -90, -30, -58, -93, -101, -83, -83,
    -- layer=1 filter=138 channel=102
    -83, -78, -47, -34, -22, -43, -3, -21, -12,
    -- layer=1 filter=138 channel=103
    -38, -73, -33, 38, 9, -4, -39, -33, -35,
    -- layer=1 filter=138 channel=104
    24, -5, 20, 33, 49, -12, -66, -24, -11,
    -- layer=1 filter=138 channel=105
    -72, -68, -71, -28, -48, -69, -31, -33, -71,
    -- layer=1 filter=138 channel=106
    -14, -35, -46, 12, -22, -22, -56, -43, -31,
    -- layer=1 filter=138 channel=107
    0, -5, 0, -2, 4, -9, -12, 0, 2,
    -- layer=1 filter=138 channel=108
    58, 34, 9, 40, 11, 4, 13, -7, 48,
    -- layer=1 filter=138 channel=109
    -3, 8, 5, 0, 6, -8, 8, -8, 0,
    -- layer=1 filter=138 channel=110
    -19, 3, -22, -29, -17, -17, -22, -9, -21,
    -- layer=1 filter=138 channel=111
    -60, -84, -75, -12, -17, 2, -26, -83, -34,
    -- layer=1 filter=138 channel=112
    -47, -45, -43, 24, 21, 18, -74, -17, -14,
    -- layer=1 filter=138 channel=113
    24, 39, 38, 1, 29, 50, 17, 30, 10,
    -- layer=1 filter=138 channel=114
    80, 62, 32, -71, -99, -57, -11, 65, 89,
    -- layer=1 filter=138 channel=115
    -71, -18, -53, -66, -63, -64, -24, 4, -33,
    -- layer=1 filter=138 channel=116
    -4, -8, -8, -4, -4, -4, -1, -9, -9,
    -- layer=1 filter=138 channel=117
    -84, -32, -63, 10, 8, 7, -77, -83, -57,
    -- layer=1 filter=138 channel=118
    -35, -78, -56, 20, 2, 8, -16, -39, -43,
    -- layer=1 filter=138 channel=119
    36, -3, -16, 13, 21, 11, 10, -27, 2,
    -- layer=1 filter=138 channel=120
    -2, 23, -17, -38, -37, -54, -6, 37, 16,
    -- layer=1 filter=138 channel=121
    -53, -27, -20, -25, -32, -14, 6, -14, -89,
    -- layer=1 filter=138 channel=122
    -5, 9, -2, -6, 5, 3, -10, 5, -3,
    -- layer=1 filter=138 channel=123
    -49, -31, -2, -23, -3, 6, -16, -32, -53,
    -- layer=1 filter=138 channel=124
    5, -1, -8, 6, -16, -22, 2, -4, -10,
    -- layer=1 filter=138 channel=125
    -28, 6, -25, -42, -28, -27, 12, 12, -30,
    -- layer=1 filter=138 channel=126
    57, 25, -5, -27, -104, -79, -14, 38, 25,
    -- layer=1 filter=138 channel=127
    -60, -82, -59, -13, 8, 25, -11, -58, -43,
    -- layer=1 filter=139 channel=0
    -18, -30, -18, -5, -7, -5, -12, -1, -9,
    -- layer=1 filter=139 channel=1
    1, 25, 18, -7, -10, -4, 3, 2, 7,
    -- layer=1 filter=139 channel=2
    -35, -29, -20, 6, -8, -13, -2, -3, -6,
    -- layer=1 filter=139 channel=3
    6, 4, 8, 8, 7, -4, -8, -1, 2,
    -- layer=1 filter=139 channel=4
    7, 3, 9, -10, -8, -3, -1, 2, -3,
    -- layer=1 filter=139 channel=5
    12, 31, 15, 1, -9, -6, -24, -14, -28,
    -- layer=1 filter=139 channel=6
    -10, -13, -6, -30, -20, -12, -22, -24, -12,
    -- layer=1 filter=139 channel=7
    -5, -10, -8, -9, -9, -10, 5, -16, 2,
    -- layer=1 filter=139 channel=8
    17, 25, 12, 0, 3, 4, 2, -5, -21,
    -- layer=1 filter=139 channel=9
    -14, 0, -10, -22, -16, 4, -19, 2, 7,
    -- layer=1 filter=139 channel=10
    3, -11, -2, -16, 0, -10, -9, -14, -1,
    -- layer=1 filter=139 channel=11
    -14, -15, -19, -22, -31, -17, 1, -18, -23,
    -- layer=1 filter=139 channel=12
    4, 4, -14, -7, -32, 6, 0, -26, -27,
    -- layer=1 filter=139 channel=13
    0, -6, 8, -21, 0, -2, -11, -19, -6,
    -- layer=1 filter=139 channel=14
    -8, -12, -19, -11, -9, -20, -26, -2, -21,
    -- layer=1 filter=139 channel=15
    9, 16, 10, -22, -21, 7, -7, -15, 9,
    -- layer=1 filter=139 channel=16
    22, 28, 15, 3, -2, -8, -8, -15, -14,
    -- layer=1 filter=139 channel=17
    -28, -29, -9, -13, -17, -16, -15, 0, 1,
    -- layer=1 filter=139 channel=18
    -2, 5, 4, -17, -27, -7, 4, -30, -21,
    -- layer=1 filter=139 channel=19
    -1, 4, -16, -16, -16, 3, -23, 0, -10,
    -- layer=1 filter=139 channel=20
    -8, -5, 4, -1, -10, 1, -24, -13, -4,
    -- layer=1 filter=139 channel=21
    2, -14, -8, -3, -14, -17, -24, -9, -23,
    -- layer=1 filter=139 channel=22
    -2, 3, 27, 0, -9, 3, -24, -6, -5,
    -- layer=1 filter=139 channel=23
    -11, 2, 4, -6, -12, 7, 1, -44, -1,
    -- layer=1 filter=139 channel=24
    -3, -15, -13, -19, -18, -15, -17, -3, -21,
    -- layer=1 filter=139 channel=25
    16, 12, 13, 3, -12, 2, 0, -24, 8,
    -- layer=1 filter=139 channel=26
    -16, -16, -17, -12, -14, -15, -14, -6, 5,
    -- layer=1 filter=139 channel=27
    -37, -25, -23, -31, -25, -29, -10, -5, 13,
    -- layer=1 filter=139 channel=28
    0, -14, 2, -5, 0, -11, -11, -23, -1,
    -- layer=1 filter=139 channel=29
    -15, -14, -13, 0, 0, -12, -1, 3, -9,
    -- layer=1 filter=139 channel=30
    1, -7, -2, -22, -12, -14, -22, -14, -19,
    -- layer=1 filter=139 channel=31
    -1, -16, -26, -20, -24, 13, -25, -35, -38,
    -- layer=1 filter=139 channel=32
    -31, -14, -32, -13, -3, -9, -13, -17, -4,
    -- layer=1 filter=139 channel=33
    1, 0, -20, -10, -12, -6, -5, -15, 0,
    -- layer=1 filter=139 channel=34
    4, 6, -6, 2, -2, -1, -10, -7, -1,
    -- layer=1 filter=139 channel=35
    3, -1, 2, 1, 9, -10, 5, -1, 1,
    -- layer=1 filter=139 channel=36
    -28, -38, -31, -39, -33, -7, -16, -3, -16,
    -- layer=1 filter=139 channel=37
    32, 34, 12, 0, -10, -2, 4, -10, -30,
    -- layer=1 filter=139 channel=38
    -17, -17, -13, -21, 6, -3, -10, -11, -9,
    -- layer=1 filter=139 channel=39
    -11, 0, 4, 9, 1, 2, 13, 10, 8,
    -- layer=1 filter=139 channel=40
    3, 0, -3, -25, -21, -5, -12, -31, -17,
    -- layer=1 filter=139 channel=41
    -20, -2, -11, -7, -28, 9, -10, -17, 2,
    -- layer=1 filter=139 channel=42
    -34, -23, -12, -9, -10, -4, -17, -11, -9,
    -- layer=1 filter=139 channel=43
    16, 28, 12, -7, -6, 7, -4, -7, -3,
    -- layer=1 filter=139 channel=44
    -17, -17, -20, -23, -3, -21, -33, -1, -5,
    -- layer=1 filter=139 channel=45
    -7, 20, 6, -23, -5, -8, -12, -23, -14,
    -- layer=1 filter=139 channel=46
    18, 30, -6, 0, 0, 5, -19, -2, -10,
    -- layer=1 filter=139 channel=47
    -8, -23, 19, 8, -19, 15, -23, -22, 13,
    -- layer=1 filter=139 channel=48
    -14, -19, -24, 1, -7, -8, 5, -6, -4,
    -- layer=1 filter=139 channel=49
    -17, -22, -21, -13, -28, -9, -25, -17, -6,
    -- layer=1 filter=139 channel=50
    -7, 4, 6, 3, -4, -14, -9, -6, -20,
    -- layer=1 filter=139 channel=51
    -24, -7, -15, -16, -18, -12, -8, -2, -4,
    -- layer=1 filter=139 channel=52
    -12, 7, 1, -6, -1, -5, -10, -5, -1,
    -- layer=1 filter=139 channel=53
    3, -5, -10, -2, 4, 3, 8, -5, -5,
    -- layer=1 filter=139 channel=54
    22, 29, 5, -8, -10, 13, -1, -20, -10,
    -- layer=1 filter=139 channel=55
    -16, -4, -14, -17, -30, -10, -22, -16, -16,
    -- layer=1 filter=139 channel=56
    -5, 6, 8, -1, 4, 6, -5, -11, -8,
    -- layer=1 filter=139 channel=57
    -9, -3, 2, -13, -5, -12, -5, -29, -10,
    -- layer=1 filter=139 channel=58
    -13, -12, 0, 6, -20, 13, 5, -19, -5,
    -- layer=1 filter=139 channel=59
    4, 2, 7, 2, -9, -4, -10, 6, -11,
    -- layer=1 filter=139 channel=60
    -6, -2, -11, -2, 8, 6, 0, 15, -3,
    -- layer=1 filter=139 channel=61
    -5, -1, -1, 1, 3, 10, -9, -5, 0,
    -- layer=1 filter=139 channel=62
    26, 34, 10, 0, -10, 11, 8, -14, -13,
    -- layer=1 filter=139 channel=63
    -21, -18, -13, -40, -35, -21, -11, -18, -15,
    -- layer=1 filter=139 channel=64
    -18, -5, 14, 7, -2, 4, -4, 3, 4,
    -- layer=1 filter=139 channel=65
    -13, 0, 0, -13, -8, -15, -11, -2, 8,
    -- layer=1 filter=139 channel=66
    -28, -12, -14, -20, -11, -15, -4, -12, -4,
    -- layer=1 filter=139 channel=67
    -14, -24, -16, -12, -4, 0, -6, -4, 6,
    -- layer=1 filter=139 channel=68
    -23, -11, -18, -30, -4, -15, -9, 4, 3,
    -- layer=1 filter=139 channel=69
    28, 40, 10, -18, -19, -9, -28, -15, -11,
    -- layer=1 filter=139 channel=70
    -11, -3, -36, -3, -7, -5, 4, -10, -9,
    -- layer=1 filter=139 channel=71
    -5, -14, -14, -20, -10, -13, -5, -13, -31,
    -- layer=1 filter=139 channel=72
    -12, -4, -8, -26, -11, -7, -24, 0, -1,
    -- layer=1 filter=139 channel=73
    2, 0, 1, 5, 8, 7, 7, -1, 3,
    -- layer=1 filter=139 channel=74
    -6, 0, -14, -9, -5, 5, -14, -9, -38,
    -- layer=1 filter=139 channel=75
    22, -6, -27, -13, -11, 11, -13, -21, -21,
    -- layer=1 filter=139 channel=76
    -11, 2, 0, -6, -6, 5, -11, -6, -11,
    -- layer=1 filter=139 channel=77
    6, -7, -17, -10, 4, -6, -13, -11, -3,
    -- layer=1 filter=139 channel=78
    5, -14, -19, -27, -11, -7, -6, -14, -14,
    -- layer=1 filter=139 channel=79
    16, 10, 19, -8, -15, 11, -14, -8, -29,
    -- layer=1 filter=139 channel=80
    10, -3, -3, 0, 0, 0, -2, -8, -9,
    -- layer=1 filter=139 channel=81
    0, -7, -2, -9, 0, -16, 0, -15, -4,
    -- layer=1 filter=139 channel=82
    -20, -16, -23, 9, -10, -2, -14, 1, -9,
    -- layer=1 filter=139 channel=83
    -1, 3, 2, -6, 2, 1, -26, 2, -14,
    -- layer=1 filter=139 channel=84
    2, 0, 12, -17, -15, -23, -4, -16, -21,
    -- layer=1 filter=139 channel=85
    5, 3, 29, -4, -28, 15, 15, -22, -3,
    -- layer=1 filter=139 channel=86
    -14, -20, -5, -3, -8, -2, -9, -16, -8,
    -- layer=1 filter=139 channel=87
    16, 1, -13, -27, -6, 1, -17, -18, 12,
    -- layer=1 filter=139 channel=88
    -38, -27, -31, -23, -18, -18, -5, 2, -17,
    -- layer=1 filter=139 channel=89
    -14, -13, -16, -24, -10, -33, -10, -4, -19,
    -- layer=1 filter=139 channel=90
    -17, -10, -17, -28, -9, -17, -13, -7, -10,
    -- layer=1 filter=139 channel=91
    -17, -7, -6, 0, -17, -5, -18, -1, 2,
    -- layer=1 filter=139 channel=92
    -32, -25, 3, -8, -2, -2, 0, 12, 5,
    -- layer=1 filter=139 channel=93
    -7, -10, -21, -2, -4, -10, -15, 2, -8,
    -- layer=1 filter=139 channel=94
    -20, -19, -9, -13, -19, -9, -10, -12, 0,
    -- layer=1 filter=139 channel=95
    -4, -1, -8, -16, -29, -4, -16, -17, -17,
    -- layer=1 filter=139 channel=96
    3, 3, 6, -7, -7, -9, -1, -8, 3,
    -- layer=1 filter=139 channel=97
    -12, -16, -10, -6, -7, -22, -10, -11, 2,
    -- layer=1 filter=139 channel=98
    25, 22, 27, 16, 2, -7, 17, 6, -2,
    -- layer=1 filter=139 channel=99
    -3, -4, -3, -23, -9, -23, -26, -7, -9,
    -- layer=1 filter=139 channel=100
    -22, -12, -17, -19, -25, -24, -22, -25, -20,
    -- layer=1 filter=139 channel=101
    -16, -20, -22, -12, -15, -24, -21, -4, -18,
    -- layer=1 filter=139 channel=102
    -8, -9, -12, -6, -12, 4, 5, 7, 2,
    -- layer=1 filter=139 channel=103
    -1, -3, 7, -30, -38, -41, -20, -29, -38,
    -- layer=1 filter=139 channel=104
    -5, -1, -13, -1, -4, 5, 11, -13, 15,
    -- layer=1 filter=139 channel=105
    -22, -26, -24, -4, -9, -6, -3, -11, -16,
    -- layer=1 filter=139 channel=106
    -30, -15, -19, -32, -10, -30, -12, -20, -6,
    -- layer=1 filter=139 channel=107
    5, -3, -9, 5, 5, 10, -10, -11, -1,
    -- layer=1 filter=139 channel=108
    -19, -22, -7, -20, -5, -6, -23, 0, -3,
    -- layer=1 filter=139 channel=109
    10, -1, -10, -4, 2, 1, -6, 0, -1,
    -- layer=1 filter=139 channel=110
    2, 0, -2, 6, -8, -9, -11, -8, 7,
    -- layer=1 filter=139 channel=111
    14, 1, 4, -29, -28, -20, -2, -17, -23,
    -- layer=1 filter=139 channel=112
    -5, -3, 2, -10, -6, -9, -5, -20, -35,
    -- layer=1 filter=139 channel=113
    -3, -1, -20, -13, -7, -27, -8, -24, -12,
    -- layer=1 filter=139 channel=114
    27, 26, 11, -10, -12, -14, -1, -7, -31,
    -- layer=1 filter=139 channel=115
    -10, -7, -7, 0, -20, -14, -9, -12, -1,
    -- layer=1 filter=139 channel=116
    -7, 0, 6, -9, 0, 9, -8, 0, 4,
    -- layer=1 filter=139 channel=117
    0, 16, 10, -10, -15, -25, -4, -16, -18,
    -- layer=1 filter=139 channel=118
    8, 0, 1, -12, -7, -15, -7, -24, -33,
    -- layer=1 filter=139 channel=119
    -32, -26, -21, -20, -12, -8, -16, 0, -6,
    -- layer=1 filter=139 channel=120
    0, 7, -5, -10, -10, -17, -10, -12, -20,
    -- layer=1 filter=139 channel=121
    7, -18, -16, -18, -6, -4, -37, -11, -15,
    -- layer=1 filter=139 channel=122
    -3, -4, 4, -4, 8, 3, 5, 5, -6,
    -- layer=1 filter=139 channel=123
    -21, -25, -22, -14, -29, -24, -22, -34, -20,
    -- layer=1 filter=139 channel=124
    -2, 7, 5, 2, 2, 6, -6, -7, -10,
    -- layer=1 filter=139 channel=125
    0, -2, -29, -12, -14, -17, -12, -24, -27,
    -- layer=1 filter=139 channel=126
    -7, 0, -3, 6, -8, -1, 13, 7, -7,
    -- layer=1 filter=139 channel=127
    16, -4, -2, -10, -8, -2, -7, -23, -16,
    -- layer=1 filter=140 channel=0
    2, 2, -2, -10, 1, -1, -19, 9, -4,
    -- layer=1 filter=140 channel=1
    -4, -6, -6, -10, -6, -1, -5, -11, -14,
    -- layer=1 filter=140 channel=2
    0, 0, 0, -3, -7, 6, -4, 1, 0,
    -- layer=1 filter=140 channel=3
    -1, -4, 8, 3, 2, 5, 0, 1, -8,
    -- layer=1 filter=140 channel=4
    -10, 3, 6, 0, 8, -10, -1, 0, 6,
    -- layer=1 filter=140 channel=5
    -3, 4, 2, -4, -4, 9, 1, -11, -4,
    -- layer=1 filter=140 channel=6
    -12, 1, -9, 4, -9, -11, -12, -5, -8,
    -- layer=1 filter=140 channel=7
    0, 4, -3, 1, 15, 5, -16, 16, 0,
    -- layer=1 filter=140 channel=8
    -12, 2, -11, 6, -6, -1, -8, 2, -10,
    -- layer=1 filter=140 channel=9
    0, -7, -8, -13, -11, -2, 14, -6, 1,
    -- layer=1 filter=140 channel=10
    -12, -7, -6, -10, 3, -6, -4, 6, -7,
    -- layer=1 filter=140 channel=11
    -13, 10, -5, 2, -4, -14, 12, -7, -2,
    -- layer=1 filter=140 channel=12
    -2, 7, -1, 2, 0, 3, 1, 1, -4,
    -- layer=1 filter=140 channel=13
    -7, -9, 0, -15, 0, -12, 3, -3, -12,
    -- layer=1 filter=140 channel=14
    4, -1, -8, -9, 4, -4, 8, -4, 2,
    -- layer=1 filter=140 channel=15
    2, 2, 14, 12, -7, 0, -15, -8, -3,
    -- layer=1 filter=140 channel=16
    4, 3, 4, -2, -2, -11, -14, -4, -4,
    -- layer=1 filter=140 channel=17
    0, 10, -7, -1, -3, -10, -15, -2, -6,
    -- layer=1 filter=140 channel=18
    -2, -17, 3, -2, 15, -2, -1, -12, 3,
    -- layer=1 filter=140 channel=19
    -14, -18, -11, 0, 2, 6, -10, -14, -3,
    -- layer=1 filter=140 channel=20
    -17, 0, -2, -10, -9, -8, -5, -15, 0,
    -- layer=1 filter=140 channel=21
    4, 0, 0, -4, 3, -4, -15, 3, 2,
    -- layer=1 filter=140 channel=22
    -2, -7, -18, -7, -12, -6, -3, 2, -12,
    -- layer=1 filter=140 channel=23
    0, -8, 10, -1, 3, -3, -13, -9, 4,
    -- layer=1 filter=140 channel=24
    -8, -3, 0, -9, -7, -16, -3, -13, 1,
    -- layer=1 filter=140 channel=25
    0, 4, -5, 5, 5, -5, 0, -3, 1,
    -- layer=1 filter=140 channel=26
    -9, -8, -5, -4, -7, 3, -5, -5, -8,
    -- layer=1 filter=140 channel=27
    17, 7, 5, 2, 0, -8, -8, 9, -1,
    -- layer=1 filter=140 channel=28
    -15, -7, -3, -7, -10, -14, -7, -5, -5,
    -- layer=1 filter=140 channel=29
    0, -7, 13, -7, 5, -9, -9, -4, 0,
    -- layer=1 filter=140 channel=30
    -12, -8, -3, -17, 0, -5, -6, 0, 0,
    -- layer=1 filter=140 channel=31
    -11, 3, -14, -18, 6, 3, -5, -6, -11,
    -- layer=1 filter=140 channel=32
    5, -4, -6, -3, 1, 0, 0, 3, -3,
    -- layer=1 filter=140 channel=33
    5, 10, 2, -2, 10, -10, 11, -2, -13,
    -- layer=1 filter=140 channel=34
    7, 0, -10, -3, -7, -11, -7, 1, -5,
    -- layer=1 filter=140 channel=35
    6, -3, 7, 9, 8, 0, 7, -5, -2,
    -- layer=1 filter=140 channel=36
    -8, -1, 9, 0, -3, -11, -7, 8, -6,
    -- layer=1 filter=140 channel=37
    4, -4, 0, 2, 5, -3, 4, -2, -3,
    -- layer=1 filter=140 channel=38
    -17, -4, -3, 0, -15, -17, -14, -5, -3,
    -- layer=1 filter=140 channel=39
    6, 11, 4, -6, 0, -4, -19, 1, 7,
    -- layer=1 filter=140 channel=40
    -3, 2, -5, 2, 6, -16, 10, -5, -16,
    -- layer=1 filter=140 channel=41
    8, -4, -1, 1, 1, -2, 4, -12, 0,
    -- layer=1 filter=140 channel=42
    -7, -1, -1, -8, 15, 6, 2, 6, -11,
    -- layer=1 filter=140 channel=43
    -2, -1, 3, 2, -9, -10, -9, 4, 3,
    -- layer=1 filter=140 channel=44
    -4, -14, -16, 4, -6, -12, 5, -7, -20,
    -- layer=1 filter=140 channel=45
    5, 3, -6, -7, -3, -10, -9, 0, -4,
    -- layer=1 filter=140 channel=46
    -9, 4, 11, 0, 6, 6, -15, -6, -7,
    -- layer=1 filter=140 channel=47
    -2, -11, -3, -1, 2, -11, 0, -13, -11,
    -- layer=1 filter=140 channel=48
    -18, -14, -14, -12, -6, -7, -17, -15, -3,
    -- layer=1 filter=140 channel=49
    -5, -1, -2, -12, 4, -9, -5, -14, 0,
    -- layer=1 filter=140 channel=50
    -5, 0, -8, 0, -3, 4, -6, -7, -9,
    -- layer=1 filter=140 channel=51
    -11, 1, 2, -3, -14, -4, -7, -2, -16,
    -- layer=1 filter=140 channel=52
    8, -8, 0, 4, 2, -9, 10, 4, 0,
    -- layer=1 filter=140 channel=53
    8, 2, -3, -5, -1, 4, -4, -1, 0,
    -- layer=1 filter=140 channel=54
    -8, -5, -5, -11, 0, 4, -10, 4, 0,
    -- layer=1 filter=140 channel=55
    4, 3, 11, 5, 0, -9, -8, -7, 8,
    -- layer=1 filter=140 channel=56
    0, 0, -5, 2, -8, -5, 3, 4, 6,
    -- layer=1 filter=140 channel=57
    -12, 4, -12, -2, -1, -5, -7, 6, -1,
    -- layer=1 filter=140 channel=58
    -4, -7, -9, -5, 5, -5, -9, -3, -4,
    -- layer=1 filter=140 channel=59
    2, -10, 7, -4, -4, -5, -10, -7, 1,
    -- layer=1 filter=140 channel=60
    -3, -10, 9, 0, 2, -1, 8, -8, -3,
    -- layer=1 filter=140 channel=61
    1, -2, 2, -4, 0, -10, 0, 9, 1,
    -- layer=1 filter=140 channel=62
    -11, -12, -11, -8, -7, -1, -12, -10, -15,
    -- layer=1 filter=140 channel=63
    2, -1, 3, 1, 5, -6, 2, -9, 4,
    -- layer=1 filter=140 channel=64
    -2, -12, -15, -1, -8, -9, -6, -3, -14,
    -- layer=1 filter=140 channel=65
    -7, -12, -1, -8, -5, -12, -12, -15, 2,
    -- layer=1 filter=140 channel=66
    -6, 14, -1, -1, 5, -13, -4, 6, 5,
    -- layer=1 filter=140 channel=67
    0, -8, -5, -9, -15, 2, -11, 2, -8,
    -- layer=1 filter=140 channel=68
    -8, -16, -16, -6, -11, 0, 0, -12, -17,
    -- layer=1 filter=140 channel=69
    1, -10, 9, -1, -10, 0, -5, 0, -3,
    -- layer=1 filter=140 channel=70
    -11, -2, -3, -2, 0, -11, 0, -10, -12,
    -- layer=1 filter=140 channel=71
    0, -2, -2, 0, -2, -13, 1, 0, 3,
    -- layer=1 filter=140 channel=72
    1, -1, 10, -9, -4, -1, 6, -12, 7,
    -- layer=1 filter=140 channel=73
    -2, -5, -6, 4, 0, -9, 6, -9, 6,
    -- layer=1 filter=140 channel=74
    -13, -13, -6, -5, 8, 4, -6, -6, -1,
    -- layer=1 filter=140 channel=75
    -9, -5, -11, -4, 0, -15, -12, -13, -7,
    -- layer=1 filter=140 channel=76
    1, 3, -2, -2, 12, 9, 3, 2, 0,
    -- layer=1 filter=140 channel=77
    -4, 0, -17, -15, -2, -4, -15, 0, -1,
    -- layer=1 filter=140 channel=78
    0, -6, 1, 5, -6, 5, -4, 7, 0,
    -- layer=1 filter=140 channel=79
    -8, -5, -14, 2, -7, -7, -14, -6, 3,
    -- layer=1 filter=140 channel=80
    3, -6, 8, -3, 5, -5, 3, -4, -3,
    -- layer=1 filter=140 channel=81
    0, -11, -1, -8, 1, -7, 1, -11, -8,
    -- layer=1 filter=140 channel=82
    -11, -16, -6, 0, 0, -1, -5, 7, 0,
    -- layer=1 filter=140 channel=83
    2, -9, -4, -2, -8, 6, -9, -3, -7,
    -- layer=1 filter=140 channel=84
    -22, -24, 1, -6, -1, 9, 4, -3, 1,
    -- layer=1 filter=140 channel=85
    -5, -5, 1, -8, -7, 0, -2, -7, 5,
    -- layer=1 filter=140 channel=86
    -7, -2, 0, 8, -2, -4, -15, 2, -10,
    -- layer=1 filter=140 channel=87
    -8, -1, 4, -3, 1, -1, 5, -1, -9,
    -- layer=1 filter=140 channel=88
    2, 3, 0, 1, 5, 0, 3, -9, -10,
    -- layer=1 filter=140 channel=89
    3, 0, -14, -2, 0, -3, -7, 3, -12,
    -- layer=1 filter=140 channel=90
    -10, -9, 0, 6, -18, 4, 7, -5, -11,
    -- layer=1 filter=140 channel=91
    -16, -18, -7, -1, -1, 0, 4, 0, -12,
    -- layer=1 filter=140 channel=92
    0, 6, -10, -1, -5, -10, 6, 6, -16,
    -- layer=1 filter=140 channel=93
    3, -9, -8, -2, -5, -7, -3, -3, -11,
    -- layer=1 filter=140 channel=94
    9, 0, -8, -5, -5, -3, -11, 1, -3,
    -- layer=1 filter=140 channel=95
    -7, -14, -15, 3, -3, -10, -13, -13, -2,
    -- layer=1 filter=140 channel=96
    -7, -10, 5, -9, -5, -4, -11, -7, 3,
    -- layer=1 filter=140 channel=97
    -10, 0, -11, -6, -17, 2, -5, -7, -2,
    -- layer=1 filter=140 channel=98
    -2, -7, 1, -1, -11, -11, 4, -4, -3,
    -- layer=1 filter=140 channel=99
    -5, -11, -8, -7, -7, 2, -9, -12, 2,
    -- layer=1 filter=140 channel=100
    -9, 8, 0, -8, -7, 0, 0, -8, 9,
    -- layer=1 filter=140 channel=101
    -12, -17, -15, -8, -18, -16, 3, -3, -2,
    -- layer=1 filter=140 channel=102
    -12, 3, -5, -10, -3, 0, -17, -2, -2,
    -- layer=1 filter=140 channel=103
    -11, -2, -10, -2, -5, -9, 4, 0, 2,
    -- layer=1 filter=140 channel=104
    -5, -5, -11, 3, -7, 2, -2, 7, 5,
    -- layer=1 filter=140 channel=105
    -4, 12, -8, 0, 9, -13, -13, 3, -10,
    -- layer=1 filter=140 channel=106
    -3, -4, -16, -6, -17, 2, 3, -8, -4,
    -- layer=1 filter=140 channel=107
    4, 6, 0, -6, 0, -7, 5, 10, -1,
    -- layer=1 filter=140 channel=108
    -3, -19, -10, -1, 3, -16, 4, -3, -17,
    -- layer=1 filter=140 channel=109
    0, 0, 7, 4, -1, 5, 1, 5, 9,
    -- layer=1 filter=140 channel=110
    7, -11, 0, -7, 3, -6, -3, -6, 6,
    -- layer=1 filter=140 channel=111
    -3, -8, -12, -10, 1, -9, 13, -5, 4,
    -- layer=1 filter=140 channel=112
    -14, 9, 1, -9, 4, 3, 3, -5, 3,
    -- layer=1 filter=140 channel=113
    -4, 4, -7, -14, 12, 2, 0, 8, -9,
    -- layer=1 filter=140 channel=114
    -8, 0, -3, 14, 5, 13, -10, -6, -14,
    -- layer=1 filter=140 channel=115
    4, 0, -10, -13, 5, 1, -18, 15, 5,
    -- layer=1 filter=140 channel=116
    2, -9, 9, 10, 6, 4, -6, 4, 2,
    -- layer=1 filter=140 channel=117
    0, -11, -3, -15, 11, 0, 2, -3, 6,
    -- layer=1 filter=140 channel=118
    -8, -17, -13, 0, 4, -3, 0, -3, 3,
    -- layer=1 filter=140 channel=119
    -3, -6, -3, -8, -2, -16, 2, -2, -9,
    -- layer=1 filter=140 channel=120
    2, -6, -11, -2, 3, 0, 2, 4, 1,
    -- layer=1 filter=140 channel=121
    7, -5, 5, -6, 5, -10, -11, 5, -3,
    -- layer=1 filter=140 channel=122
    -10, -1, 0, -1, -4, 6, -4, -4, 0,
    -- layer=1 filter=140 channel=123
    11, 8, -9, 2, 0, -12, -11, 6, 0,
    -- layer=1 filter=140 channel=124
    -9, 0, -1, 2, 1, 1, -7, 0, 6,
    -- layer=1 filter=140 channel=125
    0, -6, -14, -10, -3, -10, -9, -6, 3,
    -- layer=1 filter=140 channel=126
    -1, -3, 0, -3, -8, -3, 2, 0, -4,
    -- layer=1 filter=140 channel=127
    -16, -22, -10, 0, -4, -7, -5, -13, -9,
    -- layer=1 filter=141 channel=0
    -50, -65, -37, -44, -30, -33, -23, -21, -34,
    -- layer=1 filter=141 channel=1
    11, 11, -26, -23, -21, -3, -21, -1, -21,
    -- layer=1 filter=141 channel=2
    53, 79, 64, 64, 63, 62, 63, 58, 20,
    -- layer=1 filter=141 channel=3
    -6, 5, 0, -14, 0, 11, 2, 8, 0,
    -- layer=1 filter=141 channel=4
    9, -14, 12, -12, -5, -8, -20, -22, -16,
    -- layer=1 filter=141 channel=5
    50, 42, 10, -25, -5, -6, -10, -7, -12,
    -- layer=1 filter=141 channel=6
    -29, -15, 6, -26, -4, -8, -35, -20, -1,
    -- layer=1 filter=141 channel=7
    14, 17, 9, -21, 29, 12, -14, 18, 24,
    -- layer=1 filter=141 channel=8
    49, 29, 11, -19, -2, -6, -1, -10, -10,
    -- layer=1 filter=141 channel=9
    40, -10, -15, -25, -4, 11, 12, -8, 4,
    -- layer=1 filter=141 channel=10
    20, 35, 13, -9, 35, 35, -13, 45, 41,
    -- layer=1 filter=141 channel=11
    9, 5, -8, 11, 8, -29, 1, -9, -16,
    -- layer=1 filter=141 channel=12
    13, -32, -1, -60, 4, -1, 17, 29, -16,
    -- layer=1 filter=141 channel=13
    1, 5, 9, 3, 1, -1, -8, 4, 12,
    -- layer=1 filter=141 channel=14
    0, 35, 10, -59, 23, -16, -20, 41, 5,
    -- layer=1 filter=141 channel=15
    49, 67, 25, 26, 22, 24, 6, -1, 27,
    -- layer=1 filter=141 channel=16
    54, 33, 24, -8, -4, -3, -3, -3, 1,
    -- layer=1 filter=141 channel=17
    -70, -60, -58, -35, -26, -61, -27, -48, -33,
    -- layer=1 filter=141 channel=18
    -3, 3, -12, -100, -82, -68, -38, -43, -16,
    -- layer=1 filter=141 channel=19
    1, -5, -12, -34, -55, -30, -29, -46, -24,
    -- layer=1 filter=141 channel=20
    -14, -8, 13, -20, -18, -9, -29, -21, 6,
    -- layer=1 filter=141 channel=21
    -15, -22, 1, 3, -7, 17, -13, 19, 20,
    -- layer=1 filter=141 channel=22
    0, -8, 3, 13, 13, 4, -6, -11, 6,
    -- layer=1 filter=141 channel=23
    28, 0, -8, 43, 38, 67, 32, 7, 88,
    -- layer=1 filter=141 channel=24
    7, 0, 7, 19, 24, 4, 22, 19, 20,
    -- layer=1 filter=141 channel=25
    52, 5, 6, -13, 28, 26, -16, 5, 38,
    -- layer=1 filter=141 channel=26
    -8, 39, -8, 6, 32, -8, 5, 11, 10,
    -- layer=1 filter=141 channel=27
    22, 0, 18, 26, 24, 8, 26, 26, 29,
    -- layer=1 filter=141 channel=28
    -4, 12, -14, -46, 9, -3, -28, 22, 6,
    -- layer=1 filter=141 channel=29
    16, 11, 35, 33, 19, 26, 5, 29, 10,
    -- layer=1 filter=141 channel=30
    -43, -25, -45, -116, -106, -52, -44, -50, -52,
    -- layer=1 filter=141 channel=31
    32, 51, 31, 16, 22, 32, 17, 28, 3,
    -- layer=1 filter=141 channel=32
    16, 29, -42, 11, 34, 23, -4, 12, 28,
    -- layer=1 filter=141 channel=33
    -13, -15, -18, -15, 0, 17, 4, 9, 24,
    -- layer=1 filter=141 channel=34
    3, -4, -9, -9, -11, 11, -6, -12, 21,
    -- layer=1 filter=141 channel=35
    16, 20, 7, -21, 4, 0, -3, -16, -10,
    -- layer=1 filter=141 channel=36
    -12, -7, -17, -6, -20, -33, 9, 6, -32,
    -- layer=1 filter=141 channel=37
    46, 34, 23, -15, 10, 8, 6, -5, 4,
    -- layer=1 filter=141 channel=38
    -24, -9, 10, -21, -4, 0, -7, -12, 1,
    -- layer=1 filter=141 channel=39
    -41, -56, -38, -43, -35, -50, -13, -14, -42,
    -- layer=1 filter=141 channel=40
    19, 35, 38, -27, 0, 15, -13, 3, -4,
    -- layer=1 filter=141 channel=41
    24, 22, -35, -23, 0, -2, -11, 13, 65,
    -- layer=1 filter=141 channel=42
    54, 75, 90, 40, 64, 61, 47, 52, 36,
    -- layer=1 filter=141 channel=43
    41, 12, 7, 5, -1, 30, -1, 8, 0,
    -- layer=1 filter=141 channel=44
    -2, 19, -17, 7, 27, -1, 19, 24, 2,
    -- layer=1 filter=141 channel=45
    2, 7, 6, 13, 7, -10, 13, 0, -4,
    -- layer=1 filter=141 channel=46
    53, 44, 43, -7, -5, 1, -17, -22, -4,
    -- layer=1 filter=141 channel=47
    36, 27, -1, 17, 49, 75, -7, 26, 63,
    -- layer=1 filter=141 channel=48
    -52, -44, -33, -36, -33, 9, -22, -18, 28,
    -- layer=1 filter=141 channel=49
    13, 13, 25, 5, 23, 37, 7, 24, 26,
    -- layer=1 filter=141 channel=50
    -32, 0, -23, -22, -25, -14, 7, -21, -7,
    -- layer=1 filter=141 channel=51
    -29, -20, 3, -37, -13, 15, -23, -14, 18,
    -- layer=1 filter=141 channel=52
    2, -7, -18, -19, -10, -27, -19, -1, 24,
    -- layer=1 filter=141 channel=53
    -8, -40, 14, -10, -6, -12, -26, -8, -11,
    -- layer=1 filter=141 channel=54
    57, 35, 31, 11, 42, 37, -3, 19, 41,
    -- layer=1 filter=141 channel=55
    33, 42, 30, 29, 29, 33, 21, 32, 8,
    -- layer=1 filter=141 channel=56
    -12, -4, -10, 0, 1, -10, -6, 2, -12,
    -- layer=1 filter=141 channel=57
    27, 31, 28, -18, 29, 29, -17, 25, 32,
    -- layer=1 filter=141 channel=58
    30, 23, 14, 40, 51, 74, 8, 41, 74,
    -- layer=1 filter=141 channel=59
    -15, -6, 0, -18, 26, 2, -10, 2, -29,
    -- layer=1 filter=141 channel=60
    -44, -3, -28, -20, 18, -11, -18, 16, -17,
    -- layer=1 filter=141 channel=61
    -6, -17, 5, -18, -2, -19, -7, 0, -6,
    -- layer=1 filter=141 channel=62
    22, 15, 16, -31, 5, -7, -2, 0, 11,
    -- layer=1 filter=141 channel=63
    -42, -44, -20, -30, -43, -28, 3, -10, -6,
    -- layer=1 filter=141 channel=64
    -15, -32, -9, -16, -11, -13, -20, 0, 2,
    -- layer=1 filter=141 channel=65
    -40, -40, -17, -26, -1, -6, -11, -7, 8,
    -- layer=1 filter=141 channel=66
    -27, -55, -57, -20, -25, -21, -2, -7, -11,
    -- layer=1 filter=141 channel=67
    7, -31, -18, 20, -10, -10, 8, -19, 11,
    -- layer=1 filter=141 channel=68
    0, 16, 1, 20, 42, 11, 12, 21, -3,
    -- layer=1 filter=141 channel=69
    62, 69, 38, 2, 5, -7, 18, 8, 12,
    -- layer=1 filter=141 channel=70
    19, -7, 21, -10, 9, 15, -9, 14, 4,
    -- layer=1 filter=141 channel=71
    -4, -17, -19, 8, 5, 16, 23, 15, 40,
    -- layer=1 filter=141 channel=72
    -17, -14, -31, -100, -58, -38, -30, -89, -40,
    -- layer=1 filter=141 channel=73
    11, 3, 1, 4, -10, 12, 6, 12, 21,
    -- layer=1 filter=141 channel=74
    -24, -10, -36, -71, 18, -26, -25, 15, 41,
    -- layer=1 filter=141 channel=75
    0, 16, 19, -90, 10, -53, 11, -3, -24,
    -- layer=1 filter=141 channel=76
    -49, -62, -71, -44, -59, -56, -56, -29, 7,
    -- layer=1 filter=141 channel=77
    -39, -49, -24, -15, 13, -2, 13, 16, 17,
    -- layer=1 filter=141 channel=78
    -28, -40, -27, -44, -4, -4, -20, 4, 3,
    -- layer=1 filter=141 channel=79
    32, 13, 5, -16, 7, 13, 6, 11, 21,
    -- layer=1 filter=141 channel=80
    -10, 5, -19, 13, 0, 4, -9, -7, -24,
    -- layer=1 filter=141 channel=81
    4, -26, -16, 12, 23, 28, 32, 8, 28,
    -- layer=1 filter=141 channel=82
    -28, -35, -17, -18, -8, 1, 0, 6, 23,
    -- layer=1 filter=141 channel=83
    -38, 0, -27, -20, -26, -13, -35, -28, -55,
    -- layer=1 filter=141 channel=84
    -7, -17, -46, -48, -48, -79, -34, -18, -11,
    -- layer=1 filter=141 channel=85
    2, 19, -10, 13, 42, 50, -1, 7, 84,
    -- layer=1 filter=141 channel=86
    28, -11, -7, -16, -10, -22, -7, 0, -10,
    -- layer=1 filter=141 channel=87
    58, 25, 0, -26, -16, 23, 21, 11, -11,
    -- layer=1 filter=141 channel=88
    13, -11, 4, 24, 9, 13, 15, 2, 23,
    -- layer=1 filter=141 channel=89
    -31, -29, -39, -17, -22, -3, -11, -16, 14,
    -- layer=1 filter=141 channel=90
    -9, 10, -4, -4, 27, -23, 19, 11, 1,
    -- layer=1 filter=141 channel=91
    -21, -12, 5, -27, -18, 5, -11, -25, 7,
    -- layer=1 filter=141 channel=92
    44, 48, -15, 28, 25, 28, 4, -19, 33,
    -- layer=1 filter=141 channel=93
    -32, -38, -26, -15, -5, -7, -5, -10, 0,
    -- layer=1 filter=141 channel=94
    -49, -85, -61, -59, -53, -44, -35, -22, -27,
    -- layer=1 filter=141 channel=95
    -41, -53, -37, -122, -89, -83, -37, -41, -5,
    -- layer=1 filter=141 channel=96
    -25, -29, -25, -11, -22, -22, 3, -21, -20,
    -- layer=1 filter=141 channel=97
    -53, -68, -61, -34, -17, -30, -8, -9, -20,
    -- layer=1 filter=141 channel=98
    -3, 9, -14, -6, 14, 9, -11, -4, 3,
    -- layer=1 filter=141 channel=99
    -13, 38, 7, -7, 67, 24, 1, 82, 16,
    -- layer=1 filter=141 channel=100
    -23, -18, -35, -33, -37, -59, -14, -15, 0,
    -- layer=1 filter=141 channel=101
    -25, -34, -13, -16, -21, -7, -26, -10, 7,
    -- layer=1 filter=141 channel=102
    -75, -83, -87, -75, -62, -91, -55, -51, -51,
    -- layer=1 filter=141 channel=103
    -17, -16, -16, 5, -36, -28, -20, -20, -20,
    -- layer=1 filter=141 channel=104
    12, 11, -13, 15, 3, -10, -17, -1, 46,
    -- layer=1 filter=141 channel=105
    -56, -70, -49, -36, -27, -11, -21, -10, -9,
    -- layer=1 filter=141 channel=106
    0, 13, -18, 10, 3, 15, -13, -21, 8,
    -- layer=1 filter=141 channel=107
    7, -5, -9, -2, -10, -5, 4, 3, -3,
    -- layer=1 filter=141 channel=108
    17, 44, -14, 15, 25, 37, 22, 21, 23,
    -- layer=1 filter=141 channel=109
    -9, -4, 7, 1, -5, 3, -10, 3, -2,
    -- layer=1 filter=141 channel=110
    -33, -23, -9, -28, -15, 1, -4, -10, 0,
    -- layer=1 filter=141 channel=111
    -50, -54, -30, -154, -110, -66, -72, -45, -42,
    -- layer=1 filter=141 channel=112
    -48, -87, -73, -108, -62, -31, -60, -28, 4,
    -- layer=1 filter=141 channel=113
    26, 48, 50, 0, 34, 34, 4, 18, 50,
    -- layer=1 filter=141 channel=114
    75, 59, 47, -16, -5, 7, 17, 10, -10,
    -- layer=1 filter=141 channel=115
    2, -10, -14, -20, -7, 1, -9, -6, 18,
    -- layer=1 filter=141 channel=116
    -6, 0, 9, 8, -1, 10, 2, 5, -5,
    -- layer=1 filter=141 channel=117
    -57, -79, 14, -86, -76, -7, -56, -70, -11,
    -- layer=1 filter=141 channel=118
    -23, -9, -39, -78, -58, -49, -13, -13, -13,
    -- layer=1 filter=141 channel=119
    5, 12, -40, 13, 23, 9, 7, 32, 37,
    -- layer=1 filter=141 channel=120
    -9, -31, -2, -8, -4, 3, -9, 0, 31,
    -- layer=1 filter=141 channel=121
    -12, 1, 6, -2, -4, -4, 11, 12, -2,
    -- layer=1 filter=141 channel=122
    0, -7, 1, 0, 10, -7, -7, -10, -7,
    -- layer=1 filter=141 channel=123
    2, 18, 23, 16, 9, 5, 28, 1, 12,
    -- layer=1 filter=141 channel=124
    -2, 0, 27, 29, 18, 21, 1, -6, -12,
    -- layer=1 filter=141 channel=125
    18, 20, 28, 5, 22, 40, -13, 21, 32,
    -- layer=1 filter=141 channel=126
    -39, -13, -34, -23, 7, -9, -48, -39, -39,
    -- layer=1 filter=141 channel=127
    -23, 0, -30, -125, -68, -82, -29, -39, -34,
    -- layer=1 filter=142 channel=0
    3, 0, -33, 8, -28, 5, 0, 5, 26,
    -- layer=1 filter=142 channel=1
    -55, -27, -33, -73, -60, 64, -10, 36, 44,
    -- layer=1 filter=142 channel=2
    -29, 22, 0, 0, 16, -15, 32, -8, -26,
    -- layer=1 filter=142 channel=3
    9, -10, -4, -6, -3, 2, -7, 2, 10,
    -- layer=1 filter=142 channel=4
    -11, -8, -18, -9, 12, -6, -14, -6, -18,
    -- layer=1 filter=142 channel=5
    -38, -64, -9, -86, -33, 77, -11, 31, -12,
    -- layer=1 filter=142 channel=6
    23, -10, 4, 9, 41, -20, -8, -63, 11,
    -- layer=1 filter=142 channel=7
    -29, -2, -14, -67, -17, 63, 34, 83, 12,
    -- layer=1 filter=142 channel=8
    -24, -88, -29, -75, -32, 79, -9, 59, 12,
    -- layer=1 filter=142 channel=9
    -40, 41, 37, 86, 44, 37, 44, -19, 10,
    -- layer=1 filter=142 channel=10
    -24, -22, 16, -51, -1, 87, 41, 85, -5,
    -- layer=1 filter=142 channel=11
    11, 5, 17, 21, -12, 1, -21, -13, 50,
    -- layer=1 filter=142 channel=12
    -15, 18, -48, -31, -5, -28, -58, -19, -39,
    -- layer=1 filter=142 channel=13
    -15, -15, 18, 18, 36, -36, 11, -25, -5,
    -- layer=1 filter=142 channel=14
    -5, 20, -36, -37, -35, 14, -79, -32, -13,
    -- layer=1 filter=142 channel=15
    -18, -4, -111, -69, -45, -28, -58, -64, -109,
    -- layer=1 filter=142 channel=16
    -50, -77, 1, -61, -9, 102, 1, 67, -11,
    -- layer=1 filter=142 channel=17
    -23, -14, 14, -19, -10, 27, -9, 24, 15,
    -- layer=1 filter=142 channel=18
    -52, 16, -14, 11, -17, -24, -2, -48, 34,
    -- layer=1 filter=142 channel=19
    -77, -38, 74, 9, 104, 125, 80, 116, -57,
    -- layer=1 filter=142 channel=20
    -26, -19, 11, -25, -6, 51, -26, 24, 7,
    -- layer=1 filter=142 channel=21
    2, -6, -21, 3, -13, 0, -15, 6, 37,
    -- layer=1 filter=142 channel=22
    -11, -26, -3, -39, -81, 41, -46, 21, 62,
    -- layer=1 filter=142 channel=23
    -69, -41, -21, -120, -29, -51, -45, 4, -142,
    -- layer=1 filter=142 channel=24
    8, -8, 9, -1, 19, -11, 4, -8, -88,
    -- layer=1 filter=142 channel=25
    -34, -35, 27, -41, 35, 108, 61, 130, 13,
    -- layer=1 filter=142 channel=26
    -33, 19, 6, 20, -7, -102, -25, -77, -18,
    -- layer=1 filter=142 channel=27
    22, 27, 41, 1, -14, -12, -4, -28, 19,
    -- layer=1 filter=142 channel=28
    -7, -4, -15, -44, -24, 80, 29, 58, 32,
    -- layer=1 filter=142 channel=29
    -3, 4, -3, -18, -50, -12, 7, 9, 11,
    -- layer=1 filter=142 channel=30
    -65, 2, -16, 6, 4, 5, 47, -63, 8,
    -- layer=1 filter=142 channel=31
    -34, -27, -42, -47, -18, -15, -43, -97, -6,
    -- layer=1 filter=142 channel=32
    -32, 22, 16, 27, 1, -161, -1, -111, -14,
    -- layer=1 filter=142 channel=33
    19, -4, 31, 13, -31, 17, 0, 3, 36,
    -- layer=1 filter=142 channel=34
    59, 50, 15, 35, 27, -17, 17, -23, 13,
    -- layer=1 filter=142 channel=35
    -6, -5, -20, -24, -23, -23, -31, -23, -10,
    -- layer=1 filter=142 channel=36
    23, 17, 21, 17, -2, -9, -7, -3, 40,
    -- layer=1 filter=142 channel=37
    -29, -50, 49, -77, 25, 100, 23, 67, -39,
    -- layer=1 filter=142 channel=38
    -8, -9, 6, 13, 9, 11, 12, -11, 4,
    -- layer=1 filter=142 channel=39
    33, 4, 26, 4, -5, 17, -23, 18, 2,
    -- layer=1 filter=142 channel=40
    -50, -6, -15, -12, 0, -4, -58, -91, -16,
    -- layer=1 filter=142 channel=41
    -47, 60, 68, 81, 62, -7, 59, 3, -43,
    -- layer=1 filter=142 channel=42
    -1, 25, 39, 19, 44, -10, 60, 33, -46,
    -- layer=1 filter=142 channel=43
    -49, -50, 5, -56, -13, 104, 8, 83, 12,
    -- layer=1 filter=142 channel=44
    -22, -8, -13, 1, -39, -160, -55, -115, 24,
    -- layer=1 filter=142 channel=45
    -13, -17, -34, -32, -48, -28, -39, -54, -25,
    -- layer=1 filter=142 channel=46
    -84, -117, -9, -42, 46, 40, 28, 48, -60,
    -- layer=1 filter=142 channel=47
    -31, 16, 12, 9, 58, -87, 32, -43, -177,
    -- layer=1 filter=142 channel=48
    -5, 15, -3, 17, -1, -28, 1, 0, -22,
    -- layer=1 filter=142 channel=49
    5, 7, 22, 46, 44, -28, 44, -1, -25,
    -- layer=1 filter=142 channel=50
    -26, -37, -30, 6, -21, -19, -49, -25, 18,
    -- layer=1 filter=142 channel=51
    2, -1, -13, -1, -7, 35, 35, 36, -10,
    -- layer=1 filter=142 channel=52
    -14, 2, 9, 2, 16, -32, 14, 20, -1,
    -- layer=1 filter=142 channel=53
    5, 3, 8, 3, 1, -5, 12, 17, 3,
    -- layer=1 filter=142 channel=54
    -21, -46, 40, -38, 47, 130, 59, 146, -26,
    -- layer=1 filter=142 channel=55
    35, 17, 34, -7, 13, -15, -10, -4, 15,
    -- layer=1 filter=142 channel=56
    -6, -9, -3, 7, 3, -8, 4, -9, -9,
    -- layer=1 filter=142 channel=57
    -12, -27, 11, -43, -4, 75, 31, 65, -16,
    -- layer=1 filter=142 channel=58
    -81, -22, 25, -60, 54, 7, 49, 79, -136,
    -- layer=1 filter=142 channel=59
    -4, 3, -1, -24, 0, 16, 9, 20, 25,
    -- layer=1 filter=142 channel=60
    22, -21, 0, 16, 5, 14, -11, 12, -12,
    -- layer=1 filter=142 channel=61
    -3, -7, 4, -8, 3, 10, -9, 0, 9,
    -- layer=1 filter=142 channel=62
    -23, -55, 28, -75, 17, 112, 4, 86, -28,
    -- layer=1 filter=142 channel=63
    0, 15, 2, 17, -9, -31, -9, -14, 46,
    -- layer=1 filter=142 channel=64
    22, 7, -14, 11, -31, 10, -16, 14, 44,
    -- layer=1 filter=142 channel=65
    19, -6, -22, -9, -20, 2, -26, -21, 4,
    -- layer=1 filter=142 channel=66
    13, 10, -17, -14, -10, 1, -22, 27, 45,
    -- layer=1 filter=142 channel=67
    45, 58, 17, 17, 18, -27, 46, 11, -10,
    -- layer=1 filter=142 channel=68
    -23, 8, 5, 7, -26, -149, -50, -113, 50,
    -- layer=1 filter=142 channel=69
    -43, -42, -56, -67, -25, 20, -25, -12, -80,
    -- layer=1 filter=142 channel=70
    33, -1, 1, 36, 42, -32, 58, -87, -43,
    -- layer=1 filter=142 channel=71
    8, -21, -18, -15, -13, 10, -3, 29, -9,
    -- layer=1 filter=142 channel=72
    -66, 0, 26, 24, 39, 57, 83, -11, 12,
    -- layer=1 filter=142 channel=73
    6, 3, -8, -3, -4, 18, -2, -3, 10,
    -- layer=1 filter=142 channel=74
    -12, -32, -13, 10, 18, -66, -57, -39, 92,
    -- layer=1 filter=142 channel=75
    -42, 0, -54, -32, -25, -49, -52, -54, -25,
    -- layer=1 filter=142 channel=76
    -15, 26, 22, 48, 38, -54, 8, -6, 23,
    -- layer=1 filter=142 channel=77
    -4, 0, -20, -25, -33, 3, -7, 2, 2,
    -- layer=1 filter=142 channel=78
    -1, 0, -20, -17, -2, 19, 18, 17, 15,
    -- layer=1 filter=142 channel=79
    -26, -60, 23, -67, 22, 82, 0, 75, -32,
    -- layer=1 filter=142 channel=80
    10, 1, 46, -29, 10, 27, 15, -2, 23,
    -- layer=1 filter=142 channel=81
    4, -23, -3, -20, 12, 2, -8, 38, -28,
    -- layer=1 filter=142 channel=82
    13, 6, -7, 21, -12, -18, 2, 12, -13,
    -- layer=1 filter=142 channel=83
    -31, -51, -43, -60, -103, -72, -56, -48, -32,
    -- layer=1 filter=142 channel=84
    -33, 21, 46, 75, 42, -15, 62, -34, 89,
    -- layer=1 filter=142 channel=85
    -5, -6, 56, -25, 47, 13, 72, 68, -110,
    -- layer=1 filter=142 channel=86
    17, -10, -5, -29, -14, 20, -37, 2, 60,
    -- layer=1 filter=142 channel=87
    -47, -3, 62, 45, 80, 91, 83, 49, -26,
    -- layer=1 filter=142 channel=88
    -3, -6, 0, 13, 13, -22, 10, 4, -4,
    -- layer=1 filter=142 channel=89
    7, 17, -14, 40, 7, -53, -9, -37, 27,
    -- layer=1 filter=142 channel=90
    -43, -42, -69, -34, -90, -150, -68, -126, -31,
    -- layer=1 filter=142 channel=91
    -5, 4, -7, -17, 3, 2, 19, -7, -2,
    -- layer=1 filter=142 channel=92
    -9, -13, -76, -23, -44, -92, -2, -71, -65,
    -- layer=1 filter=142 channel=93
    9, 1, -18, -16, -10, -10, -4, 4, 4,
    -- layer=1 filter=142 channel=94
    13, 12, -17, 0, -29, 10, -10, -5, 48,
    -- layer=1 filter=142 channel=95
    1, 17, 6, 35, 21, -67, 6, -44, 63,
    -- layer=1 filter=142 channel=96
    5, 21, 10, -8, 9, -25, -12, -21, 0,
    -- layer=1 filter=142 channel=97
    3, 0, -17, -18, -37, 21, -23, 19, 28,
    -- layer=1 filter=142 channel=98
    -57, -52, 0, -68, -14, 96, -10, 87, 4,
    -- layer=1 filter=142 channel=99
    -42, -76, -69, -112, -129, 0, -101, -52, -6,
    -- layer=1 filter=142 channel=100
    5, 8, 7, 4, -17, -18, 3, -17, 45,
    -- layer=1 filter=142 channel=101
    -1, 5, 3, 17, 6, -29, 0, -20, 29,
    -- layer=1 filter=142 channel=102
    14, 6, -18, -5, -27, 10, -18, -42, 11,
    -- layer=1 filter=142 channel=103
    16, -10, 13, 14, -9, 7, -2, -16, 12,
    -- layer=1 filter=142 channel=104
    -24, -15, -23, -41, -29, -63, -21, -5, -115,
    -- layer=1 filter=142 channel=105
    20, 6, -9, -1, -32, 17, -20, 17, 19,
    -- layer=1 filter=142 channel=106
    -11, 16, 17, 23, 13, -83, -18, -88, 20,
    -- layer=1 filter=142 channel=107
    4, -2, 17, 14, 7, 20, 6, 18, 20,
    -- layer=1 filter=142 channel=108
    -34, 3, -12, -1, -21, -173, -37, -117, -65,
    -- layer=1 filter=142 channel=109
    -10, 5, -8, 7, 9, 8, -1, 6, 2,
    -- layer=1 filter=142 channel=110
    -14, 3, -10, -8, -26, 2, -7, -4, 3,
    -- layer=1 filter=142 channel=111
    -50, 26, 1, 42, 3, -34, -5, -82, -3,
    -- layer=1 filter=142 channel=112
    -4, 14, 1, 26, 5, -42, 30, 3, 66,
    -- layer=1 filter=142 channel=113
    10, -17, 41, -6, 13, 1, 5, 39, -62,
    -- layer=1 filter=142 channel=114
    -3, -5, -37, -46, -33, 39, -50, -38, -20,
    -- layer=1 filter=142 channel=115
    5, -20, 5, -31, -24, 49, 0, 37, 6,
    -- layer=1 filter=142 channel=116
    -8, -8, 0, 1, -5, 0, -1, -10, 7,
    -- layer=1 filter=142 channel=117
    -40, 3, -6, -46, -55, -77, -19, -58, -15,
    -- layer=1 filter=142 channel=118
    -51, 6, 2, 28, 11, -32, 10, -72, 26,
    -- layer=1 filter=142 channel=119
    -43, 6, 34, 23, -1, -133, -10, -64, -45,
    -- layer=1 filter=142 channel=120
    -24, -13, -13, -24, 8, 44, 28, 73, -32,
    -- layer=1 filter=142 channel=121
    -25, -21, -39, -29, -69, -37, 0, -63, -23,
    -- layer=1 filter=142 channel=122
    -9, 6, 3, 8, -1, 0, 2, 2, 0,
    -- layer=1 filter=142 channel=123
    13, -6, -3, -3, -16, -54, 1, -8, -27,
    -- layer=1 filter=142 channel=124
    -7, -7, 4, -16, -22, -11, 23, 11, -14,
    -- layer=1 filter=142 channel=125
    42, -8, 6, 28, 28, -11, 57, -37, -28,
    -- layer=1 filter=142 channel=126
    -61, -37, -59, -90, -101, 26, -17, 65, 0,
    -- layer=1 filter=142 channel=127
    -39, 4, -20, 28, 9, -27, -2, -36, 45,
    -- layer=1 filter=143 channel=0
    -13, -8, 1, -49, -40, -36, -35, -29, -10,
    -- layer=1 filter=143 channel=1
    -13, -27, -64, -93, -70, -57, -22, -43, -40,
    -- layer=1 filter=143 channel=2
    1, 22, 15, 59, 56, 56, 65, 69, 65,
    -- layer=1 filter=143 channel=3
    6, 2, 8, 11, -4, 8, -4, -2, 0,
    -- layer=1 filter=143 channel=4
    18, 9, 16, 0, 14, 3, 4, 3, -9,
    -- layer=1 filter=143 channel=5
    -66, -46, -102, -103, -79, -70, -29, -36, -12,
    -- layer=1 filter=143 channel=6
    22, 28, 23, 20, 3, -11, -53, -29, -31,
    -- layer=1 filter=143 channel=7
    -11, -22, -5, -132, -71, -43, -64, -34, -22,
    -- layer=1 filter=143 channel=8
    -28, -53, -119, -95, -81, -76, -24, -45, -11,
    -- layer=1 filter=143 channel=9
    49, 26, 50, 13, 11, -5, 18, 20, 14,
    -- layer=1 filter=143 channel=10
    -11, -43, -23, -96, -50, -44, -43, -22, 5,
    -- layer=1 filter=143 channel=11
    26, 8, 8, 23, 14, 26, 25, 22, 37,
    -- layer=1 filter=143 channel=12
    32, 24, 16, 41, 4, 36, -43, -16, -21,
    -- layer=1 filter=143 channel=13
    9, -8, -20, -5, 0, -15, 0, 3, -9,
    -- layer=1 filter=143 channel=14
    10, 24, 18, -37, -8, -9, -60, 0, -42,
    -- layer=1 filter=143 channel=15
    -51, -48, -59, -52, -41, -41, 16, -35, -25,
    -- layer=1 filter=143 channel=16
    -63, -92, -97, -134, -84, -72, -10, -54, -18,
    -- layer=1 filter=143 channel=17
    -28, -13, -49, -55, -76, -46, -63, -66, -40,
    -- layer=1 filter=143 channel=18
    38, 32, 57, 19, 5, 2, -7, 0, -16,
    -- layer=1 filter=143 channel=19
    42, 16, 47, 14, 25, -10, -39, -43, 6,
    -- layer=1 filter=143 channel=20
    -9, -30, -34, -32, -13, -32, -13, -17, -23,
    -- layer=1 filter=143 channel=21
    0, -8, 5, 5, 23, 13, 8, 15, 0,
    -- layer=1 filter=143 channel=22
    -53, -41, -28, -20, -17, -20, 12, -24, -8,
    -- layer=1 filter=143 channel=23
    -1, -30, -18, -34, -42, -50, 2, -7, -18,
    -- layer=1 filter=143 channel=24
    16, 1, -1, 18, 16, 28, 22, 23, 14,
    -- layer=1 filter=143 channel=25
    -9, -51, -27, -116, -47, -59, -13, -24, 1,
    -- layer=1 filter=143 channel=26
    20, -10, 0, 4, -3, -32, 2, -18, -34,
    -- layer=1 filter=143 channel=27
    -26, -12, -12, 35, 20, 22, 37, 31, 47,
    -- layer=1 filter=143 channel=28
    -34, -77, -22, -90, -71, -41, -28, -22, -4,
    -- layer=1 filter=143 channel=29
    -29, -49, -37, -40, -46, -28, -25, -43, -22,
    -- layer=1 filter=143 channel=30
    51, 49, 43, 23, 19, 8, -54, -23, -15,
    -- layer=1 filter=143 channel=31
    48, 57, 54, 43, 33, 41, 10, 40, 48,
    -- layer=1 filter=143 channel=32
    53, 25, 21, 20, -15, -56, 16, 1, -47,
    -- layer=1 filter=143 channel=33
    1, -4, -23, 41, 32, 26, -16, -7, -19,
    -- layer=1 filter=143 channel=34
    18, 28, 23, -13, 16, 25, -1, 0, -13,
    -- layer=1 filter=143 channel=35
    14, 3, 3, -3, -8, 0, 34, 0, 0,
    -- layer=1 filter=143 channel=36
    6, 2, -4, 18, 5, 1, 10, 0, 15,
    -- layer=1 filter=143 channel=37
    -72, -76, -61, -115, -71, -42, -11, -32, 7,
    -- layer=1 filter=143 channel=38
    11, -8, -5, 16, 15, 0, 0, 16, 10,
    -- layer=1 filter=143 channel=39
    -42, -35, -48, -30, -13, -35, -13, -8, 10,
    -- layer=1 filter=143 channel=40
    44, 36, 34, 15, -4, 6, -38, 4, -6,
    -- layer=1 filter=143 channel=41
    44, 46, 25, 42, -12, -1, 18, 17, -30,
    -- layer=1 filter=143 channel=42
    7, 13, 25, 55, 48, 51, 61, 81, 65,
    -- layer=1 filter=143 channel=43
    -42, -35, -52, -122, -67, -51, -24, -59, -13,
    -- layer=1 filter=143 channel=44
    12, -12, -25, -5, -38, -69, -1, -30, -65,
    -- layer=1 filter=143 channel=45
    -9, -17, -31, -27, -1, -13, -6, -27, -34,
    -- layer=1 filter=143 channel=46
    11, -1, 33, -13, 6, 0, -21, 16, 20,
    -- layer=1 filter=143 channel=47
    35, 18, 16, 28, 17, 20, 46, 28, 20,
    -- layer=1 filter=143 channel=48
    -5, -10, -12, -5, -3, -8, -18, -27, -28,
    -- layer=1 filter=143 channel=49
    25, 29, 29, 37, 10, 25, 30, 55, 37,
    -- layer=1 filter=143 channel=50
    55, 21, 4, -1, 7, -12, 16, 9, 3,
    -- layer=1 filter=143 channel=51
    29, -1, 4, -12, 7, -3, 0, 13, 2,
    -- layer=1 filter=143 channel=52
    -3, -6, 8, -4, -28, -30, -15, -24, -8,
    -- layer=1 filter=143 channel=53
    1, 0, -6, 6, -4, 0, 1, -5, -13,
    -- layer=1 filter=143 channel=54
    -25, -45, -12, -56, -11, -30, 4, -5, 43,
    -- layer=1 filter=143 channel=55
    18, -5, 2, 32, 23, 27, 33, 42, 36,
    -- layer=1 filter=143 channel=56
    -5, -9, 7, -1, -6, -9, -9, 8, -10,
    -- layer=1 filter=143 channel=57
    -21, -35, -5, -35, -13, -31, -10, -11, 9,
    -- layer=1 filter=143 channel=58
    -38, -43, -21, -37, -26, -37, -31, -21, 0,
    -- layer=1 filter=143 channel=59
    -7, -16, -16, -2, -4, -11, -1, -2, -28,
    -- layer=1 filter=143 channel=60
    -21, -37, 0, -28, 24, -14, -12, 14, 18,
    -- layer=1 filter=143 channel=61
    4, -8, 2, 5, 3, -8, 7, 12, 1,
    -- layer=1 filter=143 channel=62
    -53, -96, -112, -155, -99, -80, -29, -68, -29,
    -- layer=1 filter=143 channel=63
    20, 12, 23, -1, -4, -5, 12, 14, 4,
    -- layer=1 filter=143 channel=64
    10, -14, -18, -29, -16, -7, -29, -15, -9,
    -- layer=1 filter=143 channel=65
    -17, -43, -41, -23, -10, -24, -16, -29, -34,
    -- layer=1 filter=143 channel=66
    -5, -8, 1, -24, -19, -18, -19, -12, -11,
    -- layer=1 filter=143 channel=67
    29, 18, 10, 7, -12, -30, -6, -25, -30,
    -- layer=1 filter=143 channel=68
    15, -9, -3, -6, -58, -78, -32, -28, -71,
    -- layer=1 filter=143 channel=69
    -37, -43, -70, -46, -49, -28, 16, -26, -32,
    -- layer=1 filter=143 channel=70
    51, 48, 42, 5, -16, -16, -20, -11, -4,
    -- layer=1 filter=143 channel=71
    -12, -3, -12, 6, 20, 19, 13, 16, 4,
    -- layer=1 filter=143 channel=72
    59, 38, 42, 26, 27, -6, -24, 4, -20,
    -- layer=1 filter=143 channel=73
    -9, -1, -2, 0, -8, 2, -21, 0, -5,
    -- layer=1 filter=143 channel=74
    34, 28, 55, 1, -39, -49, -80, 3, -45,
    -- layer=1 filter=143 channel=75
    47, 42, 56, 23, 10, 35, -6, 44, 20,
    -- layer=1 filter=143 channel=76
    26, 10, 14, 1, -47, -18, -30, -6, -20,
    -- layer=1 filter=143 channel=77
    -12, -17, -13, 3, 0, -4, -1, 5, 8,
    -- layer=1 filter=143 channel=78
    -6, -16, 0, -13, -33, -12, 0, -19, 3,
    -- layer=1 filter=143 channel=79
    -73, -94, -93, -102, -75, -68, -13, -40, -16,
    -- layer=1 filter=143 channel=80
    9, 4, -29, -16, -33, 13, -10, -20, -37,
    -- layer=1 filter=143 channel=81
    -32, -22, -17, 0, -5, -2, -7, -6, 14,
    -- layer=1 filter=143 channel=82
    0, 7, -10, 6, 11, 7, 7, 14, 3,
    -- layer=1 filter=143 channel=83
    -33, -33, -22, -38, -44, -71, -40, -39, -59,
    -- layer=1 filter=143 channel=84
    43, 41, 42, 14, -25, -36, -42, -20, -61,
    -- layer=1 filter=143 channel=85
    12, 16, 0, 11, -10, -6, 4, 0, 31,
    -- layer=1 filter=143 channel=86
    16, -11, -2, -2, 5, 7, -6, -10, -10,
    -- layer=1 filter=143 channel=87
    74, 49, 70, 34, 68, 11, -22, 13, 8,
    -- layer=1 filter=143 channel=88
    24, 25, 28, 37, 11, 23, 14, 14, 15,
    -- layer=1 filter=143 channel=89
    5, 10, -1, 11, -3, 10, 0, 17, -9,
    -- layer=1 filter=143 channel=90
    -6, -30, -55, -30, -65, -84, -14, -54, -85,
    -- layer=1 filter=143 channel=91
    41, 18, 27, 14, 15, -2, -1, 10, 11,
    -- layer=1 filter=143 channel=92
    -16, -26, -50, -12, -23, -54, 32, -33, -30,
    -- layer=1 filter=143 channel=93
    -2, 0, -4, -2, -7, 0, 4, -1, -15,
    -- layer=1 filter=143 channel=94
    -19, -16, -6, -42, -33, -39, -25, -33, -50,
    -- layer=1 filter=143 channel=95
    54, 43, 50, -7, -35, -9, -30, -16, -41,
    -- layer=1 filter=143 channel=96
    -19, -15, -13, 11, -4, -22, -12, -15, -20,
    -- layer=1 filter=143 channel=97
    -35, -36, -34, -47, -41, -46, -49, -55, -36,
    -- layer=1 filter=143 channel=98
    -45, -59, -67, -106, -51, -54, -48, -52, -20,
    -- layer=1 filter=143 channel=99
    -32, -51, -18, -107, -61, -59, -90, -36, -35,
    -- layer=1 filter=143 channel=100
    26, -9, 19, 27, 15, 19, 30, 18, 22,
    -- layer=1 filter=143 channel=101
    27, 21, 5, 5, -9, -6, 3, 17, -9,
    -- layer=1 filter=143 channel=102
    -6, -14, -11, -34, -25, -33, -50, -44, -37,
    -- layer=1 filter=143 channel=103
    26, 6, 15, 24, 15, 12, 40, 30, 32,
    -- layer=1 filter=143 channel=104
    76, 14, 31, 19, 4, 4, 10, -1, -19,
    -- layer=1 filter=143 channel=105
    -12, -24, -13, -40, -42, -45, -55, -46, -34,
    -- layer=1 filter=143 channel=106
    37, 22, 9, 0, -8, -23, 9, 4, -9,
    -- layer=1 filter=143 channel=107
    -6, 1, -6, 7, 21, 14, 10, 8, -5,
    -- layer=1 filter=143 channel=108
    25, -1, -16, 15, -29, -37, 27, -4, -46,
    -- layer=1 filter=143 channel=109
    10, 0, 11, -7, -1, 7, 1, 6, -2,
    -- layer=1 filter=143 channel=110
    8, 6, 7, -1, -14, 10, -15, -3, 0,
    -- layer=1 filter=143 channel=111
    50, 52, 53, -8, -38, -33, -84, -43, -79,
    -- layer=1 filter=143 channel=112
    35, 36, 35, -16, -68, -21, -29, -78, -75,
    -- layer=1 filter=143 channel=113
    -18, -3, 5, 4, 8, 17, 34, 32, 24,
    -- layer=1 filter=143 channel=114
    -48, -64, -52, -60, -42, -42, 1, -26, 0,
    -- layer=1 filter=143 channel=115
    -23, -34, -20, -38, -41, -47, -19, -43, -9,
    -- layer=1 filter=143 channel=116
    0, 3, -2, 6, -2, 6, 0, 1, 10,
    -- layer=1 filter=143 channel=117
    38, 39, 35, -51, -71, -51, -97, -105, -101,
    -- layer=1 filter=143 channel=118
    46, 34, 53, 16, -15, -26, -55, -40, -44,
    -- layer=1 filter=143 channel=119
    30, 8, 9, 9, -31, -44, 1, -26, -53,
    -- layer=1 filter=143 channel=120
    20, -10, -3, -13, 6, 0, 15, -2, 22,
    -- layer=1 filter=143 channel=121
    59, 28, 29, 36, 35, 57, 32, 65, 46,
    -- layer=1 filter=143 channel=122
    -6, -4, 6, 1, 2, 8, -5, 7, 5,
    -- layer=1 filter=143 channel=123
    22, 8, 16, 17, 24, 22, 49, 49, 45,
    -- layer=1 filter=143 channel=124
    -21, -8, 0, 2, 4, -3, -11, 9, -3,
    -- layer=1 filter=143 channel=125
    61, 27, 40, -10, -11, -7, 9, 13, 7,
    -- layer=1 filter=143 channel=126
    -60, -41, -62, -74, -49, -69, -71, -61, -17,
    -- layer=1 filter=143 channel=127
    66, 46, 59, 34, -3, -5, -27, -23, -35,
    -- layer=1 filter=144 channel=0
    7, 10, 4, 13, 2, 0, 6, 8, 5,
    -- layer=1 filter=144 channel=1
    -11, -14, -5, 17, 6, 3, 6, -7, -17,
    -- layer=1 filter=144 channel=2
    37, 36, 14, 14, -21, 1, 25, 24, -12,
    -- layer=1 filter=144 channel=3
    -8, 6, 9, 4, 2, 10, 0, 7, 5,
    -- layer=1 filter=144 channel=4
    9, 2, 7, 10, 1, 9, -7, -3, -5,
    -- layer=1 filter=144 channel=5
    19, 14, 19, -6, 15, -6, -2, -34, -27,
    -- layer=1 filter=144 channel=6
    13, 10, 1, -47, -39, 14, -33, 7, 55,
    -- layer=1 filter=144 channel=7
    -1, 17, -31, 13, 33, 4, 20, 34, 22,
    -- layer=1 filter=144 channel=8
    -6, 5, 17, 22, 33, 16, 16, -11, 7,
    -- layer=1 filter=144 channel=9
    6, -10, -4, 17, -53, 7, -33, 63, -15,
    -- layer=1 filter=144 channel=10
    -3, 22, -5, 8, 26, -15, 16, 35, 27,
    -- layer=1 filter=144 channel=11
    -3, -9, -17, 19, 12, -9, 11, 0, -11,
    -- layer=1 filter=144 channel=12
    -1, -3, -13, 20, -28, 0, -32, 26, 37,
    -- layer=1 filter=144 channel=13
    1, -40, -1, -27, 4, 9, 6, 42, 45,
    -- layer=1 filter=144 channel=14
    10, 14, -52, 0, 24, -25, -32, 31, 4,
    -- layer=1 filter=144 channel=15
    -40, -16, -16, -39, -14, 27, 10, 6, 14,
    -- layer=1 filter=144 channel=16
    -1, 4, 12, 6, 20, -5, 26, 16, 14,
    -- layer=1 filter=144 channel=17
    16, -2, 22, 30, 9, 14, 6, 14, 24,
    -- layer=1 filter=144 channel=18
    4, -16, 9, 8, 12, -20, 11, -11, 1,
    -- layer=1 filter=144 channel=19
    17, 27, 10, -47, -13, -43, 5, 12, 6,
    -- layer=1 filter=144 channel=20
    -26, -17, -5, -38, -18, 3, 7, 19, 32,
    -- layer=1 filter=144 channel=21
    -39, -57, -27, -61, -43, -25, -37, -21, -44,
    -- layer=1 filter=144 channel=22
    -12, -29, -4, 16, 13, 23, 16, 34, 52,
    -- layer=1 filter=144 channel=23
    0, 28, 5, 16, 46, 28, 55, 29, 22,
    -- layer=1 filter=144 channel=24
    -15, -37, -7, -54, -9, -34, -11, -25, 0,
    -- layer=1 filter=144 channel=25
    -16, 19, -26, 13, 2, -15, 15, 31, 27,
    -- layer=1 filter=144 channel=26
    4, -44, -17, -33, 22, 16, 15, 29, 34,
    -- layer=1 filter=144 channel=27
    5, 3, -25, 4, -14, -7, -1, -8, -22,
    -- layer=1 filter=144 channel=28
    -21, 7, -25, -6, -2, -30, 8, 33, 29,
    -- layer=1 filter=144 channel=29
    -7, -11, -30, 11, -19, 0, -9, -30, -30,
    -- layer=1 filter=144 channel=30
    2, -25, 17, -25, -14, -23, 2, -20, -4,
    -- layer=1 filter=144 channel=31
    -16, -15, -20, -19, -28, -2, -23, -7, 12,
    -- layer=1 filter=144 channel=32
    -4, -31, -13, -18, 25, 1, 15, 16, 4,
    -- layer=1 filter=144 channel=33
    -8, -1, -3, -3, 9, 2, 33, 4, 12,
    -- layer=1 filter=144 channel=34
    28, 2, -31, 19, 19, 7, -14, 13, 9,
    -- layer=1 filter=144 channel=35
    -16, 0, -14, -13, -4, -15, 0, -11, 1,
    -- layer=1 filter=144 channel=36
    17, 22, 1, 25, 21, 14, 22, 15, 11,
    -- layer=1 filter=144 channel=37
    7, 19, -4, -7, 8, -24, 15, -16, -14,
    -- layer=1 filter=144 channel=38
    -34, -24, -4, -57, -20, -7, -14, 10, 43,
    -- layer=1 filter=144 channel=39
    14, -1, 7, 20, 21, -1, 0, 1, -3,
    -- layer=1 filter=144 channel=40
    -50, -46, -33, -40, -36, -42, -35, 0, 34,
    -- layer=1 filter=144 channel=41
    46, -29, 17, -3, 14, -18, 22, 29, -17,
    -- layer=1 filter=144 channel=42
    26, 32, 25, 19, 24, -8, -2, -19, -22,
    -- layer=1 filter=144 channel=43
    -25, 14, 6, 0, 31, -7, 6, 4, -15,
    -- layer=1 filter=144 channel=44
    -2, -15, -11, -5, 47, 16, 24, 36, 25,
    -- layer=1 filter=144 channel=45
    -21, -32, -17, -58, -9, -12, 0, -13, 8,
    -- layer=1 filter=144 channel=46
    29, 43, 42, -59, -49, -14, 13, 3, -12,
    -- layer=1 filter=144 channel=47
    -3, 34, 8, 14, 10, 33, 24, -1, -14,
    -- layer=1 filter=144 channel=48
    -16, -12, -4, -24, 3, 0, -26, -9, 10,
    -- layer=1 filter=144 channel=49
    -5, -4, -25, -1, -13, -6, -8, 1, -3,
    -- layer=1 filter=144 channel=50
    5, -6, 10, 2, -3, -7, -24, -12, -8,
    -- layer=1 filter=144 channel=51
    -46, -28, -18, -32, -15, -26, -19, 0, 24,
    -- layer=1 filter=144 channel=52
    12, 1, -18, 4, 1, 13, -5, 7, 16,
    -- layer=1 filter=144 channel=53
    8, 7, -9, 1, 8, -6, -11, -15, -14,
    -- layer=1 filter=144 channel=54
    -7, 33, -1, -8, 11, -39, 14, 21, 34,
    -- layer=1 filter=144 channel=55
    17, -7, -34, 30, 11, -13, -4, -42, -42,
    -- layer=1 filter=144 channel=56
    2, 1, -6, -5, -6, -8, 3, 9, 7,
    -- layer=1 filter=144 channel=57
    -14, -8, -29, -5, 5, -7, 5, 29, 40,
    -- layer=1 filter=144 channel=58
    9, 40, 0, 27, 27, 6, 34, 6, 39,
    -- layer=1 filter=144 channel=59
    3, 6, 3, 11, -11, 4, -9, -7, -6,
    -- layer=1 filter=144 channel=60
    -5, -20, -17, -21, -12, -11, -11, -7, -6,
    -- layer=1 filter=144 channel=61
    3, 7, -9, 3, -7, -7, 0, -7, 0,
    -- layer=1 filter=144 channel=62
    6, 0, 7, 1, 28, -20, 12, -3, 11,
    -- layer=1 filter=144 channel=63
    5, 7, -19, 18, -5, -1, 14, 0, -18,
    -- layer=1 filter=144 channel=64
    2, -10, -1, -4, 2, -4, -3, 0, -11,
    -- layer=1 filter=144 channel=65
    -10, -1, 0, -31, -10, 16, -7, -2, 2,
    -- layer=1 filter=144 channel=66
    7, 17, 0, 9, 0, -9, -9, 7, -20,
    -- layer=1 filter=144 channel=67
    -43, -37, -46, -16, -8, -1, -14, 22, -16,
    -- layer=1 filter=144 channel=68
    23, -20, 1, -26, 48, 1, 10, 36, 19,
    -- layer=1 filter=144 channel=69
    4, -14, -6, -36, 15, 8, 24, -1, 3,
    -- layer=1 filter=144 channel=70
    -24, -18, 5, -4, -25, 1, -38, -23, 5,
    -- layer=1 filter=144 channel=71
    -26, 3, -8, -40, 0, -30, -2, 0, -29,
    -- layer=1 filter=144 channel=72
    13, -4, 2, -48, -32, -26, 10, 7, -3,
    -- layer=1 filter=144 channel=73
    -11, -3, 0, -5, 7, -6, -10, 4, -2,
    -- layer=1 filter=144 channel=74
    -3, 20, 20, -26, 3, -7, -12, 7, -10,
    -- layer=1 filter=144 channel=75
    8, -11, -7, -8, -33, -46, -13, 1, 4,
    -- layer=1 filter=144 channel=76
    -3, -8, 0, -22, 10, 14, -8, 21, 0,
    -- layer=1 filter=144 channel=77
    -27, -33, -12, -5, 1, -1, -25, -19, -3,
    -- layer=1 filter=144 channel=78
    4, 7, 1, -4, 2, -2, 1, 25, -5,
    -- layer=1 filter=144 channel=79
    1, -4, 0, 15, 6, -1, 30, 4, 13,
    -- layer=1 filter=144 channel=80
    1, 5, 0, 9, 1, 0, 6, -1, 9,
    -- layer=1 filter=144 channel=81
    -20, -23, -22, 3, 7, -19, -5, -26, -18,
    -- layer=1 filter=144 channel=82
    -70, -56, -23, -46, -37, 6, -46, -46, -12,
    -- layer=1 filter=144 channel=83
    0, -24, 6, 0, 9, 3, 5, -10, 33,
    -- layer=1 filter=144 channel=84
    -18, -23, 19, 8, 23, -15, 2, 11, -3,
    -- layer=1 filter=144 channel=85
    0, 28, 16, 27, 54, 24, 24, 22, 23,
    -- layer=1 filter=144 channel=86
    1, 17, 0, 20, 5, -4, 14, 6, 0,
    -- layer=1 filter=144 channel=87
    11, 35, 31, 30, -2, -11, -25, 32, -26,
    -- layer=1 filter=144 channel=88
    -30, -2, -19, -16, -21, -19, 1, -12, 1,
    -- layer=1 filter=144 channel=89
    -54, -29, -23, -34, -18, -10, -32, -8, -19,
    -- layer=1 filter=144 channel=90
    28, -27, -17, -26, 21, 13, 19, 6, 25,
    -- layer=1 filter=144 channel=91
    -30, -32, -21, -32, -38, 1, -21, -20, 24,
    -- layer=1 filter=144 channel=92
    26, -4, -20, -27, 2, 18, -10, 19, -9,
    -- layer=1 filter=144 channel=93
    -13, -15, 2, -3, 0, 4, -13, -20, -2,
    -- layer=1 filter=144 channel=94
    11, 21, 11, 21, 12, 20, 16, 8, 0,
    -- layer=1 filter=144 channel=95
    -6, -1, 33, 1, 19, -5, -18, 25, -2,
    -- layer=1 filter=144 channel=96
    10, 15, -1, 4, 14, 18, 5, 13, 13,
    -- layer=1 filter=144 channel=97
    -2, 4, -5, 21, 18, 14, -5, 5, -5,
    -- layer=1 filter=144 channel=98
    -15, -15, 5, 32, 37, -1, 7, 12, 7,
    -- layer=1 filter=144 channel=99
    -29, -26, -16, -10, 1, 10, 8, 36, 28,
    -- layer=1 filter=144 channel=100
    5, 4, 1, 6, 12, 0, 7, 2, -16,
    -- layer=1 filter=144 channel=101
    -42, -22, -5, -21, -28, 14, -29, -7, 14,
    -- layer=1 filter=144 channel=102
    0, 25, 30, 3, 17, 12, 13, 9, 12,
    -- layer=1 filter=144 channel=103
    19, -4, -19, 6, -3, -11, -7, -20, -18,
    -- layer=1 filter=144 channel=104
    -15, 8, -3, 21, 10, 30, 29, 28, 2,
    -- layer=1 filter=144 channel=105
    4, 11, 0, 15, 3, 4, -6, 4, -11,
    -- layer=1 filter=144 channel=106
    -44, -33, -17, -40, -17, -6, -20, 30, 12,
    -- layer=1 filter=144 channel=107
    6, 0, -3, 17, 7, 15, 17, 6, 2,
    -- layer=1 filter=144 channel=108
    0, -62, -1, -27, 25, 33, 16, 8, 23,
    -- layer=1 filter=144 channel=109
    1, -8, 6, -5, 3, -1, -7, -5, 0,
    -- layer=1 filter=144 channel=110
    -8, -7, -2, 0, 9, -6, -13, 1, -5,
    -- layer=1 filter=144 channel=111
    0, -18, 31, 10, 32, -13, -17, -1, -8,
    -- layer=1 filter=144 channel=112
    -3, 5, 11, 48, 34, 15, -2, -7, 1,
    -- layer=1 filter=144 channel=113
    10, 26, 23, 12, 20, 13, 13, 20, 50,
    -- layer=1 filter=144 channel=114
    2, 8, -5, -13, 17, -9, 24, -28, -24,
    -- layer=1 filter=144 channel=115
    1, 28, 3, 13, 24, -2, 20, 6, 8,
    -- layer=1 filter=144 channel=116
    10, -2, -6, 6, -1, -5, 1, -2, 0,
    -- layer=1 filter=144 channel=117
    -22, 11, 25, 33, 25, 8, -28, -28, -11,
    -- layer=1 filter=144 channel=118
    -14, -12, 11, -22, -15, -15, -19, 0, -16,
    -- layer=1 filter=144 channel=119
    23, -45, -4, -31, 20, 0, 18, 4, 24,
    -- layer=1 filter=144 channel=120
    -43, -26, -35, -9, -22, -17, -4, -10, 7,
    -- layer=1 filter=144 channel=121
    5, -6, -25, -22, -46, -39, -7, 5, -9,
    -- layer=1 filter=144 channel=122
    5, -10, -5, 6, -10, 5, -10, 8, 1,
    -- layer=1 filter=144 channel=123
    18, 1, -31, -1, -27, -30, 17, -16, -24,
    -- layer=1 filter=144 channel=124
    -15, -15, -17, 5, -4, -8, -12, -5, -7,
    -- layer=1 filter=144 channel=125
    -22, -23, -25, -77, -34, -11, -26, -2, 54,
    -- layer=1 filter=144 channel=126
    -14, -27, -9, 49, 48, 11, -37, -38, 7,
    -- layer=1 filter=144 channel=127
    -11, -12, 26, -9, -9, -7, -6, 7, -10,
    -- layer=1 filter=145 channel=0
    -1, 0, -2, -3, 1, -3, 2, 7, -11,
    -- layer=1 filter=145 channel=1
    3, -4, 8, 0, -12, -9, 5, 1, 5,
    -- layer=1 filter=145 channel=2
    -10, 7, -2, 2, 6, -9, 0, 3, -10,
    -- layer=1 filter=145 channel=3
    -8, 0, -10, 1, 2, 9, -6, -5, -7,
    -- layer=1 filter=145 channel=4
    -5, 0, 4, 4, 2, 0, 0, 1, 7,
    -- layer=1 filter=145 channel=5
    -10, -6, 7, -4, 9, 1, -7, -2, -1,
    -- layer=1 filter=145 channel=6
    -11, 1, 5, -10, -1, -4, -7, -7, 6,
    -- layer=1 filter=145 channel=7
    7, 0, -2, 1, -1, 11, 2, -10, -10,
    -- layer=1 filter=145 channel=8
    0, -7, -3, 1, -5, -4, 0, -1, -6,
    -- layer=1 filter=145 channel=9
    5, -1, 4, -1, 6, 1, -6, -9, 6,
    -- layer=1 filter=145 channel=10
    0, -10, 7, 7, -5, -10, 7, 3, -11,
    -- layer=1 filter=145 channel=11
    6, 6, 2, -7, 9, 6, 9, -2, -1,
    -- layer=1 filter=145 channel=12
    -4, -4, -7, -8, 8, 4, 5, 4, 2,
    -- layer=1 filter=145 channel=13
    6, 0, -8, -9, 3, 7, -1, 7, 3,
    -- layer=1 filter=145 channel=14
    3, -10, -3, 4, 4, -2, -6, -10, 6,
    -- layer=1 filter=145 channel=15
    -2, -9, 5, 0, 0, -7, 4, 0, -11,
    -- layer=1 filter=145 channel=16
    -2, 7, -7, 3, -8, -3, -1, -9, -8,
    -- layer=1 filter=145 channel=17
    -3, 1, 4, -4, 0, -3, -7, 0, -6,
    -- layer=1 filter=145 channel=18
    -5, -8, 0, 6, 0, -11, 0, -2, -2,
    -- layer=1 filter=145 channel=19
    -6, -3, 0, -4, -5, -3, 3, -5, -7,
    -- layer=1 filter=145 channel=20
    -10, -6, 7, -2, -10, -10, 7, -11, -3,
    -- layer=1 filter=145 channel=21
    -1, -10, 4, -1, -9, 0, 0, 1, -11,
    -- layer=1 filter=145 channel=22
    -5, -5, 5, 5, 1, 8, -9, 6, 5,
    -- layer=1 filter=145 channel=23
    -4, 7, 0, -10, 0, 7, 0, -10, 8,
    -- layer=1 filter=145 channel=24
    0, -6, 6, -1, -4, -7, 6, 4, -1,
    -- layer=1 filter=145 channel=25
    -11, -9, -9, 4, 1, 8, 3, -4, 10,
    -- layer=1 filter=145 channel=26
    -14, 2, -3, 3, -10, 5, 3, 6, -8,
    -- layer=1 filter=145 channel=27
    -7, -2, 3, 1, 1, -10, -8, -3, -7,
    -- layer=1 filter=145 channel=28
    0, 0, -10, 8, -1, -6, -10, -12, -12,
    -- layer=1 filter=145 channel=29
    6, -8, -8, 8, -2, 0, 5, -6, 5,
    -- layer=1 filter=145 channel=30
    -4, 0, -1, -10, -3, 8, 6, -7, 8,
    -- layer=1 filter=145 channel=31
    0, -1, -4, 0, 5, 3, 10, 0, 7,
    -- layer=1 filter=145 channel=32
    2, -8, 0, -5, 3, -9, -1, -11, -10,
    -- layer=1 filter=145 channel=33
    -1, -3, 0, -8, -1, -6, 0, 8, -3,
    -- layer=1 filter=145 channel=34
    0, -3, -6, -3, 5, 3, -3, 0, 7,
    -- layer=1 filter=145 channel=35
    -9, -10, -8, -3, 0, -10, -12, -2, -11,
    -- layer=1 filter=145 channel=36
    5, -10, 6, -5, 0, 0, 5, -8, -8,
    -- layer=1 filter=145 channel=37
    1, 0, 3, 4, -3, 3, -7, 0, 5,
    -- layer=1 filter=145 channel=38
    -2, -9, -10, 0, -7, -9, -3, 3, -9,
    -- layer=1 filter=145 channel=39
    8, 5, 1, 5, -1, -6, 0, -3, 3,
    -- layer=1 filter=145 channel=40
    -5, 5, -1, -7, 0, -1, 1, -2, -8,
    -- layer=1 filter=145 channel=41
    -7, 3, 3, 0, 9, -8, -2, 4, -2,
    -- layer=1 filter=145 channel=42
    6, 0, 4, 9, -6, 3, 7, -2, -1,
    -- layer=1 filter=145 channel=43
    -9, 1, 0, -2, -7, 0, 1, 2, 0,
    -- layer=1 filter=145 channel=44
    -9, -11, 8, 4, -6, -2, 7, 7, 1,
    -- layer=1 filter=145 channel=45
    -3, -9, -12, 3, 0, -4, 7, 0, 0,
    -- layer=1 filter=145 channel=46
    -6, 8, -3, -5, -1, -3, -1, -8, -8,
    -- layer=1 filter=145 channel=47
    1, -9, -3, -11, -3, 4, 0, 2, -12,
    -- layer=1 filter=145 channel=48
    -9, 6, 0, 7, -10, -11, -9, 3, 1,
    -- layer=1 filter=145 channel=49
    0, 7, -9, 0, -8, -8, 0, -8, -3,
    -- layer=1 filter=145 channel=50
    -8, 4, 7, -8, 0, -1, -7, 5, -2,
    -- layer=1 filter=145 channel=51
    -1, 5, 7, 0, -7, -3, -8, 2, 4,
    -- layer=1 filter=145 channel=52
    -9, 8, -10, -6, 0, -11, 0, -4, -6,
    -- layer=1 filter=145 channel=53
    -8, -9, 7, 2, -10, -1, 7, 5, -5,
    -- layer=1 filter=145 channel=54
    -8, 0, -2, 9, 2, 4, 4, 6, -7,
    -- layer=1 filter=145 channel=55
    -5, 11, -7, -10, 10, -9, -4, -1, -2,
    -- layer=1 filter=145 channel=56
    3, 6, -3, 8, -10, -6, 1, 9, 0,
    -- layer=1 filter=145 channel=57
    -6, 8, -10, 8, 0, -5, 2, -1, 6,
    -- layer=1 filter=145 channel=58
    -9, -4, -13, 8, 3, 0, -10, 7, 3,
    -- layer=1 filter=145 channel=59
    -5, -12, 0, -9, 4, -2, -2, -11, -6,
    -- layer=1 filter=145 channel=60
    4, 8, 0, 6, 2, 10, -5, 9, -3,
    -- layer=1 filter=145 channel=61
    1, -5, -4, -4, 8, -3, -1, -10, 11,
    -- layer=1 filter=145 channel=62
    7, 2, 7, -12, -10, 3, -9, -6, -1,
    -- layer=1 filter=145 channel=63
    3, -7, 0, 0, -2, 1, 8, 8, -6,
    -- layer=1 filter=145 channel=64
    6, 4, 0, -1, -4, 2, 0, 0, 3,
    -- layer=1 filter=145 channel=65
    0, 3, 5, 6, -4, 3, -12, 6, 5,
    -- layer=1 filter=145 channel=66
    -8, -11, -10, -9, -2, 7, -8, -8, -12,
    -- layer=1 filter=145 channel=67
    4, -12, 6, -11, -9, -3, 0, 0, 4,
    -- layer=1 filter=145 channel=68
    -2, -4, 1, -7, 6, -5, 0, -7, 0,
    -- layer=1 filter=145 channel=69
    2, -7, -8, 1, -8, 1, -5, -1, -2,
    -- layer=1 filter=145 channel=70
    -9, 1, 0, -3, -9, 1, 9, 6, 2,
    -- layer=1 filter=145 channel=71
    3, -2, 2, -2, -9, 3, 6, -8, -1,
    -- layer=1 filter=145 channel=72
    -3, 3, 0, 7, 4, 8, 5, 0, -3,
    -- layer=1 filter=145 channel=73
    -1, 0, 8, 2, -9, -5, -12, -4, 2,
    -- layer=1 filter=145 channel=74
    -2, 7, -3, -2, 3, 1, 2, -5, 1,
    -- layer=1 filter=145 channel=75
    -8, -5, 9, 0, -6, -1, -10, -10, -4,
    -- layer=1 filter=145 channel=76
    -6, 2, -8, 8, -12, -7, -4, 7, 0,
    -- layer=1 filter=145 channel=77
    0, -9, 8, 7, 1, -11, 4, -2, -7,
    -- layer=1 filter=145 channel=78
    7, -4, 6, -4, 8, 4, -8, -9, -12,
    -- layer=1 filter=145 channel=79
    3, -3, -4, -1, -4, 6, 1, 0, 0,
    -- layer=1 filter=145 channel=80
    -8, -6, -5, -9, 5, -9, 5, 0, -8,
    -- layer=1 filter=145 channel=81
    8, -9, 2, -11, 6, 5, -10, 4, 8,
    -- layer=1 filter=145 channel=82
    0, 7, 6, 3, -6, -1, -6, -7, 7,
    -- layer=1 filter=145 channel=83
    8, 8, -10, 6, 5, 3, 5, -8, 5,
    -- layer=1 filter=145 channel=84
    -7, 2, -9, -8, -6, 5, -2, 3, 6,
    -- layer=1 filter=145 channel=85
    -6, -4, 6, 3, 4, 9, 8, -4, -10,
    -- layer=1 filter=145 channel=86
    -4, 6, -2, 0, 6, -8, -5, -5, -8,
    -- layer=1 filter=145 channel=87
    -6, 0, -5, 3, 4, -9, -3, -6, 2,
    -- layer=1 filter=145 channel=88
    2, 0, -5, -10, 8, -8, -4, 6, -7,
    -- layer=1 filter=145 channel=89
    -10, 4, -4, -4, -11, 3, 5, -6, -6,
    -- layer=1 filter=145 channel=90
    -7, 0, -12, 5, -5, -2, 0, -12, 2,
    -- layer=1 filter=145 channel=91
    -8, 0, 1, 2, 3, 7, -10, 0, 2,
    -- layer=1 filter=145 channel=92
    0, -10, 3, -11, -3, -1, 5, -7, 8,
    -- layer=1 filter=145 channel=93
    -2, -6, 0, -9, -7, -2, -7, -4, 8,
    -- layer=1 filter=145 channel=94
    -2, -8, -2, -8, 6, 3, -4, -6, 5,
    -- layer=1 filter=145 channel=95
    0, 6, 1, 0, -1, 3, -11, 6, 0,
    -- layer=1 filter=145 channel=96
    -9, -1, -11, -5, -11, -7, 5, -8, -8,
    -- layer=1 filter=145 channel=97
    2, -12, 7, 0, -6, -5, 5, 7, -3,
    -- layer=1 filter=145 channel=98
    -9, -9, 4, 2, -8, -9, -2, -10, 0,
    -- layer=1 filter=145 channel=99
    6, 2, 4, 2, -8, -5, 0, -7, 2,
    -- layer=1 filter=145 channel=100
    4, -10, -2, 1, 0, -3, -1, -10, 4,
    -- layer=1 filter=145 channel=101
    6, 1, 5, 1, 5, -1, -1, 8, 4,
    -- layer=1 filter=145 channel=102
    -9, -6, 0, -1, 8, -7, -3, -8, 8,
    -- layer=1 filter=145 channel=103
    -7, -8, -3, 2, -6, -8, -3, -4, -8,
    -- layer=1 filter=145 channel=104
    2, -10, 5, 6, -1, -1, -6, -2, 8,
    -- layer=1 filter=145 channel=105
    8, 0, 4, -1, -5, -10, -3, -6, 7,
    -- layer=1 filter=145 channel=106
    -11, -9, -3, 6, -4, 7, 1, -10, -7,
    -- layer=1 filter=145 channel=107
    -5, -10, -2, -2, 2, 3, -1, -3, -5,
    -- layer=1 filter=145 channel=108
    4, 0, -9, -12, -6, 8, 1, -9, -9,
    -- layer=1 filter=145 channel=109
    -2, 1, 2, -5, -9, -5, 0, 7, -2,
    -- layer=1 filter=145 channel=110
    6, -3, 2, 8, -6, -12, -3, -8, 3,
    -- layer=1 filter=145 channel=111
    5, -9, -1, -6, 3, -5, -7, 1, -3,
    -- layer=1 filter=145 channel=112
    2, 1, -9, 0, -3, 4, -6, 0, 1,
    -- layer=1 filter=145 channel=113
    -3, 3, 4, 6, -11, 1, -2, 0, -6,
    -- layer=1 filter=145 channel=114
    -1, -7, -7, -10, 7, 4, 3, -7, -9,
    -- layer=1 filter=145 channel=115
    -9, -3, 2, -5, -8, 4, 3, 4, 2,
    -- layer=1 filter=145 channel=116
    5, -5, 5, 0, 1, 6, 1, -3, -3,
    -- layer=1 filter=145 channel=117
    -3, 2, -3, -9, 3, 8, 0, -8, -9,
    -- layer=1 filter=145 channel=118
    -8, 6, 3, 4, 1, -2, -6, 7, -5,
    -- layer=1 filter=145 channel=119
    -12, -5, -2, -7, 7, 8, 5, -8, 3,
    -- layer=1 filter=145 channel=120
    -2, 6, 2, -12, -3, -4, 3, -10, 6,
    -- layer=1 filter=145 channel=121
    3, 9, -3, -5, 0, 6, -3, -7, -6,
    -- layer=1 filter=145 channel=122
    -4, 0, 0, 3, 8, -3, 4, -9, -4,
    -- layer=1 filter=145 channel=123
    4, -6, 2, 5, -11, 3, 3, -3, -12,
    -- layer=1 filter=145 channel=124
    5, -1, -2, 2, -1, 7, 6, -2, 5,
    -- layer=1 filter=145 channel=125
    8, -1, 0, -2, -8, 8, 5, -7, 3,
    -- layer=1 filter=145 channel=126
    -11, -7, 3, 8, -2, 0, 7, -5, -6,
    -- layer=1 filter=145 channel=127
    6, 4, -1, 0, 8, -1, 0, 2, -10,
    -- layer=1 filter=146 channel=0
    -13, -9, 1, -17, -2, -15, -29, 0, -8,
    -- layer=1 filter=146 channel=1
    -39, 14, 0, -48, -43, -4, 10, -9, 0,
    -- layer=1 filter=146 channel=2
    49, 28, 2, 45, 10, -2, 34, 15, 1,
    -- layer=1 filter=146 channel=3
    0, -1, 10, -9, -8, 8, -6, 13, 7,
    -- layer=1 filter=146 channel=4
    6, 2, -3, -3, -13, -13, -18, -6, -14,
    -- layer=1 filter=146 channel=5
    -74, -16, -24, -44, -16, 17, 13, 5, 23,
    -- layer=1 filter=146 channel=6
    24, 29, 16, 41, 34, 20, 11, -5, -21,
    -- layer=1 filter=146 channel=7
    -8, 17, 37, -13, 6, 35, -6, 31, -5,
    -- layer=1 filter=146 channel=8
    -26, 5, -12, -46, -50, -25, 7, -7, -4,
    -- layer=1 filter=146 channel=9
    7, 26, -29, 13, -12, -11, -37, -33, -3,
    -- layer=1 filter=146 channel=10
    3, 3, 25, -3, 24, 8, -2, 53, 15,
    -- layer=1 filter=146 channel=11
    14, -37, -26, 31, 11, -15, 28, 44, 5,
    -- layer=1 filter=146 channel=12
    -64, 17, -38, -28, -32, 22, -5, -16, -28,
    -- layer=1 filter=146 channel=13
    21, 36, -1, 9, 16, 2, -5, -23, -36,
    -- layer=1 filter=146 channel=14
    -46, -40, 4, -62, -45, -16, -1, 0, -35,
    -- layer=1 filter=146 channel=15
    -24, 9, -7, -9, -24, -19, 12, -14, 30,
    -- layer=1 filter=146 channel=16
    -48, 24, -11, -60, -33, -15, -15, -3, -11,
    -- layer=1 filter=146 channel=17
    33, -9, 24, -5, -32, -47, -35, -49, -49,
    -- layer=1 filter=146 channel=18
    -68, -35, -9, -44, -17, -7, -30, 7, -23,
    -- layer=1 filter=146 channel=19
    -88, -41, -26, -68, -32, -45, -14, -36, 17,
    -- layer=1 filter=146 channel=20
    20, 46, 23, 10, 26, 7, 0, -23, -30,
    -- layer=1 filter=146 channel=21
    -27, -8, 15, -14, 4, 5, 1, 8, 2,
    -- layer=1 filter=146 channel=22
    41, 45, 13, 11, 6, -8, -6, -20, -42,
    -- layer=1 filter=146 channel=23
    -32, 35, -14, -17, -48, -18, 50, 22, 16,
    -- layer=1 filter=146 channel=24
    -28, -73, -76, -32, -32, -47, 15, -32, 13,
    -- layer=1 filter=146 channel=25
    -23, 30, 17, -21, 16, 19, -11, 22, -13,
    -- layer=1 filter=146 channel=26
    35, -1, -14, 6, -56, -16, 20, -46, -18,
    -- layer=1 filter=146 channel=27
    70, 13, -18, 54, 1, -30, 66, 35, -1,
    -- layer=1 filter=146 channel=28
    -45, -4, 18, -44, -13, 12, -49, 17, -22,
    -- layer=1 filter=146 channel=29
    29, -21, 3, 48, 19, 24, 34, 18, -8,
    -- layer=1 filter=146 channel=30
    -57, -28, 4, -16, -20, 14, -5, -16, -28,
    -- layer=1 filter=146 channel=31
    5, 24, 10, 33, 34, 31, 17, 20, 6,
    -- layer=1 filter=146 channel=32
    3, -21, -28, 41, -20, 25, 49, 18, 13,
    -- layer=1 filter=146 channel=33
    -6, -17, -13, -23, -29, -18, 3, -14, -7,
    -- layer=1 filter=146 channel=34
    -44, -64, -44, -37, -52, -41, -5, -25, -44,
    -- layer=1 filter=146 channel=35
    0, 7, 12, 13, -4, 9, 4, -31, 27,
    -- layer=1 filter=146 channel=36
    2, -52, -27, 30, 0, -34, 27, 34, 17,
    -- layer=1 filter=146 channel=37
    -83, -1, -7, -41, 19, 8, 12, 48, 49,
    -- layer=1 filter=146 channel=38
    31, 33, 22, 2, 32, 1, 0, -5, -27,
    -- layer=1 filter=146 channel=39
    5, -12, -24, -2, -22, -39, -4, -2, 4,
    -- layer=1 filter=146 channel=40
    37, 45, 33, 35, 45, 38, 4, 18, -6,
    -- layer=1 filter=146 channel=41
    -24, -21, -44, 9, -45, -17, 7, -6, 3,
    -- layer=1 filter=146 channel=42
    62, 39, 20, 32, 44, -7, 2, 31, -11,
    -- layer=1 filter=146 channel=43
    -40, 20, -16, -47, -37, -2, -15, 14, -9,
    -- layer=1 filter=146 channel=44
    31, -19, -15, 33, -41, -9, 46, -8, 12,
    -- layer=1 filter=146 channel=45
    -7, 0, -7, -5, -19, -17, 21, -6, 13,
    -- layer=1 filter=146 channel=46
    -39, -46, -37, -46, -35, -27, 28, -11, 6,
    -- layer=1 filter=146 channel=47
    -19, 10, -1, 14, 10, 16, 47, 46, 14,
    -- layer=1 filter=146 channel=48
    11, 14, 16, -2, 6, -7, -15, 11, -9,
    -- layer=1 filter=146 channel=49
    23, 29, 8, 38, 24, 10, 30, 4, 4,
    -- layer=1 filter=146 channel=50
    -15, -9, -15, -11, -7, -9, -19, -30, -5,
    -- layer=1 filter=146 channel=51
    9, 18, 17, 3, 23, -3, -11, 11, -19,
    -- layer=1 filter=146 channel=52
    -1, 5, -5, 12, -9, -12, -11, -1, 0,
    -- layer=1 filter=146 channel=53
    3, -15, -21, -1, -4, -14, -6, 3, -12,
    -- layer=1 filter=146 channel=54
    -28, -3, 16, 9, 1, 25, 3, 29, 10,
    -- layer=1 filter=146 channel=55
    -11, -66, -60, -6, -28, -9, 21, 30, 34,
    -- layer=1 filter=146 channel=56
    -3, 10, 7, -7, 0, -3, -7, 1, 10,
    -- layer=1 filter=146 channel=57
    39, 38, 53, 6, 51, 10, -8, 42, -6,
    -- layer=1 filter=146 channel=58
    5, 42, 10, -15, 17, -23, 60, 60, 24,
    -- layer=1 filter=146 channel=59
    3, -12, -2, -15, -15, 6, -24, -8, -22,
    -- layer=1 filter=146 channel=60
    -10, -19, -18, -10, -17, 2, -3, -7, 9,
    -- layer=1 filter=146 channel=61
    4, 7, 7, -1, -12, -10, 8, 11, -19,
    -- layer=1 filter=146 channel=62
    -27, 21, -22, -60, -28, -38, -20, -19, 1,
    -- layer=1 filter=146 channel=63
    -30, -59, -39, -11, -41, -23, 7, 31, 0,
    -- layer=1 filter=146 channel=64
    -6, 25, 11, -11, 0, -11, -20, -20, -7,
    -- layer=1 filter=146 channel=65
    -7, 21, 15, -4, 1, 8, -19, -21, -8,
    -- layer=1 filter=146 channel=66
    -12, -35, -14, 8, -34, -11, 30, -1, 15,
    -- layer=1 filter=146 channel=67
    7, 18, 33, 0, 44, 22, 14, 0, -4,
    -- layer=1 filter=146 channel=68
    28, -25, -15, 30, -51, 13, 43, 2, 23,
    -- layer=1 filter=146 channel=69
    -31, -15, -14, -41, -53, -38, 7, -22, 16,
    -- layer=1 filter=146 channel=70
    -6, -5, 3, 14, 29, 33, 1, 13, -9,
    -- layer=1 filter=146 channel=71
    -60, -62, -42, -43, -58, -35, -20, -9, -14,
    -- layer=1 filter=146 channel=72
    -62, -18, -36, -49, -62, -13, -53, -66, -54,
    -- layer=1 filter=146 channel=73
    -3, -8, -4, -7, 3, 0, -8, -14, 4,
    -- layer=1 filter=146 channel=74
    34, 8, -6, 7, 12, 41, 18, 8, 26,
    -- layer=1 filter=146 channel=75
    -94, -29, -12, -51, -74, -13, -63, -44, -68,
    -- layer=1 filter=146 channel=76
    0, -16, -15, 17, -22, 8, 13, -20, -16,
    -- layer=1 filter=146 channel=77
    -46, -9, 1, -49, -9, 0, 12, 15, 24,
    -- layer=1 filter=146 channel=78
    -11, -22, -18, -22, -16, 0, -26, 0, -23,
    -- layer=1 filter=146 channel=79
    -32, 34, -14, -43, -33, -39, -11, -23, -7,
    -- layer=1 filter=146 channel=80
    2, -9, 0, 21, 9, 24, -12, 30, 25,
    -- layer=1 filter=146 channel=81
    -82, -59, -35, -99, -104, -52, -8, -22, 21,
    -- layer=1 filter=146 channel=82
    -4, 5, 19, -5, 15, -1, -8, 16, 8,
    -- layer=1 filter=146 channel=83
    -23, -3, 4, -17, -74, -10, 12, -33, 20,
    -- layer=1 filter=146 channel=84
    9, -15, -16, 20, -17, 23, 8, 2, -12,
    -- layer=1 filter=146 channel=85
    -27, 30, 13, -29, 15, -39, 20, 24, 19,
    -- layer=1 filter=146 channel=86
    8, -20, -9, -4, -28, -20, -8, -9, -13,
    -- layer=1 filter=146 channel=87
    -10, 8, 6, -36, -4, 4, 2, -22, 43,
    -- layer=1 filter=146 channel=88
    9, 19, -5, 18, 25, -9, 10, 4, 7,
    -- layer=1 filter=146 channel=89
    9, 13, 3, 2, 1, 4, 12, -11, -1,
    -- layer=1 filter=146 channel=90
    0, -41, -4, 0, -69, -2, 41, -20, 41,
    -- layer=1 filter=146 channel=91
    13, 38, 36, 23, 26, 28, -14, -1, -24,
    -- layer=1 filter=146 channel=92
    4, -9, -26, -2, -34, -11, 16, 1, 55,
    -- layer=1 filter=146 channel=93
    -19, -22, -14, -20, -20, -25, -3, -8, -7,
    -- layer=1 filter=146 channel=94
    -19, -6, 6, -9, -22, -4, -35, -26, -18,
    -- layer=1 filter=146 channel=95
    -27, -9, -13, 2, -31, 17, -1, -26, -41,
    -- layer=1 filter=146 channel=96
    -23, -11, -33, -11, -9, -14, 22, 25, 33,
    -- layer=1 filter=146 channel=97
    -15, -23, -5, -48, -31, -24, -26, -22, -17,
    -- layer=1 filter=146 channel=98
    2, 39, 13, -49, -34, -28, -29, 10, -22,
    -- layer=1 filter=146 channel=99
    -10, -40, 15, -19, -5, -5, -15, 33, 20,
    -- layer=1 filter=146 channel=100
    0, -22, -37, -4, -3, -1, 28, 21, 0,
    -- layer=1 filter=146 channel=101
    23, 39, 23, 7, 15, 18, -7, -7, -26,
    -- layer=1 filter=146 channel=102
    5, 19, 33, -16, 7, 16, -49, -36, -29,
    -- layer=1 filter=146 channel=103
    19, -3, -8, 29, 8, -2, 14, 50, 23,
    -- layer=1 filter=146 channel=104
    -15, 35, 14, -17, -17, -2, 5, 3, 9,
    -- layer=1 filter=146 channel=105
    -19, -31, 7, -36, -30, -13, -43, -6, 4,
    -- layer=1 filter=146 channel=106
    42, 36, 18, 44, 14, 13, 34, -16, -9,
    -- layer=1 filter=146 channel=107
    5, 0, 1, 3, 11, -2, -14, 1, -16,
    -- layer=1 filter=146 channel=108
    7, -35, -46, 25, -65, -35, 46, -11, 0,
    -- layer=1 filter=146 channel=109
    -8, 7, 0, -10, -9, 0, -10, 0, -8,
    -- layer=1 filter=146 channel=110
    -15, 2, -2, 2, 7, -2, -4, -7, 0,
    -- layer=1 filter=146 channel=111
    -26, -30, -3, -41, -16, -2, -13, -8, -39,
    -- layer=1 filter=146 channel=112
    -39, -32, -12, -31, -29, 16, -15, -14, -12,
    -- layer=1 filter=146 channel=113
    14, 7, -14, 15, 17, -17, -7, 16, -28,
    -- layer=1 filter=146 channel=114
    -3, -34, 8, -12, -8, 52, 42, 20, 34,
    -- layer=1 filter=146 channel=115
    -7, 11, 19, -7, -15, -18, -31, -10, -18,
    -- layer=1 filter=146 channel=116
    0, -3, 6, 6, 4, -9, 8, 7, -3,
    -- layer=1 filter=146 channel=117
    -63, -71, -30, -72, -31, -18, -45, -3, -14,
    -- layer=1 filter=146 channel=118
    -6, -8, 11, 1, 13, 46, 23, 0, -2,
    -- layer=1 filter=146 channel=119
    0, -49, -49, 18, -58, -14, 41, 0, 7,
    -- layer=1 filter=146 channel=120
    -17, 24, 23, -21, 8, 3, -7, 18, -2,
    -- layer=1 filter=146 channel=121
    -68, -64, -32, -72, -56, -24, -21, -27, -42,
    -- layer=1 filter=146 channel=122
    9, 9, -3, -5, -1, 9, 4, -1, -7,
    -- layer=1 filter=146 channel=123
    -33, -62, -39, -31, -66, -26, 13, 23, -7,
    -- layer=1 filter=146 channel=124
    3, -1, 6, 10, 2, 0, -4, 13, 9,
    -- layer=1 filter=146 channel=125
    14, 0, -10, 0, 41, 5, 0, 15, -4,
    -- layer=1 filter=146 channel=126
    -49, 6, -2, -99, -39, -37, 12, 36, 46,
    -- layer=1 filter=146 channel=127
    -25, 0, 19, 2, 15, 33, 6, 14, 4,
    -- layer=1 filter=147 channel=0
    13, 0, 7, -4, 5, -7, 0, -20, -20,
    -- layer=1 filter=147 channel=1
    1, -2, 15, 43, 16, -7, -18, -12, 15,
    -- layer=1 filter=147 channel=2
    15, -14, -11, 9, -10, -8, 28, -16, -16,
    -- layer=1 filter=147 channel=3
    9, -12, -13, -8, -10, 3, 10, 0, 5,
    -- layer=1 filter=147 channel=4
    9, 14, 8, -8, 5, -7, -3, 8, 8,
    -- layer=1 filter=147 channel=5
    -31, 12, -3, 30, 3, -15, -50, 4, 7,
    -- layer=1 filter=147 channel=6
    -9, -8, 1, -17, -2, -4, 30, 4, -13,
    -- layer=1 filter=147 channel=7
    -33, -13, 3, 34, -28, -43, -20, -2, 29,
    -- layer=1 filter=147 channel=8
    -18, 8, 9, 53, 0, 0, -32, -1, 23,
    -- layer=1 filter=147 channel=9
    34, 42, 5, 36, -17, 1, 29, 17, -5,
    -- layer=1 filter=147 channel=10
    -38, -22, -12, 26, -6, -16, -37, 23, 22,
    -- layer=1 filter=147 channel=11
    -4, 9, 19, 8, 10, 10, -1, -12, -8,
    -- layer=1 filter=147 channel=12
    -22, -62, -56, -29, -55, -55, -21, -17, -1,
    -- layer=1 filter=147 channel=13
    -5, -3, -4, -1, 0, 20, 13, 0, -4,
    -- layer=1 filter=147 channel=14
    -46, -33, -5, -22, -27, -37, -19, -2, -13,
    -- layer=1 filter=147 channel=15
    -28, -55, -21, -20, -58, -36, -36, -36, -32,
    -- layer=1 filter=147 channel=16
    1, 14, 13, 49, 10, -19, -30, 15, 0,
    -- layer=1 filter=147 channel=17
    -7, -8, -6, -5, -1, -16, -8, -16, -24,
    -- layer=1 filter=147 channel=18
    8, -11, -9, -21, 2, 13, -3, 2, -29,
    -- layer=1 filter=147 channel=19
    79, 115, 25, 129, 60, 75, 51, 116, 33,
    -- layer=1 filter=147 channel=20
    -7, -3, 13, 19, 9, 13, -8, -10, 7,
    -- layer=1 filter=147 channel=21
    6, 13, 14, 4, 4, -6, -12, -39, -9,
    -- layer=1 filter=147 channel=22
    -18, 8, 11, 21, 24, 8, -1, 4, 12,
    -- layer=1 filter=147 channel=23
    -9, 24, -14, -27, -70, -50, -9, -13, -1,
    -- layer=1 filter=147 channel=24
    20, 18, -8, 12, -7, 11, -15, -15, -24,
    -- layer=1 filter=147 channel=25
    -2, 34, 7, 85, 7, -20, -12, 42, 38,
    -- layer=1 filter=147 channel=26
    -17, -3, -5, 7, -22, 12, 11, 10, -10,
    -- layer=1 filter=147 channel=27
    18, 37, 40, 5, 2, 17, 1, -15, -13,
    -- layer=1 filter=147 channel=28
    -15, 28, 5, 33, -2, -40, -17, -2, 1,
    -- layer=1 filter=147 channel=29
    3, -1, 8, -11, -11, -26, -22, -13, -10,
    -- layer=1 filter=147 channel=30
    1, -16, -8, 4, -3, 37, 23, 26, 0,
    -- layer=1 filter=147 channel=31
    -16, -37, 10, -23, -6, 19, -4, 8, 10,
    -- layer=1 filter=147 channel=32
    -11, -27, -18, 11, -4, 11, 35, 16, 6,
    -- layer=1 filter=147 channel=33
    1, 16, 25, 23, 1, 8, -2, -4, -4,
    -- layer=1 filter=147 channel=34
    -8, -9, 6, -7, 0, -5, 4, 9, -10,
    -- layer=1 filter=147 channel=35
    1, 3, -7, 7, -10, -13, 0, -2, -1,
    -- layer=1 filter=147 channel=36
    0, 15, 8, 2, 7, 8, 2, -6, -1,
    -- layer=1 filter=147 channel=37
    16, 30, 0, 60, 8, 3, -34, 30, 8,
    -- layer=1 filter=147 channel=38
    -9, -12, 13, 11, 1, 0, -2, 5, -6,
    -- layer=1 filter=147 channel=39
    22, 13, 10, 0, 1, -5, -13, -13, 1,
    -- layer=1 filter=147 channel=40
    -22, -13, 15, 0, 17, 15, 30, 16, -22,
    -- layer=1 filter=147 channel=41
    12, 21, -32, 46, -4, 25, 66, 57, 13,
    -- layer=1 filter=147 channel=42
    -11, 8, -19, -2, -16, -24, 28, 10, -5,
    -- layer=1 filter=147 channel=43
    -6, 18, -1, 42, 15, -38, -33, 25, 20,
    -- layer=1 filter=147 channel=44
    3, -20, -4, 19, -6, -2, 5, 1, -9,
    -- layer=1 filter=147 channel=45
    4, -19, -10, 6, -19, -9, -35, -7, -20,
    -- layer=1 filter=147 channel=46
    15, 66, 28, 43, 26, 30, 5, 65, -3,
    -- layer=1 filter=147 channel=47
    -4, -10, -20, 3, -37, 9, 40, 19, 13,
    -- layer=1 filter=147 channel=48
    19, 20, 11, -3, -2, -6, -13, -28, -32,
    -- layer=1 filter=147 channel=49
    5, 2, -15, -10, -11, 8, 2, 4, -32,
    -- layer=1 filter=147 channel=50
    3, -3, 20, 3, 1, 4, -5, -1, -15,
    -- layer=1 filter=147 channel=51
    -3, 0, 10, 22, -1, -2, -2, -17, -1,
    -- layer=1 filter=147 channel=52
    8, -16, -7, -5, 7, -8, 3, 13, 15,
    -- layer=1 filter=147 channel=53
    -20, -19, 10, 3, -16, -6, -20, -10, -9,
    -- layer=1 filter=147 channel=54
    29, 53, 3, 84, 29, -11, 8, 71, 40,
    -- layer=1 filter=147 channel=55
    18, 2, 6, -3, -17, -1, 0, -13, 22,
    -- layer=1 filter=147 channel=56
    -3, 1, -8, 8, 1, 1, 10, -6, -10,
    -- layer=1 filter=147 channel=57
    -30, -21, -18, 23, -16, -11, -29, 10, 25,
    -- layer=1 filter=147 channel=58
    18, 12, -3, 24, -32, -18, -1, 34, 52,
    -- layer=1 filter=147 channel=59
    -4, 9, -13, -11, -12, -11, 3, 12, -6,
    -- layer=1 filter=147 channel=60
    18, 4, 18, 10, 4, 3, 10, 19, 14,
    -- layer=1 filter=147 channel=61
    -13, 12, -16, 7, -6, 4, 3, 4, -3,
    -- layer=1 filter=147 channel=62
    10, 22, 14, 63, 0, -30, -36, 18, 0,
    -- layer=1 filter=147 channel=63
    9, 17, 20, 8, 0, 13, 2, -17, -23,
    -- layer=1 filter=147 channel=64
    -8, 1, 7, 5, 1, -5, -10, -10, -6,
    -- layer=1 filter=147 channel=65
    19, 0, 18, 23, -5, -16, -20, -26, -38,
    -- layer=1 filter=147 channel=66
    11, 24, 9, -6, -9, -21, 0, -19, -13,
    -- layer=1 filter=147 channel=67
    16, 16, 10, 3, 1, -6, -7, -10, -17,
    -- layer=1 filter=147 channel=68
    0, -24, 5, 33, -7, 4, 28, 7, -2,
    -- layer=1 filter=147 channel=69
    -4, -32, -33, -4, -49, -12, -50, -14, -10,
    -- layer=1 filter=147 channel=70
    -14, -16, 1, -19, -4, 11, 10, -9, -11,
    -- layer=1 filter=147 channel=71
    24, 32, 33, 25, 0, -25, -23, -31, -6,
    -- layer=1 filter=147 channel=72
    9, 30, -12, 60, 13, 58, 44, 63, 10,
    -- layer=1 filter=147 channel=73
    5, 8, 1, 4, -10, 0, 4, 0, -16,
    -- layer=1 filter=147 channel=74
    8, -13, -1, 20, 6, -6, 31, 17, -9,
    -- layer=1 filter=147 channel=75
    -44, -59, -17, -50, -54, -40, -26, -37, -14,
    -- layer=1 filter=147 channel=76
    3, 0, 9, 0, 11, -10, 14, -16, -20,
    -- layer=1 filter=147 channel=77
    31, 22, 6, 12, 7, -25, -19, -12, -20,
    -- layer=1 filter=147 channel=78
    19, 1, 11, 15, 11, -13, -5, 7, 17,
    -- layer=1 filter=147 channel=79
    0, 19, 0, 43, 8, -22, -41, -3, 11,
    -- layer=1 filter=147 channel=80
    -1, 9, -5, 12, 7, 4, 7, 10, 7,
    -- layer=1 filter=147 channel=81
    21, 20, -1, -2, 2, -32, -47, -17, -28,
    -- layer=1 filter=147 channel=82
    17, 7, 9, 1, 4, -1, -8, -24, -31,
    -- layer=1 filter=147 channel=83
    -2, -48, -22, -10, -32, -25, -42, -9, -16,
    -- layer=1 filter=147 channel=84
    40, 3, 28, 39, 44, 30, 50, 26, -24,
    -- layer=1 filter=147 channel=85
    15, 41, -6, 22, -35, -19, 13, 36, 27,
    -- layer=1 filter=147 channel=86
    4, 19, 6, 6, 2, -9, -2, -7, 3,
    -- layer=1 filter=147 channel=87
    61, 69, -4, 97, 31, 61, 41, 114, 24,
    -- layer=1 filter=147 channel=88
    -1, 21, 6, 10, 2, 4, 0, -12, -20,
    -- layer=1 filter=147 channel=89
    27, 14, 6, -4, 2, -19, 7, -21, -32,
    -- layer=1 filter=147 channel=90
    -19, -51, -10, -5, -51, 1, -6, -20, -14,
    -- layer=1 filter=147 channel=91
    -10, -4, 0, 3, -3, 15, 3, -3, 0,
    -- layer=1 filter=147 channel=92
    -14, -57, -38, -28, -57, -17, -4, -12, 21,
    -- layer=1 filter=147 channel=93
    6, 16, -5, 15, -10, -21, -26, -32, -24,
    -- layer=1 filter=147 channel=94
    -6, 0, -3, -1, 1, 0, -10, -19, -26,
    -- layer=1 filter=147 channel=95
    19, 7, 33, 35, 45, 9, 54, 19, -25,
    -- layer=1 filter=147 channel=96
    10, 21, 13, -1, -6, 7, 4, -9, 9,
    -- layer=1 filter=147 channel=97
    10, 5, 11, 8, -8, -20, -24, -18, -14,
    -- layer=1 filter=147 channel=98
    -15, 7, -23, 29, 6, -41, -36, 0, 25,
    -- layer=1 filter=147 channel=99
    -4, -24, -25, 0, -21, -35, -25, -2, -41,
    -- layer=1 filter=147 channel=100
    6, -7, 8, 7, 6, 13, 4, 0, -10,
    -- layer=1 filter=147 channel=101
    -3, -5, 0, -5, 14, -12, 13, -11, -13,
    -- layer=1 filter=147 channel=102
    3, -16, -5, -6, 2, -22, 10, -28, -34,
    -- layer=1 filter=147 channel=103
    3, 16, 8, 1, 7, 29, -9, -3, -4,
    -- layer=1 filter=147 channel=104
    -20, 21, -6, 10, -25, -7, 27, 22, 7,
    -- layer=1 filter=147 channel=105
    2, -2, 14, -5, -4, -18, -20, -26, -13,
    -- layer=1 filter=147 channel=106
    -9, -20, -7, 12, 21, 0, 18, 3, -26,
    -- layer=1 filter=147 channel=107
    0, 1, -1, -2, -6, -15, 11, 12, 11,
    -- layer=1 filter=147 channel=108
    -12, -44, -15, 3, -36, -28, 3, 9, -8,
    -- layer=1 filter=147 channel=109
    -6, -4, -4, -12, 6, -6, -3, -10, -2,
    -- layer=1 filter=147 channel=110
    10, 0, 0, 0, 0, 6, -11, 4, 1,
    -- layer=1 filter=147 channel=111
    11, -25, 12, -15, -4, 24, 18, -13, -47,
    -- layer=1 filter=147 channel=112
    35, -7, 8, -5, 21, 3, 36, -22, -22,
    -- layer=1 filter=147 channel=113
    14, 23, 20, 0, -11, 6, 5, -4, -22,
    -- layer=1 filter=147 channel=114
    -15, -17, -8, 15, -17, -25, -41, -35, -29,
    -- layer=1 filter=147 channel=115
    -15, 2, 13, -3, -8, -17, -19, -12, 2,
    -- layer=1 filter=147 channel=116
    -12, 1, -4, 0, 3, 1, 1, -1, 0,
    -- layer=1 filter=147 channel=117
    8, -46, -24, 10, 21, -1, 3, -34, -13,
    -- layer=1 filter=147 channel=118
    9, 0, 15, 2, 19, 15, 40, 16, -23,
    -- layer=1 filter=147 channel=119
    -8, -7, -5, 27, -10, 9, 38, 5, 9,
    -- layer=1 filter=147 channel=120
    -1, 15, -6, 12, -11, -7, -33, 0, 11,
    -- layer=1 filter=147 channel=121
    -5, 8, -2, 3, -2, 8, -21, 10, 0,
    -- layer=1 filter=147 channel=122
    -1, -9, -5, -4, -2, 5, 9, -1, -6,
    -- layer=1 filter=147 channel=123
    -16, 2, -1, -7, -3, 8, -10, 7, 0,
    -- layer=1 filter=147 channel=124
    -3, 0, -10, 0, -11, -2, -5, 3, -1,
    -- layer=1 filter=147 channel=125
    -17, -38, -4, -17, -7, -6, -20, 7, 6,
    -- layer=1 filter=147 channel=126
    14, -12, -48, 17, -3, -26, -34, 21, 28,
    -- layer=1 filter=147 channel=127
    10, -11, 26, 13, 29, 14, 31, 20, -22,
    -- layer=1 filter=148 channel=0
    -10, -7, -13, 2, 3, 1, -5, -7, -5,
    -- layer=1 filter=148 channel=1
    -10, 8, -4, 8, -8, 0, 0, -10, -10,
    -- layer=1 filter=148 channel=2
    -7, -14, -6, 8, 13, -1, 9, 6, 19,
    -- layer=1 filter=148 channel=3
    -10, 7, 2, -8, 4, 0, -8, 8, -2,
    -- layer=1 filter=148 channel=4
    5, -11, 3, -3, 1, -4, 6, 3, -3,
    -- layer=1 filter=148 channel=5
    -4, 0, -4, -18, -16, -24, -18, -10, 4,
    -- layer=1 filter=148 channel=6
    -2, -1, -1, -16, -22, -2, 0, -5, -5,
    -- layer=1 filter=148 channel=7
    7, -9, -9, -8, -7, -6, -20, -5, -6,
    -- layer=1 filter=148 channel=8
    -5, 4, 1, -10, -5, -14, -20, -13, -13,
    -- layer=1 filter=148 channel=9
    -1, 1, -4, 1, 7, -1, -8, -5, 4,
    -- layer=1 filter=148 channel=10
    2, -14, -7, -4, -6, -2, -2, -16, 0,
    -- layer=1 filter=148 channel=11
    -1, -13, -5, -9, -16, -13, -16, -23, -8,
    -- layer=1 filter=148 channel=12
    13, 6, 9, 7, -4, 30, 6, 14, 2,
    -- layer=1 filter=148 channel=13
    -16, -7, -19, -16, -5, 0, -4, -14, -9,
    -- layer=1 filter=148 channel=14
    3, 2, -10, 8, 0, 9, -3, 1, -15,
    -- layer=1 filter=148 channel=15
    -12, -11, -2, -3, 0, -4, -10, -4, -10,
    -- layer=1 filter=148 channel=16
    1, -3, -7, -5, -16, -17, 0, -7, -11,
    -- layer=1 filter=148 channel=17
    -3, -13, -7, -8, -10, -3, 6, 0, 4,
    -- layer=1 filter=148 channel=18
    6, 1, 6, -18, -3, 9, -3, -12, -17,
    -- layer=1 filter=148 channel=19
    4, -8, -2, -13, -13, -17, -11, -16, -11,
    -- layer=1 filter=148 channel=20
    -3, -17, -17, -10, -17, -18, -21, -2, -2,
    -- layer=1 filter=148 channel=21
    -9, -9, -3, -3, -16, -2, -7, -3, -17,
    -- layer=1 filter=148 channel=22
    0, -8, -23, -3, -19, -8, -24, -21, -5,
    -- layer=1 filter=148 channel=23
    -9, -15, -10, -8, -15, -13, -10, -9, 2,
    -- layer=1 filter=148 channel=24
    -12, -7, -19, -6, -11, -13, 3, -15, -7,
    -- layer=1 filter=148 channel=25
    -5, -24, -17, -23, -18, -7, -12, -7, -16,
    -- layer=1 filter=148 channel=26
    -8, -19, -26, -15, -14, -10, 5, -12, -11,
    -- layer=1 filter=148 channel=27
    10, -8, 0, -25, -19, -20, -23, -19, -12,
    -- layer=1 filter=148 channel=28
    2, -11, 0, -2, -3, -19, -20, -26, -10,
    -- layer=1 filter=148 channel=29
    5, -8, -1, -4, -17, 4, -11, -5, -12,
    -- layer=1 filter=148 channel=30
    11, -1, 9, -24, -11, -3, -11, -22, -6,
    -- layer=1 filter=148 channel=31
    12, 20, 16, -12, -1, -9, -14, -6, -6,
    -- layer=1 filter=148 channel=32
    1, -10, -18, 6, 7, 0, -7, -8, -22,
    -- layer=1 filter=148 channel=33
    -3, -1, -14, -10, -5, -10, -5, -6, -3,
    -- layer=1 filter=148 channel=34
    5, -9, -12, -2, 0, 6, -3, 3, 0,
    -- layer=1 filter=148 channel=35
    7, -2, -3, -7, 5, 1, 7, -10, 7,
    -- layer=1 filter=148 channel=36
    -9, -15, -1, -24, -8, -18, -2, -9, -16,
    -- layer=1 filter=148 channel=37
    3, -14, -3, -9, -19, -4, -13, -4, 5,
    -- layer=1 filter=148 channel=38
    1, 0, -10, -8, -9, -8, -15, -22, -20,
    -- layer=1 filter=148 channel=39
    0, 8, 6, 3, -1, -9, -9, 0, -11,
    -- layer=1 filter=148 channel=40
    4, -5, 14, 0, -1, -2, -16, -10, -11,
    -- layer=1 filter=148 channel=41
    -13, -17, -17, -1, -2, -13, -9, -4, -18,
    -- layer=1 filter=148 channel=42
    16, -14, -4, 20, 8, 11, 9, 14, 6,
    -- layer=1 filter=148 channel=43
    -1, -14, -4, -17, -16, -12, -15, -6, -12,
    -- layer=1 filter=148 channel=44
    0, -1, -12, 4, -20, -16, -1, -15, -14,
    -- layer=1 filter=148 channel=45
    -3, -13, -6, 0, -6, -4, 0, -1, 2,
    -- layer=1 filter=148 channel=46
    29, 16, 9, 10, 17, 29, 3, 12, -1,
    -- layer=1 filter=148 channel=47
    -13, -5, 1, -6, 3, -6, 1, 2, 5,
    -- layer=1 filter=148 channel=48
    -6, 5, 0, 0, -5, 2, -14, -1, -10,
    -- layer=1 filter=148 channel=49
    -3, -4, -7, -2, -13, -12, -16, -9, 0,
    -- layer=1 filter=148 channel=50
    -6, 0, 8, 2, 0, -11, -9, -7, 3,
    -- layer=1 filter=148 channel=51
    2, -2, 3, -16, -12, 3, -2, -9, -11,
    -- layer=1 filter=148 channel=52
    -2, 0, -3, -9, -6, 2, 2, 6, 10,
    -- layer=1 filter=148 channel=53
    -10, 9, 7, 6, 8, -12, 1, 3, -3,
    -- layer=1 filter=148 channel=54
    -6, -11, 0, 2, -3, -4, 0, -4, -6,
    -- layer=1 filter=148 channel=55
    -12, -12, -16, -4, -10, -4, -9, 2, -14,
    -- layer=1 filter=148 channel=56
    -7, -8, -10, -2, -10, -5, 1, -6, -10,
    -- layer=1 filter=148 channel=57
    -11, -18, -9, -24, -14, -1, -8, -18, -3,
    -- layer=1 filter=148 channel=58
    -15, -1, -14, 7, 16, 7, -1, -2, -6,
    -- layer=1 filter=148 channel=59
    8, 7, 0, 8, -10, 4, 1, -10, -10,
    -- layer=1 filter=148 channel=60
    0, 5, 0, -1, -3, 6, 4, -2, 5,
    -- layer=1 filter=148 channel=61
    10, 0, -5, -9, -10, -4, 10, -7, -4,
    -- layer=1 filter=148 channel=62
    -9, -7, -17, -9, -19, -4, -13, -6, -8,
    -- layer=1 filter=148 channel=63
    -2, -12, -13, -5, -19, -13, -5, -14, -23,
    -- layer=1 filter=148 channel=64
    -3, 0, -5, -2, -8, -2, -12, -4, 0,
    -- layer=1 filter=148 channel=65
    3, -15, -10, -7, 3, 0, 0, -2, -13,
    -- layer=1 filter=148 channel=66
    -21, -9, -12, 0, -18, -14, -16, -14, -15,
    -- layer=1 filter=148 channel=67
    -2, 0, -8, 1, -5, -11, 6, 12, 12,
    -- layer=1 filter=148 channel=68
    0, -13, -25, -5, -8, -18, -3, -11, -16,
    -- layer=1 filter=148 channel=69
    -6, -16, -7, 4, -14, -4, 2, -4, -3,
    -- layer=1 filter=148 channel=70
    9, 27, 34, -15, -8, -8, -17, -7, 0,
    -- layer=1 filter=148 channel=71
    3, -1, 3, -15, -13, 0, -7, -23, -1,
    -- layer=1 filter=148 channel=72
    3, 8, -17, -13, 6, 7, -14, -10, 0,
    -- layer=1 filter=148 channel=73
    -3, -3, 4, -10, -2, -2, -1, -8, -9,
    -- layer=1 filter=148 channel=74
    1, -12, -10, -9, -16, -3, -6, -7, -15,
    -- layer=1 filter=148 channel=75
    6, 17, -4, 10, 1, 19, 0, 5, -1,
    -- layer=1 filter=148 channel=76
    -7, 0, -5, -7, -5, -7, -6, -1, -10,
    -- layer=1 filter=148 channel=77
    0, 0, 4, -5, -2, 4, -11, 0, -4,
    -- layer=1 filter=148 channel=78
    8, -6, 3, 7, -11, 5, -6, -4, -9,
    -- layer=1 filter=148 channel=79
    -8, -5, -22, -7, -4, -14, -12, -2, 0,
    -- layer=1 filter=148 channel=80
    -8, -9, -7, -1, 10, 1, 1, 4, -7,
    -- layer=1 filter=148 channel=81
    -11, -6, -4, -8, -15, -10, -12, -3, -8,
    -- layer=1 filter=148 channel=82
    -14, 2, -5, -14, -2, -13, -3, 0, -8,
    -- layer=1 filter=148 channel=83
    -6, -7, 2, 7, -15, -6, -6, -1, -11,
    -- layer=1 filter=148 channel=84
    -3, -11, 6, 1, -6, -1, -11, -10, -10,
    -- layer=1 filter=148 channel=85
    -6, -13, -4, -8, 7, 3, 1, 0, 5,
    -- layer=1 filter=148 channel=86
    7, 1, 1, -10, -3, -11, -8, -9, 0,
    -- layer=1 filter=148 channel=87
    0, -5, 7, -9, 0, -9, -7, -15, 0,
    -- layer=1 filter=148 channel=88
    -9, -7, -6, -3, 0, -3, -3, -3, -10,
    -- layer=1 filter=148 channel=89
    -15, 4, -16, 5, -3, 0, -12, -11, -21,
    -- layer=1 filter=148 channel=90
    2, 2, -8, 9, -8, -6, -2, -4, -15,
    -- layer=1 filter=148 channel=91
    -2, -9, 2, -2, -16, -8, -15, -7, -14,
    -- layer=1 filter=148 channel=92
    -13, -5, -16, 3, -6, -9, -4, -10, -5,
    -- layer=1 filter=148 channel=93
    -17, -13, -16, -22, -13, -20, -24, -23, -16,
    -- layer=1 filter=148 channel=94
    -5, -14, -17, 3, -15, 0, -4, -15, -8,
    -- layer=1 filter=148 channel=95
    -10, 0, -11, 0, -16, -6, -16, -14, 1,
    -- layer=1 filter=148 channel=96
    -1, -3, 9, 0, -12, 0, -5, -7, 5,
    -- layer=1 filter=148 channel=97
    -4, -15, -6, -11, -21, -27, -5, -7, -4,
    -- layer=1 filter=148 channel=98
    -9, -1, -29, -18, -20, -8, -4, -1, 0,
    -- layer=1 filter=148 channel=99
    -9, -6, 0, 6, -14, 0, -3, -1, -17,
    -- layer=1 filter=148 channel=100
    -12, -15, -10, -16, -7, -9, -10, 2, -11,
    -- layer=1 filter=148 channel=101
    0, -8, -11, 1, -12, -7, -6, -5, -24,
    -- layer=1 filter=148 channel=102
    -18, -16, -17, -7, -15, -14, -1, 0, -3,
    -- layer=1 filter=148 channel=103
    -16, -6, -1, -26, -26, -18, 0, -9, -9,
    -- layer=1 filter=148 channel=104
    9, 4, 7, -7, -4, -4, -7, 4, 10,
    -- layer=1 filter=148 channel=105
    -5, -5, -12, -8, -7, -15, -8, -12, -17,
    -- layer=1 filter=148 channel=106
    -8, -6, -17, -3, -10, -12, -1, -24, -27,
    -- layer=1 filter=148 channel=107
    -2, -7, 4, -9, -7, 3, -11, -5, 1,
    -- layer=1 filter=148 channel=108
    -3, -5, -8, 7, -8, -22, 4, -8, -9,
    -- layer=1 filter=148 channel=109
    -11, 0, -1, -3, 9, -3, -2, -3, 3,
    -- layer=1 filter=148 channel=110
    -4, 2, 2, -6, -10, -11, -9, -6, 2,
    -- layer=1 filter=148 channel=111
    -8, 6, 3, -18, -9, -6, -23, -13, -9,
    -- layer=1 filter=148 channel=112
    -11, 3, 4, -3, -10, 7, 3, 5, -1,
    -- layer=1 filter=148 channel=113
    6, 3, -7, 7, -5, -5, -12, -7, -7,
    -- layer=1 filter=148 channel=114
    13, -18, 8, -9, -13, -14, -10, -2, -2,
    -- layer=1 filter=148 channel=115
    -3, -14, -11, -4, -4, -10, -3, -9, -22,
    -- layer=1 filter=148 channel=116
    -6, -6, 9, -7, -5, 10, 11, -3, 1,
    -- layer=1 filter=148 channel=117
    -8, 12, 11, -9, 2, -9, -9, 4, -6,
    -- layer=1 filter=148 channel=118
    2, 5, -3, -19, -13, 0, -1, -22, -10,
    -- layer=1 filter=148 channel=119
    -6, -9, -14, -1, -4, -4, -4, -7, -15,
    -- layer=1 filter=148 channel=120
    0, -16, -18, -11, -5, -18, -18, -11, -16,
    -- layer=1 filter=148 channel=121
    9, 0, 2, 2, -2, -7, 3, -5, 0,
    -- layer=1 filter=148 channel=122
    10, -4, -9, 0, -1, -7, -10, -4, 9,
    -- layer=1 filter=148 channel=123
    -10, 6, -10, -6, -13, 4, -7, -12, -4,
    -- layer=1 filter=148 channel=124
    -5, -4, 7, -9, -8, -10, 1, 3, 0,
    -- layer=1 filter=148 channel=125
    -3, 0, 12, 0, -8, -11, -3, -15, -11,
    -- layer=1 filter=148 channel=126
    6, -4, -5, -7, -9, 0, -16, -1, 2,
    -- layer=1 filter=148 channel=127
    0, -3, -5, -13, -5, 0, -17, -18, 3,
    -- layer=1 filter=149 channel=0
    8, 8, -8, 2, 0, 1, -7, 2, -9,
    -- layer=1 filter=149 channel=1
    -1, -9, -3, -11, -16, -5, -14, -8, -9,
    -- layer=1 filter=149 channel=2
    -11, -3, -2, 4, -4, -7, 25, 7, -17,
    -- layer=1 filter=149 channel=3
    5, -9, -6, -10, 2, 3, -8, -6, 3,
    -- layer=1 filter=149 channel=4
    0, 7, 1, 2, 0, -11, 3, -7, 1,
    -- layer=1 filter=149 channel=5
    -7, -25, -32, -13, -18, -6, -3, -18, -22,
    -- layer=1 filter=149 channel=6
    -2, 0, 6, -3, -10, -6, -7, -5, 1,
    -- layer=1 filter=149 channel=7
    -18, -22, -19, -3, -17, -10, -26, 5, 0,
    -- layer=1 filter=149 channel=8
    -1, -3, -21, 0, -1, -3, -19, -9, -12,
    -- layer=1 filter=149 channel=9
    0, 2, -7, 11, 7, -3, 9, 4, -18,
    -- layer=1 filter=149 channel=10
    -19, -25, -2, -13, -8, 9, -20, -7, 9,
    -- layer=1 filter=149 channel=11
    -4, 10, -6, -4, -9, -8, 8, -17, 2,
    -- layer=1 filter=149 channel=12
    22, 3, -2, 10, 1, -3, -5, 6, 8,
    -- layer=1 filter=149 channel=13
    -2, -5, -10, -3, -5, -12, -6, -7, -14,
    -- layer=1 filter=149 channel=14
    1, -10, -10, -6, -3, -2, -25, 19, 0,
    -- layer=1 filter=149 channel=15
    -3, -8, -20, 0, 1, -15, 2, -2, -3,
    -- layer=1 filter=149 channel=16
    -12, -14, -16, -7, -9, 3, 0, -12, -29,
    -- layer=1 filter=149 channel=17
    -4, -2, -20, 0, -12, -22, 0, -22, -22,
    -- layer=1 filter=149 channel=18
    4, 6, -18, -1, -14, 1, -7, 4, -4,
    -- layer=1 filter=149 channel=19
    -8, 4, -5, -2, -10, -5, -2, 9, 4,
    -- layer=1 filter=149 channel=20
    -20, -22, 0, -18, -14, -5, -22, -19, -15,
    -- layer=1 filter=149 channel=21
    -3, -8, -3, 0, 0, -4, -12, -4, -5,
    -- layer=1 filter=149 channel=22
    -1, -9, -14, -18, -5, -15, -17, -13, -14,
    -- layer=1 filter=149 channel=23
    6, 0, 1, -9, 8, 1, -22, -10, -10,
    -- layer=1 filter=149 channel=24
    -12, -3, -11, -12, -14, -1, 0, 0, -19,
    -- layer=1 filter=149 channel=25
    -15, -3, -6, -11, -10, -3, -22, -21, -4,
    -- layer=1 filter=149 channel=26
    2, 5, -9, -6, -5, -3, 16, -17, -6,
    -- layer=1 filter=149 channel=27
    -3, -5, -16, 3, -20, -15, 12, -5, -7,
    -- layer=1 filter=149 channel=28
    -21, -8, -5, -21, -1, 1, -13, -19, -13,
    -- layer=1 filter=149 channel=29
    0, -7, -2, -5, -3, -11, -1, -18, -1,
    -- layer=1 filter=149 channel=30
    7, -5, -2, -10, -16, -12, -14, 4, -9,
    -- layer=1 filter=149 channel=31
    -8, -10, -19, 5, -12, 0, -10, -8, -18,
    -- layer=1 filter=149 channel=32
    5, 10, 4, -5, -1, -12, -3, -2, 1,
    -- layer=1 filter=149 channel=33
    2, -3, 6, -1, 1, 3, -1, -10, 14,
    -- layer=1 filter=149 channel=34
    -2, -5, 8, -8, 3, -1, 7, 7, -3,
    -- layer=1 filter=149 channel=35
    -3, -10, 1, -7, -7, 8, 0, -9, -1,
    -- layer=1 filter=149 channel=36
    3, -4, -14, 0, -16, 0, 9, -13, -7,
    -- layer=1 filter=149 channel=37
    -14, -11, -30, -26, -4, 5, -16, -23, -27,
    -- layer=1 filter=149 channel=38
    -1, -19, -10, -7, -18, -19, -15, -11, -19,
    -- layer=1 filter=149 channel=39
    -12, -4, -1, 3, -6, -4, -4, 0, 0,
    -- layer=1 filter=149 channel=40
    -6, -8, -8, 5, -12, -28, -7, -11, -5,
    -- layer=1 filter=149 channel=41
    0, 4, 1, -8, 0, -9, 3, -7, -10,
    -- layer=1 filter=149 channel=42
    -11, -20, -8, 6, -6, 0, -5, 4, -18,
    -- layer=1 filter=149 channel=43
    8, -16, -13, -9, -4, 1, -6, -13, -17,
    -- layer=1 filter=149 channel=44
    -2, -9, -4, -5, -6, -20, 11, -10, -8,
    -- layer=1 filter=149 channel=45
    -3, -13, -16, 6, -9, -10, -15, -13, -6,
    -- layer=1 filter=149 channel=46
    0, 12, -1, 4, 1, 5, -10, 14, -20,
    -- layer=1 filter=149 channel=47
    -19, 0, -1, -12, 4, 12, 3, -6, 0,
    -- layer=1 filter=149 channel=48
    -6, -14, -13, -9, -12, -10, -5, 0, -14,
    -- layer=1 filter=149 channel=49
    -14, -13, -8, -16, -3, -9, 0, -15, -6,
    -- layer=1 filter=149 channel=50
    -11, -2, -8, 2, 3, -10, 6, -8, -6,
    -- layer=1 filter=149 channel=51
    -19, -16, -4, -25, -1, -19, -13, -15, -17,
    -- layer=1 filter=149 channel=52
    1, 5, 0, 10, -4, 5, 1, -10, 4,
    -- layer=1 filter=149 channel=53
    -11, 2, -7, 6, -11, 3, -8, -8, -6,
    -- layer=1 filter=149 channel=54
    -21, -2, -9, -9, 5, 5, -17, 2, -4,
    -- layer=1 filter=149 channel=55
    -12, -1, -3, -16, -4, -14, -10, -16, -9,
    -- layer=1 filter=149 channel=56
    6, 0, 0, -9, -4, 6, 2, -4, -6,
    -- layer=1 filter=149 channel=57
    -15, -20, -20, -11, -20, -8, -21, -17, 6,
    -- layer=1 filter=149 channel=58
    -8, 9, -1, -13, 11, -9, -3, 4, 0,
    -- layer=1 filter=149 channel=59
    3, -9, 6, -7, -11, -9, 5, -7, 7,
    -- layer=1 filter=149 channel=60
    0, -8, -7, -2, 7, -9, 1, 8, 9,
    -- layer=1 filter=149 channel=61
    6, 9, -2, 12, 0, -12, -9, 1, -1,
    -- layer=1 filter=149 channel=62
    -6, -21, -15, -19, -14, -10, -4, -12, -10,
    -- layer=1 filter=149 channel=63
    8, 4, -1, 0, 5, -9, -2, -5, -6,
    -- layer=1 filter=149 channel=64
    7, 5, 5, 5, 5, 6, -6, 4, 6,
    -- layer=1 filter=149 channel=65
    -6, -6, 4, 0, 5, 4, -12, -4, 1,
    -- layer=1 filter=149 channel=66
    -4, -9, -12, -14, -1, -5, -7, -7, -7,
    -- layer=1 filter=149 channel=67
    -6, -20, -10, -11, 7, -2, -22, -7, -4,
    -- layer=1 filter=149 channel=68
    8, -2, -12, 18, 7, -6, 18, -1, -11,
    -- layer=1 filter=149 channel=69
    12, -12, -25, -13, -20, -4, -16, -17, -11,
    -- layer=1 filter=149 channel=70
    -24, -6, -8, -2, 0, 3, -13, -3, 0,
    -- layer=1 filter=149 channel=71
    -10, -13, -10, -16, -8, -8, -6, 0, 1,
    -- layer=1 filter=149 channel=72
    7, 1, -8, 7, -3, -3, -10, -5, 3,
    -- layer=1 filter=149 channel=73
    -1, 0, 8, 0, -2, -12, 4, 6, 6,
    -- layer=1 filter=149 channel=74
    4, 2, -20, -4, 4, -5, 1, -4, -4,
    -- layer=1 filter=149 channel=75
    8, 6, -2, 7, -16, -13, 5, 7, 1,
    -- layer=1 filter=149 channel=76
    1, 2, 2, 0, -11, 2, 0, 0, 3,
    -- layer=1 filter=149 channel=77
    -12, -3, -9, 9, 2, -7, -7, 1, 0,
    -- layer=1 filter=149 channel=78
    4, -12, -1, -8, -10, -9, -8, 2, -12,
    -- layer=1 filter=149 channel=79
    0, -3, -10, -21, -16, -8, -14, -23, -14,
    -- layer=1 filter=149 channel=80
    1, 8, -7, 2, 8, -8, -9, 10, -3,
    -- layer=1 filter=149 channel=81
    -2, 1, -2, -16, -6, -5, -10, -9, -15,
    -- layer=1 filter=149 channel=82
    -7, -3, -17, -15, -17, -12, -16, -5, -11,
    -- layer=1 filter=149 channel=83
    0, -9, -12, -5, -12, -13, 3, -17, -20,
    -- layer=1 filter=149 channel=84
    -10, -1, -5, -2, 9, -8, 4, -13, -7,
    -- layer=1 filter=149 channel=85
    -16, 8, -5, -20, 4, -11, -11, 10, -18,
    -- layer=1 filter=149 channel=86
    -13, -9, -4, 0, -17, -18, -20, -9, -23,
    -- layer=1 filter=149 channel=87
    4, 1, 6, 7, -7, -9, 2, 13, -2,
    -- layer=1 filter=149 channel=88
    -5, -3, 1, -16, 0, -5, -19, -12, -4,
    -- layer=1 filter=149 channel=89
    -8, -3, -17, -2, -1, -17, -6, -11, -15,
    -- layer=1 filter=149 channel=90
    7, -3, -1, -1, -8, -15, -2, -17, -19,
    -- layer=1 filter=149 channel=91
    -21, -13, -15, -17, -23, -13, -11, -17, -21,
    -- layer=1 filter=149 channel=92
    0, -7, -8, 1, -10, -12, 1, -19, -6,
    -- layer=1 filter=149 channel=93
    -19, -7, -1, -6, -3, -4, -11, -14, -9,
    -- layer=1 filter=149 channel=94
    -4, -10, -5, -2, 4, 3, -13, -3, -9,
    -- layer=1 filter=149 channel=95
    1, 5, -1, 4, 3, -4, 18, -7, 3,
    -- layer=1 filter=149 channel=96
    0, -7, -7, 4, -7, -6, 8, -10, -9,
    -- layer=1 filter=149 channel=97
    0, 0, 0, -3, 3, -2, -19, -14, -8,
    -- layer=1 filter=149 channel=98
    2, -18, -26, -2, -5, 4, -6, -12, -8,
    -- layer=1 filter=149 channel=99
    -21, -9, -5, -12, -2, -7, -2, 0, -3,
    -- layer=1 filter=149 channel=100
    9, 3, -8, 5, 5, 8, -5, -3, -11,
    -- layer=1 filter=149 channel=101
    -6, -15, -18, -15, -7, -13, -23, -6, -8,
    -- layer=1 filter=149 channel=102
    -7, -15, -3, 0, -8, -11, 0, -8, -10,
    -- layer=1 filter=149 channel=103
    7, 7, 1, -8, -4, 5, 4, -7, 5,
    -- layer=1 filter=149 channel=104
    -1, -9, -7, -4, 4, 6, 6, 7, -11,
    -- layer=1 filter=149 channel=105
    -14, -15, -16, -10, -7, -16, -1, -16, -11,
    -- layer=1 filter=149 channel=106
    0, -6, -8, -8, -17, -10, -17, -15, -1,
    -- layer=1 filter=149 channel=107
    3, -3, 7, -5, -9, -8, -9, 1, -5,
    -- layer=1 filter=149 channel=108
    1, -1, -15, -9, 8, -8, -4, -9, -22,
    -- layer=1 filter=149 channel=109
    -1, 6, 10, -3, 3, 0, -9, 3, -3,
    -- layer=1 filter=149 channel=110
    7, 1, -6, -11, -2, -7, 3, 3, 7,
    -- layer=1 filter=149 channel=111
    5, 6, -9, 6, -9, -12, 9, -2, -1,
    -- layer=1 filter=149 channel=112
    -12, -5, -10, 0, 3, 5, 7, 1, -8,
    -- layer=1 filter=149 channel=113
    -18, -21, 2, -17, -17, -9, -14, -5, -19,
    -- layer=1 filter=149 channel=114
    5, -14, -20, -9, -11, -14, -18, -10, -15,
    -- layer=1 filter=149 channel=115
    -5, -7, -14, -9, -11, -17, -13, -5, -21,
    -- layer=1 filter=149 channel=116
    -8, 7, -2, 10, -2, -9, 10, -8, -6,
    -- layer=1 filter=149 channel=117
    -5, 0, -4, -1, -1, 0, -3, -5, 3,
    -- layer=1 filter=149 channel=118
    0, -12, -4, 9, -7, 0, 0, -21, -6,
    -- layer=1 filter=149 channel=119
    2, -5, -1, -7, -2, 0, 3, -15, -11,
    -- layer=1 filter=149 channel=120
    -18, -13, -4, -17, -4, -14, -16, -14, -18,
    -- layer=1 filter=149 channel=121
    5, -1, 6, 5, -3, 0, 0, 2, -13,
    -- layer=1 filter=149 channel=122
    -5, 9, -7, 4, -3, -4, -3, 1, -3,
    -- layer=1 filter=149 channel=123
    -7, -3, -9, -14, -3, -13, 2, 13, -2,
    -- layer=1 filter=149 channel=124
    -11, -3, -8, 8, 0, -5, -2, 0, 0,
    -- layer=1 filter=149 channel=125
    -1, -6, -11, -10, -9, -2, -8, -18, -7,
    -- layer=1 filter=149 channel=126
    7, -11, -19, -4, -3, -13, -12, -13, -1,
    -- layer=1 filter=149 channel=127
    -7, -1, -8, -4, -20, -22, -2, -6, -17,
    -- layer=1 filter=150 channel=0
    -12, -1, -8, -10, -4, -11, -1, -2, -1,
    -- layer=1 filter=150 channel=1
    -3, -3, -7, -8, -8, 2, -11, -9, -3,
    -- layer=1 filter=150 channel=2
    -9, 4, 5, -8, 5, 2, 2, -9, 9,
    -- layer=1 filter=150 channel=3
    5, -2, 1, 8, 0, -9, 3, 7, 9,
    -- layer=1 filter=150 channel=4
    4, 0, -10, -7, -11, 0, 3, -12, 0,
    -- layer=1 filter=150 channel=5
    2, 2, -10, -4, -11, 6, -7, 10, 4,
    -- layer=1 filter=150 channel=6
    4, 5, -2, 1, -8, 2, 6, -5, 5,
    -- layer=1 filter=150 channel=7
    -10, 4, -4, 4, 7, -3, 0, 3, 7,
    -- layer=1 filter=150 channel=8
    3, -6, -5, 6, 1, 6, -11, -12, -10,
    -- layer=1 filter=150 channel=9
    -4, 2, 0, -10, -12, -11, -7, -3, 4,
    -- layer=1 filter=150 channel=10
    -7, -8, -4, 2, 7, -8, -7, -1, -2,
    -- layer=1 filter=150 channel=11
    4, -7, -6, -8, -2, 8, 0, 3, 5,
    -- layer=1 filter=150 channel=12
    -3, -10, 5, 5, -2, -1, 3, 6, 6,
    -- layer=1 filter=150 channel=13
    -1, 2, -1, 0, 8, 8, -3, -4, -2,
    -- layer=1 filter=150 channel=14
    -11, 1, -7, -1, 0, -3, -1, 8, -6,
    -- layer=1 filter=150 channel=15
    -8, 2, -8, 1, 0, -9, 9, 1, 5,
    -- layer=1 filter=150 channel=16
    -9, -11, -5, -12, -11, -2, -9, -8, 1,
    -- layer=1 filter=150 channel=17
    -8, -7, 3, -9, 6, 6, -9, -6, 4,
    -- layer=1 filter=150 channel=18
    -11, 0, -12, -13, 5, 0, -1, 4, 5,
    -- layer=1 filter=150 channel=19
    -12, -1, 0, 7, -5, -2, -8, 2, 2,
    -- layer=1 filter=150 channel=20
    -10, -3, -5, 2, -11, 5, 2, 2, 9,
    -- layer=1 filter=150 channel=21
    -5, -10, 2, -9, 6, 8, 4, 4, 4,
    -- layer=1 filter=150 channel=22
    -9, 6, -12, -8, 4, 1, -7, 4, -9,
    -- layer=1 filter=150 channel=23
    1, -1, -5, 0, 3, -1, 5, 0, -4,
    -- layer=1 filter=150 channel=24
    7, 1, -5, -10, -9, 3, 1, -5, -10,
    -- layer=1 filter=150 channel=25
    7, -9, 3, -3, 5, -11, 6, 0, -5,
    -- layer=1 filter=150 channel=26
    -5, -8, 7, 0, -10, -2, -10, 1, -4,
    -- layer=1 filter=150 channel=27
    -2, 3, 0, 10, 8, 7, 10, 1, 8,
    -- layer=1 filter=150 channel=28
    -2, -9, 2, -1, 2, 7, 6, 4, 2,
    -- layer=1 filter=150 channel=29
    -7, 7, 0, 1, 6, 4, 0, -3, 0,
    -- layer=1 filter=150 channel=30
    -5, 9, 0, 7, 2, -10, -10, 5, -2,
    -- layer=1 filter=150 channel=31
    7, 4, 6, -5, -3, -7, -4, 4, -7,
    -- layer=1 filter=150 channel=32
    8, 1, 2, -8, 3, -12, -8, 5, -5,
    -- layer=1 filter=150 channel=33
    4, -9, -3, -9, 0, 8, 7, -8, 9,
    -- layer=1 filter=150 channel=34
    -6, 6, 5, -6, 1, -1, -8, -9, -5,
    -- layer=1 filter=150 channel=35
    -5, 0, 7, -12, 2, 0, -3, -5, 6,
    -- layer=1 filter=150 channel=36
    -1, -2, 3, -8, 3, 0, 0, -1, 7,
    -- layer=1 filter=150 channel=37
    -5, 0, 10, -7, -4, 7, 1, 7, 1,
    -- layer=1 filter=150 channel=38
    -7, 6, 7, -2, -9, 6, -9, 0, -2,
    -- layer=1 filter=150 channel=39
    -5, 4, 3, -2, -1, -8, 7, -9, 0,
    -- layer=1 filter=150 channel=40
    -7, 2, 1, -2, 0, -2, -9, -2, -11,
    -- layer=1 filter=150 channel=41
    3, 5, -8, -9, -1, -2, -7, 0, 5,
    -- layer=1 filter=150 channel=42
    7, 0, 1, -7, -4, 10, 8, 10, -5,
    -- layer=1 filter=150 channel=43
    2, 6, 5, -6, 6, 3, -8, -8, 3,
    -- layer=1 filter=150 channel=44
    3, 2, 6, -6, 7, -5, 3, -4, 7,
    -- layer=1 filter=150 channel=45
    0, -5, -7, -6, 4, -5, 10, -4, -3,
    -- layer=1 filter=150 channel=46
    -6, -10, 11, -2, -6, -7, -10, 3, -2,
    -- layer=1 filter=150 channel=47
    7, -2, 6, 1, -10, 1, -11, -9, -6,
    -- layer=1 filter=150 channel=48
    4, -5, 5, -3, -6, 7, 7, -5, 6,
    -- layer=1 filter=150 channel=49
    1, -6, 6, 8, 9, -3, 4, 4, 5,
    -- layer=1 filter=150 channel=50
    -6, 2, -1, -5, 3, -2, -9, 8, -1,
    -- layer=1 filter=150 channel=51
    9, 3, 0, -10, -3, 6, 2, 0, -2,
    -- layer=1 filter=150 channel=52
    -11, -1, 10, 6, 7, 0, 4, -4, 12,
    -- layer=1 filter=150 channel=53
    -6, 0, -1, 8, 5, -6, -12, 1, -1,
    -- layer=1 filter=150 channel=54
    0, 0, -7, -4, 1, -10, 5, -7, -4,
    -- layer=1 filter=150 channel=55
    -3, 5, 5, 5, 0, -7, -4, -7, 3,
    -- layer=1 filter=150 channel=56
    -5, 7, -5, 5, 0, 4, -5, -12, -2,
    -- layer=1 filter=150 channel=57
    4, 5, -12, -7, 2, -9, -7, -3, 5,
    -- layer=1 filter=150 channel=58
    1, -1, 4, -1, 3, 8, 8, 0, -1,
    -- layer=1 filter=150 channel=59
    -12, -6, 7, -2, 6, -4, 2, 0, -10,
    -- layer=1 filter=150 channel=60
    5, -3, -8, -3, 8, 5, -3, -5, 9,
    -- layer=1 filter=150 channel=61
    -1, 1, 2, 9, 7, 0, -2, 10, 0,
    -- layer=1 filter=150 channel=62
    -1, 3, -8, 6, -7, 5, 7, 6, -8,
    -- layer=1 filter=150 channel=63
    3, -8, 0, -6, 3, 3, 7, -1, -2,
    -- layer=1 filter=150 channel=64
    0, 0, 0, 6, -1, 0, -4, 5, -7,
    -- layer=1 filter=150 channel=65
    4, -4, 3, 3, 1, -3, -2, 2, 6,
    -- layer=1 filter=150 channel=66
    -6, -1, -4, 7, 2, -9, -12, -4, 3,
    -- layer=1 filter=150 channel=67
    -3, 5, -1, 0, -6, 1, -5, 0, 5,
    -- layer=1 filter=150 channel=68
    2, -8, 8, -5, 5, 0, -4, -4, -1,
    -- layer=1 filter=150 channel=69
    -5, 8, 9, 4, 7, -6, 0, -3, 2,
    -- layer=1 filter=150 channel=70
    6, 6, 5, -2, -8, 8, -5, 7, -8,
    -- layer=1 filter=150 channel=71
    -7, -9, 6, -4, 0, -9, -2, 8, 10,
    -- layer=1 filter=150 channel=72
    -1, -10, 4, -8, -1, -5, 3, -3, 0,
    -- layer=1 filter=150 channel=73
    1, 4, -2, 0, -8, -8, 7, -9, 2,
    -- layer=1 filter=150 channel=74
    0, -6, -9, 5, 4, 6, 2, -10, -3,
    -- layer=1 filter=150 channel=75
    1, 4, -5, -4, 7, 0, 5, 0, 6,
    -- layer=1 filter=150 channel=76
    -8, -1, 5, -9, -10, 7, -11, 2, 0,
    -- layer=1 filter=150 channel=77
    -10, -7, 1, -12, -3, 6, 7, 7, 0,
    -- layer=1 filter=150 channel=78
    -7, -7, 3, -1, 5, -5, -7, -1, -12,
    -- layer=1 filter=150 channel=79
    -2, -6, -1, -5, -11, -10, 5, 5, -6,
    -- layer=1 filter=150 channel=80
    6, 7, 0, -10, 1, 6, 0, 4, 2,
    -- layer=1 filter=150 channel=81
    0, -9, -6, 5, -4, 3, 7, -3, -6,
    -- layer=1 filter=150 channel=82
    2, -3, 8, 0, 0, 10, -4, 11, -6,
    -- layer=1 filter=150 channel=83
    1, -6, 4, 3, -8, -4, -10, 2, -7,
    -- layer=1 filter=150 channel=84
    -9, 7, -4, 0, 3, 4, -1, -4, -5,
    -- layer=1 filter=150 channel=85
    3, -7, -4, 9, -3, 3, 3, -6, 2,
    -- layer=1 filter=150 channel=86
    -3, -9, -5, -1, -4, 3, 6, -12, -8,
    -- layer=1 filter=150 channel=87
    7, 4, -5, 3, 0, -11, 0, -5, -3,
    -- layer=1 filter=150 channel=88
    -6, 0, -3, -10, -10, 2, 3, -11, -8,
    -- layer=1 filter=150 channel=89
    5, 2, 1, 8, -4, -4, 6, 3, -4,
    -- layer=1 filter=150 channel=90
    -9, 4, -7, 0, -12, 5, 4, 8, -5,
    -- layer=1 filter=150 channel=91
    0, 2, 6, 4, -8, 0, -2, 5, 3,
    -- layer=1 filter=150 channel=92
    5, -6, 1, -5, 0, -3, 4, -5, -3,
    -- layer=1 filter=150 channel=93
    -3, -9, -5, 0, -4, -9, 4, -4, -9,
    -- layer=1 filter=150 channel=94
    0, -3, -11, 4, 2, 4, -11, 0, 3,
    -- layer=1 filter=150 channel=95
    -12, 0, -4, -5, -1, 4, 5, -11, -6,
    -- layer=1 filter=150 channel=96
    5, -4, 7, -11, -3, 4, 5, 5, 0,
    -- layer=1 filter=150 channel=97
    -4, -5, 4, 7, -10, 2, -7, -7, 0,
    -- layer=1 filter=150 channel=98
    -9, -3, -9, 5, -5, -11, 0, 3, 4,
    -- layer=1 filter=150 channel=99
    6, 5, 1, -7, -7, 8, 3, 6, 0,
    -- layer=1 filter=150 channel=100
    -10, -13, -4, 7, 0, -11, 6, -2, 7,
    -- layer=1 filter=150 channel=101
    6, -6, -11, -7, -11, -5, 6, 0, -5,
    -- layer=1 filter=150 channel=102
    6, -1, -5, 0, 3, 4, -10, -4, -4,
    -- layer=1 filter=150 channel=103
    3, -3, -3, -7, 2, -9, -1, -11, 6,
    -- layer=1 filter=150 channel=104
    -11, 4, -11, -7, -6, 0, -7, -2, -10,
    -- layer=1 filter=150 channel=105
    0, -11, -3, 4, 4, -5, -2, 1, -4,
    -- layer=1 filter=150 channel=106
    4, -4, -3, 0, -7, -7, 2, -3, 5,
    -- layer=1 filter=150 channel=107
    11, 5, -6, 4, 9, -3, -6, 6, 9,
    -- layer=1 filter=150 channel=108
    -2, -1, 7, 7, 2, -7, 2, 0, 5,
    -- layer=1 filter=150 channel=109
    -1, 1, 9, -7, -4, 5, 6, 0, -2,
    -- layer=1 filter=150 channel=110
    2, 5, -4, 0, 0, 7, -2, -7, 0,
    -- layer=1 filter=150 channel=111
    2, -4, -4, 5, -8, 2, -11, -14, -2,
    -- layer=1 filter=150 channel=112
    -10, 0, -8, -10, 4, 0, -12, -11, -10,
    -- layer=1 filter=150 channel=113
    0, -2, -13, 1, 1, 6, 0, 3, 7,
    -- layer=1 filter=150 channel=114
    -2, 5, 4, -12, 1, -6, -3, 5, 5,
    -- layer=1 filter=150 channel=115
    5, 4, -1, 5, -10, -1, -9, -6, 0,
    -- layer=1 filter=150 channel=116
    4, 5, 3, 0, 7, 2, -4, -5, 8,
    -- layer=1 filter=150 channel=117
    -12, -6, -11, 2, 6, -4, 0, -7, 1,
    -- layer=1 filter=150 channel=118
    4, -6, -2, 7, 3, 2, 4, 4, -3,
    -- layer=1 filter=150 channel=119
    -11, -7, 5, 1, 8, -7, -2, 0, 2,
    -- layer=1 filter=150 channel=120
    1, -8, 1, -7, 10, -1, 9, 5, 0,
    -- layer=1 filter=150 channel=121
    -2, 7, -1, 7, -7, -3, -7, 5, -1,
    -- layer=1 filter=150 channel=122
    -7, -4, -6, -9, -4, 3, 3, -3, 7,
    -- layer=1 filter=150 channel=123
    -6, 7, 0, -9, -3, -2, -2, -1, -7,
    -- layer=1 filter=150 channel=124
    0, 7, -5, 7, -6, -11, -11, -3, -12,
    -- layer=1 filter=150 channel=125
    9, -3, -7, -2, -3, 1, 4, 1, -6,
    -- layer=1 filter=150 channel=126
    0, -4, -3, 9, 7, -3, -1, 0, 4,
    -- layer=1 filter=150 channel=127
    -8, 8, -3, -4, 3, -8, 0, -3, 2,
    -- layer=1 filter=151 channel=0
    3, -9, -5, 2, 2, -7, 0, 8, 2,
    -- layer=1 filter=151 channel=1
    -2, 3, 4, 4, 6, 7, 2, -5, 7,
    -- layer=1 filter=151 channel=2
    -6, -6, 6, -4, 4, -8, 7, 1, 4,
    -- layer=1 filter=151 channel=3
    0, -6, -2, 0, 4, -2, 4, 8, -7,
    -- layer=1 filter=151 channel=4
    -8, 4, -9, -10, -2, 4, 0, -10, -8,
    -- layer=1 filter=151 channel=5
    -2, 5, -10, -1, -11, 7, 0, -5, -2,
    -- layer=1 filter=151 channel=6
    9, 10, 0, -1, -6, -2, -5, 1, 4,
    -- layer=1 filter=151 channel=7
    0, 3, -1, -1, -3, -7, 2, -10, 1,
    -- layer=1 filter=151 channel=8
    -10, 6, -2, -6, 8, 2, 2, 4, -5,
    -- layer=1 filter=151 channel=9
    -5, 7, -2, 4, -6, -1, 4, -3, 2,
    -- layer=1 filter=151 channel=10
    -8, 1, -7, -2, 6, -2, -13, -3, -9,
    -- layer=1 filter=151 channel=11
    3, -10, 0, 5, 1, -5, -7, 4, -4,
    -- layer=1 filter=151 channel=12
    5, -2, 0, -8, 1, 5, 8, -7, 0,
    -- layer=1 filter=151 channel=13
    2, 3, -2, -8, 3, -9, 1, -10, -7,
    -- layer=1 filter=151 channel=14
    -5, -5, -5, -2, 0, -5, -1, 5, 0,
    -- layer=1 filter=151 channel=15
    10, 0, -6, 10, 4, 3, 3, -10, -9,
    -- layer=1 filter=151 channel=16
    -6, 5, -10, 5, -5, -8, 2, -2, -2,
    -- layer=1 filter=151 channel=17
    7, 1, 8, 0, -11, -5, 3, -5, -6,
    -- layer=1 filter=151 channel=18
    -10, 0, 0, -1, -3, 5, -7, -7, 0,
    -- layer=1 filter=151 channel=19
    0, 2, -1, -4, 3, 3, 3, 1, -9,
    -- layer=1 filter=151 channel=20
    -8, -5, 0, -1, -6, -8, -12, 3, 5,
    -- layer=1 filter=151 channel=21
    3, -4, -5, -4, -3, -9, 7, 1, 0,
    -- layer=1 filter=151 channel=22
    0, 7, -5, -2, -3, 4, -10, 8, -6,
    -- layer=1 filter=151 channel=23
    4, 5, -8, -2, -2, -11, 5, -6, 6,
    -- layer=1 filter=151 channel=24
    7, -3, -3, 2, -4, -9, 6, -1, -6,
    -- layer=1 filter=151 channel=25
    -3, -7, 6, -13, 9, -8, -8, -9, -3,
    -- layer=1 filter=151 channel=26
    -7, -11, -13, -5, 5, 2, 6, -3, -6,
    -- layer=1 filter=151 channel=27
    1, 0, -8, -9, 3, 6, 6, 4, -7,
    -- layer=1 filter=151 channel=28
    1, -4, -3, 5, -10, 4, -3, -7, 5,
    -- layer=1 filter=151 channel=29
    -2, 1, 10, -2, -1, 4, -4, -11, 0,
    -- layer=1 filter=151 channel=30
    -6, 2, 4, 0, 1, -6, 7, -5, -6,
    -- layer=1 filter=151 channel=31
    0, 0, 0, -9, 4, 3, -12, -1, 3,
    -- layer=1 filter=151 channel=32
    6, -11, 5, -4, -12, -7, -3, -3, -2,
    -- layer=1 filter=151 channel=33
    -10, -3, 0, -4, -6, 7, 0, -6, -5,
    -- layer=1 filter=151 channel=34
    0, 2, -2, -2, 5, 3, -5, 6, -2,
    -- layer=1 filter=151 channel=35
    -8, 0, -2, -3, 1, 6, -2, -7, 7,
    -- layer=1 filter=151 channel=36
    -1, 4, 8, 3, -9, 6, 6, 0, -6,
    -- layer=1 filter=151 channel=37
    -6, 4, 5, -9, 0, -7, -1, -8, 1,
    -- layer=1 filter=151 channel=38
    0, -6, -10, -11, -4, -9, 2, -7, 4,
    -- layer=1 filter=151 channel=39
    8, 2, 4, 0, 2, -1, 7, 0, 0,
    -- layer=1 filter=151 channel=40
    -1, -4, 5, -9, -1, -8, 6, -11, 1,
    -- layer=1 filter=151 channel=41
    -1, -2, -1, 2, -8, 4, 7, 6, 4,
    -- layer=1 filter=151 channel=42
    0, -1, -3, -10, -5, 1, 8, -2, -3,
    -- layer=1 filter=151 channel=43
    7, 1, -2, 5, 8, -1, 3, 0, 0,
    -- layer=1 filter=151 channel=44
    3, -11, -1, 0, 5, 1, -5, -4, -1,
    -- layer=1 filter=151 channel=45
    -5, -11, -5, -5, 0, -10, -5, 8, 6,
    -- layer=1 filter=151 channel=46
    -7, 8, 2, 9, 4, -12, 0, 8, 0,
    -- layer=1 filter=151 channel=47
    -3, -6, 4, 4, 0, 6, -2, -1, -6,
    -- layer=1 filter=151 channel=48
    0, -5, -3, -5, -2, -3, -7, -9, 0,
    -- layer=1 filter=151 channel=49
    -9, -5, 1, 3, -9, -1, -5, 2, 7,
    -- layer=1 filter=151 channel=50
    -6, -3, 6, 0, 0, 8, 0, -6, -1,
    -- layer=1 filter=151 channel=51
    -8, -4, -3, 2, -1, 3, -3, 0, 1,
    -- layer=1 filter=151 channel=52
    6, -6, 10, 2, 10, 0, -1, -9, -1,
    -- layer=1 filter=151 channel=53
    8, -3, -9, -5, 6, -6, -10, -8, -2,
    -- layer=1 filter=151 channel=54
    -10, 0, -8, -1, 1, 2, 7, 3, -9,
    -- layer=1 filter=151 channel=55
    -2, -1, -7, -4, -13, 4, -11, 4, -10,
    -- layer=1 filter=151 channel=56
    0, 3, 3, 1, -9, 6, -7, -9, -2,
    -- layer=1 filter=151 channel=57
    -2, 5, -6, -11, 0, -4, 7, 4, -11,
    -- layer=1 filter=151 channel=58
    4, 1, 8, 4, -7, 3, -6, -9, -1,
    -- layer=1 filter=151 channel=59
    -2, 3, 4, -11, 0, 4, -8, 7, -2,
    -- layer=1 filter=151 channel=60
    1, 0, 5, 4, -5, 9, -3, 6, 8,
    -- layer=1 filter=151 channel=61
    0, 1, 10, 2, -8, -6, -7, -6, 0,
    -- layer=1 filter=151 channel=62
    3, -8, -3, -2, -3, -10, -7, 1, -1,
    -- layer=1 filter=151 channel=63
    -8, -4, 1, 0, -6, -9, 8, -4, -7,
    -- layer=1 filter=151 channel=64
    8, 8, 2, 6, 3, 0, -9, 0, 0,
    -- layer=1 filter=151 channel=65
    -5, -10, 4, -6, 2, -5, 0, -5, 6,
    -- layer=1 filter=151 channel=66
    7, 1, -7, -7, 4, -11, -9, -7, -2,
    -- layer=1 filter=151 channel=67
    -4, -9, -6, -1, -9, 4, -8, 4, -6,
    -- layer=1 filter=151 channel=68
    7, -6, 0, 2, 4, -8, 2, 4, 1,
    -- layer=1 filter=151 channel=69
    2, -12, 8, -11, 6, -6, 7, -10, 4,
    -- layer=1 filter=151 channel=70
    -8, 3, -5, 10, 6, 9, -6, 2, -8,
    -- layer=1 filter=151 channel=71
    -5, -9, 1, -10, 6, -4, -3, 5, 4,
    -- layer=1 filter=151 channel=72
    -7, -5, -9, -8, 0, -6, 4, -1, 3,
    -- layer=1 filter=151 channel=73
    3, -5, -9, -8, 3, -11, 0, -9, -1,
    -- layer=1 filter=151 channel=74
    5, -5, -8, -11, 7, -5, -7, -2, -7,
    -- layer=1 filter=151 channel=75
    -8, 5, 0, 7, -10, 3, -1, 3, 3,
    -- layer=1 filter=151 channel=76
    -10, 0, 0, 2, -10, 5, 3, 4, -8,
    -- layer=1 filter=151 channel=77
    -1, 8, 7, 0, 7, -1, -8, -7, -11,
    -- layer=1 filter=151 channel=78
    4, -1, -8, -10, -3, -8, -6, -9, 1,
    -- layer=1 filter=151 channel=79
    8, -12, -1, -12, 6, -3, 4, 5, -4,
    -- layer=1 filter=151 channel=80
    1, 4, -11, 8, -10, -7, 8, 7, 4,
    -- layer=1 filter=151 channel=81
    0, -6, 2, -9, -3, -5, -9, 1, -6,
    -- layer=1 filter=151 channel=82
    -10, 8, 7, -2, 8, 7, 0, -9, -5,
    -- layer=1 filter=151 channel=83
    -1, 4, 6, -10, 0, -5, 2, 2, -1,
    -- layer=1 filter=151 channel=84
    0, 6, -10, 4, -11, 3, 6, -3, 4,
    -- layer=1 filter=151 channel=85
    -1, -7, -7, 4, 4, 3, -7, -9, 4,
    -- layer=1 filter=151 channel=86
    4, -4, 3, -8, -11, 0, 8, 5, 3,
    -- layer=1 filter=151 channel=87
    7, 7, -10, 6, -1, 7, -11, 0, -2,
    -- layer=1 filter=151 channel=88
    -6, -3, 1, 4, 2, 7, -4, -10, 3,
    -- layer=1 filter=151 channel=89
    -12, -1, -10, -12, 6, 0, -6, 2, -4,
    -- layer=1 filter=151 channel=90
    0, -12, -9, -5, 2, -2, -7, -8, 4,
    -- layer=1 filter=151 channel=91
    -4, -7, -9, -2, -9, 6, 0, 3, -6,
    -- layer=1 filter=151 channel=92
    -5, -7, -3, -10, -11, -5, -1, 4, 0,
    -- layer=1 filter=151 channel=93
    -11, -11, -1, 2, -10, -10, -7, -7, -12,
    -- layer=1 filter=151 channel=94
    6, -9, -1, 0, -6, 8, -6, 0, 4,
    -- layer=1 filter=151 channel=95
    0, -2, 8, -1, -6, 5, 7, -3, 1,
    -- layer=1 filter=151 channel=96
    -5, 2, 5, -11, 2, -9, -10, -1, 5,
    -- layer=1 filter=151 channel=97
    -6, 8, 2, -5, -4, -7, -3, -4, 0,
    -- layer=1 filter=151 channel=98
    4, -3, -7, -15, -4, -1, -2, 8, -8,
    -- layer=1 filter=151 channel=99
    -4, -2, -4, 3, 3, -10, 4, 5, 4,
    -- layer=1 filter=151 channel=100
    7, -11, -7, -8, 7, 0, -9, -7, 6,
    -- layer=1 filter=151 channel=101
    -6, -5, -2, 1, -1, -8, 7, 7, 4,
    -- layer=1 filter=151 channel=102
    -1, 6, -3, -9, -5, -7, -10, 0, 4,
    -- layer=1 filter=151 channel=103
    -8, -4, -10, 7, -2, -8, 2, -4, 7,
    -- layer=1 filter=151 channel=104
    1, -7, 0, 8, 9, -1, -7, -8, 5,
    -- layer=1 filter=151 channel=105
    7, 6, 6, -9, -11, 7, 1, -3, 1,
    -- layer=1 filter=151 channel=106
    2, 6, -11, 6, -10, -5, 3, 3, -5,
    -- layer=1 filter=151 channel=107
    8, -6, 10, -10, 8, 8, 1, 4, 4,
    -- layer=1 filter=151 channel=108
    2, -6, -8, -7, 1, 2, -2, -3, 9,
    -- layer=1 filter=151 channel=109
    5, 2, -11, -6, 6, -3, 4, 3, 8,
    -- layer=1 filter=151 channel=110
    4, -4, -1, 0, -7, -3, -11, -9, 6,
    -- layer=1 filter=151 channel=111
    2, 8, -8, 1, 6, 2, -5, -10, -4,
    -- layer=1 filter=151 channel=112
    -6, -6, -11, -9, -11, -11, 0, -6, 0,
    -- layer=1 filter=151 channel=113
    -5, -9, 3, 7, 1, -7, -9, 6, 3,
    -- layer=1 filter=151 channel=114
    0, -8, -10, -5, 1, -4, -4, 0, -12,
    -- layer=1 filter=151 channel=115
    6, 0, 0, 6, 1, -4, -3, 2, -10,
    -- layer=1 filter=151 channel=116
    -3, 1, 1, -4, 3, -6, 9, -4, -11,
    -- layer=1 filter=151 channel=117
    8, -7, -2, 0, -7, 0, 6, 6, -8,
    -- layer=1 filter=151 channel=118
    -11, -8, -2, -1, -5, 0, 4, 0, -3,
    -- layer=1 filter=151 channel=119
    1, -4, 1, 5, -5, 0, 9, -4, -4,
    -- layer=1 filter=151 channel=120
    2, 1, -10, 5, -3, 3, 3, -6, -1,
    -- layer=1 filter=151 channel=121
    0, -8, 6, 0, -7, -7, -11, -1, 6,
    -- layer=1 filter=151 channel=122
    1, 6, 2, 2, 9, 7, -10, 4, 0,
    -- layer=1 filter=151 channel=123
    0, -10, 4, -5, -10, -8, -6, 0, -8,
    -- layer=1 filter=151 channel=124
    0, 6, 2, -7, -1, -7, -3, 1, 2,
    -- layer=1 filter=151 channel=125
    -5, -1, 0, 0, -10, 7, 7, -6, 3,
    -- layer=1 filter=151 channel=126
    0, -6, -2, 4, 0, -11, 3, -4, 8,
    -- layer=1 filter=151 channel=127
    -7, -3, -13, -7, 1, -2, -10, -4, -6,
    -- layer=1 filter=152 channel=0
    4, -5, 0, -7, -11, -11, -6, 1, -8,
    -- layer=1 filter=152 channel=1
    -3, -2, 0, 5, 4, 5, 8, -2, -5,
    -- layer=1 filter=152 channel=2
    6, 6, -4, 2, -4, 5, 0, -1, -9,
    -- layer=1 filter=152 channel=3
    1, -5, 1, 1, -2, 3, 0, 2, -3,
    -- layer=1 filter=152 channel=4
    -10, 0, -5, -3, 0, -9, -6, -6, -11,
    -- layer=1 filter=152 channel=5
    5, 0, -5, 2, 0, -10, -2, 10, 0,
    -- layer=1 filter=152 channel=6
    -9, -1, 3, 0, -6, 6, 0, 2, 2,
    -- layer=1 filter=152 channel=7
    -7, -6, -2, 5, -10, 8, 6, 4, 0,
    -- layer=1 filter=152 channel=8
    6, -1, 3, 5, -10, -11, -3, 0, -7,
    -- layer=1 filter=152 channel=9
    0, -5, 5, -9, -6, -3, -2, 0, -13,
    -- layer=1 filter=152 channel=10
    3, -3, 1, 3, -7, -11, -2, -8, -11,
    -- layer=1 filter=152 channel=11
    -3, 0, 0, 8, 5, -11, 0, -5, 2,
    -- layer=1 filter=152 channel=12
    -6, 8, -4, 3, 0, -10, 10, 11, -10,
    -- layer=1 filter=152 channel=13
    2, -3, -11, 4, 5, -11, 4, -2, 6,
    -- layer=1 filter=152 channel=14
    0, -4, 0, 3, -7, -10, 3, 3, 0,
    -- layer=1 filter=152 channel=15
    0, -7, -11, -2, -1, -5, -1, -5, -7,
    -- layer=1 filter=152 channel=16
    -8, 4, -4, -2, -11, -12, 5, -11, 4,
    -- layer=1 filter=152 channel=17
    3, 0, -11, -12, -7, 0, -1, -7, 1,
    -- layer=1 filter=152 channel=18
    5, 0, -3, -11, -11, 0, 3, 7, -11,
    -- layer=1 filter=152 channel=19
    3, 6, -7, 6, 1, -7, -10, 0, -6,
    -- layer=1 filter=152 channel=20
    0, -5, -7, -2, -5, 0, 0, 6, -3,
    -- layer=1 filter=152 channel=21
    4, -3, -7, 1, -3, 6, 3, -4, -9,
    -- layer=1 filter=152 channel=22
    -11, -6, 7, -6, 3, -7, -10, 6, 5,
    -- layer=1 filter=152 channel=23
    -3, 6, -6, -2, -10, -9, 6, -3, 4,
    -- layer=1 filter=152 channel=24
    -13, 2, -10, 0, -3, -5, -4, -6, -6,
    -- layer=1 filter=152 channel=25
    -8, 5, -5, -2, 6, -1, 5, -11, -9,
    -- layer=1 filter=152 channel=26
    6, -10, -14, 3, 3, 8, 5, -12, 0,
    -- layer=1 filter=152 channel=27
    5, -10, -5, 4, 8, 6, 6, 8, 2,
    -- layer=1 filter=152 channel=28
    -12, -11, 0, 2, 9, 8, -6, -10, 5,
    -- layer=1 filter=152 channel=29
    -3, -7, -11, -10, 6, 7, -12, -1, -4,
    -- layer=1 filter=152 channel=30
    -6, 11, 11, -9, -2, 0, -4, 1, 7,
    -- layer=1 filter=152 channel=31
    9, 7, -10, -8, 0, -2, -3, 0, -2,
    -- layer=1 filter=152 channel=32
    -4, -5, 2, 0, 0, -7, 5, 6, 6,
    -- layer=1 filter=152 channel=33
    1, -7, -12, 0, -7, 7, 5, -5, 10,
    -- layer=1 filter=152 channel=34
    6, -6, 0, -3, 1, -7, -9, 0, -4,
    -- layer=1 filter=152 channel=35
    3, 3, 5, -1, 2, 2, 1, -5, -11,
    -- layer=1 filter=152 channel=36
    3, 6, -3, -9, -10, 7, 7, -10, -7,
    -- layer=1 filter=152 channel=37
    4, 8, -7, -11, -9, 6, 10, -4, 10,
    -- layer=1 filter=152 channel=38
    -2, -12, -5, 0, -1, 7, -11, -10, 1,
    -- layer=1 filter=152 channel=39
    -4, 0, -5, 8, 7, 0, -10, -7, -4,
    -- layer=1 filter=152 channel=40
    3, -1, -5, 12, 3, 4, -10, -7, -9,
    -- layer=1 filter=152 channel=41
    5, -4, 4, 5, 0, 1, 0, 0, 2,
    -- layer=1 filter=152 channel=42
    -8, 10, 5, -8, -4, -7, -7, 6, 4,
    -- layer=1 filter=152 channel=43
    -6, 3, -2, -1, -4, 6, -2, -3, -1,
    -- layer=1 filter=152 channel=44
    3, 1, 9, 6, -3, 8, 5, -2, -3,
    -- layer=1 filter=152 channel=45
    -6, -4, -10, 0, 3, -1, -3, 3, -12,
    -- layer=1 filter=152 channel=46
    -3, -1, 3, -9, 2, 7, 10, 9, 2,
    -- layer=1 filter=152 channel=47
    -7, -6, -5, 5, -7, 4, -10, -11, -6,
    -- layer=1 filter=152 channel=48
    -1, -3, 6, -8, -4, 1, 0, 7, 4,
    -- layer=1 filter=152 channel=49
    6, -11, -5, -10, -9, 0, 5, -1, 0,
    -- layer=1 filter=152 channel=50
    0, -1, 6, 0, -8, -1, -10, -12, 0,
    -- layer=1 filter=152 channel=51
    4, 4, -5, -5, 5, 7, -5, -10, -2,
    -- layer=1 filter=152 channel=52
    0, -8, -9, -12, -10, 7, 5, -6, -10,
    -- layer=1 filter=152 channel=53
    -12, 7, -11, 0, 8, -2, 1, 8, 7,
    -- layer=1 filter=152 channel=54
    -7, 1, 3, -11, -12, 1, 9, -8, -1,
    -- layer=1 filter=152 channel=55
    -1, -6, 8, -12, 5, 6, -5, 11, -7,
    -- layer=1 filter=152 channel=56
    -2, -1, -1, -7, 0, -11, 0, 8, -10,
    -- layer=1 filter=152 channel=57
    6, -7, 1, 2, -8, 3, 6, -6, -3,
    -- layer=1 filter=152 channel=58
    5, 0, 4, 3, 3, -9, -10, 7, -1,
    -- layer=1 filter=152 channel=59
    6, -11, -1, -2, -8, -4, 8, -6, 1,
    -- layer=1 filter=152 channel=60
    10, -7, -7, -8, 4, 2, 1, -7, -1,
    -- layer=1 filter=152 channel=61
    8, 1, -8, -2, 7, -1, 3, 0, -4,
    -- layer=1 filter=152 channel=62
    -5, 5, -3, -7, -3, -5, 8, 7, 3,
    -- layer=1 filter=152 channel=63
    2, -5, 4, -3, 2, 0, -6, -2, -6,
    -- layer=1 filter=152 channel=64
    -5, -8, -1, 7, -3, 6, -2, 6, 3,
    -- layer=1 filter=152 channel=65
    -5, -8, -7, 1, -8, 2, -1, 8, 8,
    -- layer=1 filter=152 channel=66
    -4, 7, -10, -1, 8, -7, -9, -12, -12,
    -- layer=1 filter=152 channel=67
    -11, -3, 5, 8, -9, -8, -10, 4, -6,
    -- layer=1 filter=152 channel=68
    4, -5, 3, -11, -7, 2, -4, 6, -5,
    -- layer=1 filter=152 channel=69
    0, -1, -11, 5, -13, -3, -2, 0, 4,
    -- layer=1 filter=152 channel=70
    4, 4, -11, -8, 2, -7, -10, 7, 8,
    -- layer=1 filter=152 channel=71
    -3, -2, -6, 5, -5, 0, 5, -2, 7,
    -- layer=1 filter=152 channel=72
    -5, 3, -11, -7, 7, -5, 0, 6, 2,
    -- layer=1 filter=152 channel=73
    -9, -4, -5, 4, -4, 6, -8, 7, -11,
    -- layer=1 filter=152 channel=74
    8, 2, -8, -3, -1, 1, 2, 3, -12,
    -- layer=1 filter=152 channel=75
    -8, -5, 3, 8, 4, 3, -10, -12, -12,
    -- layer=1 filter=152 channel=76
    6, -11, 9, 4, 0, 3, 0, 4, 0,
    -- layer=1 filter=152 channel=77
    -9, -6, -7, 2, 6, 7, -9, -7, 8,
    -- layer=1 filter=152 channel=78
    -4, 2, 0, -5, 3, -3, -10, 1, 6,
    -- layer=1 filter=152 channel=79
    2, -3, -1, -11, 3, -4, -6, -4, 0,
    -- layer=1 filter=152 channel=80
    -5, -8, 0, -9, 8, 0, 7, 0, -8,
    -- layer=1 filter=152 channel=81
    4, -7, -9, 6, -9, 3, -2, 2, -4,
    -- layer=1 filter=152 channel=82
    1, 6, -12, 0, -5, -8, 7, 0, 3,
    -- layer=1 filter=152 channel=83
    -1, -1, -2, 4, 4, -7, -10, -3, 8,
    -- layer=1 filter=152 channel=84
    -6, 0, 0, 5, 5, 4, -10, -8, 0,
    -- layer=1 filter=152 channel=85
    3, 3, 1, -1, -4, -11, -7, 1, -8,
    -- layer=1 filter=152 channel=86
    3, 5, 3, 1, -3, -4, -1, -3, 6,
    -- layer=1 filter=152 channel=87
    5, 0, 3, 3, -1, 2, 4, -4, 3,
    -- layer=1 filter=152 channel=88
    3, -13, 1, 3, -13, 1, -14, 3, -11,
    -- layer=1 filter=152 channel=89
    7, 2, 5, 4, -1, 0, 2, 1, 5,
    -- layer=1 filter=152 channel=90
    -2, -4, -7, 2, -8, 0, -2, 0, 7,
    -- layer=1 filter=152 channel=91
    5, -4, -7, 7, -8, 4, 0, 3, 4,
    -- layer=1 filter=152 channel=92
    0, -10, -3, 8, -4, -1, -11, -4, 0,
    -- layer=1 filter=152 channel=93
    3, -12, 7, 7, -9, 1, -9, 6, -1,
    -- layer=1 filter=152 channel=94
    5, 2, -5, 6, 2, -5, -4, 6, -7,
    -- layer=1 filter=152 channel=95
    2, 5, 0, 3, -9, -6, -2, -7, 5,
    -- layer=1 filter=152 channel=96
    5, -6, 7, 6, 4, -10, 0, 9, 7,
    -- layer=1 filter=152 channel=97
    -10, 0, -4, -9, 5, 0, 1, -10, -2,
    -- layer=1 filter=152 channel=98
    -10, 1, 4, -5, -10, 0, 6, -5, -5,
    -- layer=1 filter=152 channel=99
    5, -8, 1, -10, -10, -6, -4, 4, 8,
    -- layer=1 filter=152 channel=100
    -5, -10, -8, -10, -8, 7, -4, 7, -8,
    -- layer=1 filter=152 channel=101
    8, -8, -10, -11, 6, 1, 0, -11, -5,
    -- layer=1 filter=152 channel=102
    -8, 0, 9, -5, -6, -9, 5, -5, 3,
    -- layer=1 filter=152 channel=103
    2, -2, -9, 6, -8, -9, -7, 4, 8,
    -- layer=1 filter=152 channel=104
    5, 8, -7, -7, -3, -6, 2, -1, -4,
    -- layer=1 filter=152 channel=105
    5, 7, 1, -7, -12, -12, -9, -8, 3,
    -- layer=1 filter=152 channel=106
    -11, -8, -7, 6, -2, 7, 0, -4, 1,
    -- layer=1 filter=152 channel=107
    -7, 0, -3, -7, -3, -2, 5, 2, 5,
    -- layer=1 filter=152 channel=108
    0, -4, 5, -4, 3, 4, 4, -8, -3,
    -- layer=1 filter=152 channel=109
    -8, -3, 6, -3, 0, -5, 0, 8, 7,
    -- layer=1 filter=152 channel=110
    7, -2, 3, -1, 5, 0, 1, -10, 4,
    -- layer=1 filter=152 channel=111
    -11, 0, -11, 5, -3, -3, 5, -9, 2,
    -- layer=1 filter=152 channel=112
    -11, 6, 6, -2, 5, -2, 2, -11, -4,
    -- layer=1 filter=152 channel=113
    -8, 1, -5, 0, -11, 3, 0, 3, 7,
    -- layer=1 filter=152 channel=114
    -7, 8, -7, 5, 9, 7, -4, 10, -9,
    -- layer=1 filter=152 channel=115
    -9, -11, 2, -8, 3, 7, -8, -7, 0,
    -- layer=1 filter=152 channel=116
    0, -3, 0, 4, -7, 7, 6, 6, -11,
    -- layer=1 filter=152 channel=117
    -7, -4, 7, 7, -8, 6, 4, -2, -5,
    -- layer=1 filter=152 channel=118
    8, 5, 4, 7, 7, -9, -7, -6, 1,
    -- layer=1 filter=152 channel=119
    2, -6, 8, 0, -12, -10, -5, -11, -2,
    -- layer=1 filter=152 channel=120
    -11, -7, -1, -5, -7, 3, -8, -5, 4,
    -- layer=1 filter=152 channel=121
    6, -4, -9, -2, 5, 0, 3, -6, -4,
    -- layer=1 filter=152 channel=122
    -9, -4, -1, -3, -7, 4, 1, 7, 5,
    -- layer=1 filter=152 channel=123
    -11, 6, -8, 0, -10, -3, 6, -7, -7,
    -- layer=1 filter=152 channel=124
    4, -3, -8, 0, -4, -1, -5, -10, 3,
    -- layer=1 filter=152 channel=125
    0, -1, -1, 0, 6, 3, 4, -1, 4,
    -- layer=1 filter=152 channel=126
    -5, 6, 2, 7, 1, -2, -7, 1, 3,
    -- layer=1 filter=152 channel=127
    -7, 0, 3, -8, 4, -1, -7, -5, 4,
    -- layer=1 filter=153 channel=0
    -9, -5, -6, -6, 1, -7, -5, -11, -2,
    -- layer=1 filter=153 channel=1
    -6, 6, -8, -2, 7, -4, 0, -9, -4,
    -- layer=1 filter=153 channel=2
    -3, -6, 7, -4, -10, -11, 6, -1, 6,
    -- layer=1 filter=153 channel=3
    1, -9, -8, -8, -1, 10, 9, -1, 4,
    -- layer=1 filter=153 channel=4
    -11, -2, 1, 1, 7, -6, -11, 3, 5,
    -- layer=1 filter=153 channel=5
    2, -3, -1, -1, -2, -2, -10, -5, -6,
    -- layer=1 filter=153 channel=6
    0, 0, -9, -10, -7, -1, -5, -4, -5,
    -- layer=1 filter=153 channel=7
    -9, 2, 0, -12, -3, -6, -5, -4, 4,
    -- layer=1 filter=153 channel=8
    1, -5, 7, 6, 5, -6, -2, 1, 7,
    -- layer=1 filter=153 channel=9
    6, -6, 4, 5, 1, -8, -9, 9, 0,
    -- layer=1 filter=153 channel=10
    0, 0, -2, 0, -12, -8, 5, 3, -1,
    -- layer=1 filter=153 channel=11
    -3, 6, 2, -4, -10, -8, 7, -8, -8,
    -- layer=1 filter=153 channel=12
    7, 1, 0, 0, -9, -5, -6, 3, -8,
    -- layer=1 filter=153 channel=13
    0, -8, 4, -6, -7, -3, 0, -7, 2,
    -- layer=1 filter=153 channel=14
    6, -7, 6, -13, 1, -4, 2, -7, -4,
    -- layer=1 filter=153 channel=15
    7, 5, 11, 5, 2, 9, 2, 9, -12,
    -- layer=1 filter=153 channel=16
    3, 0, -10, 2, 8, -3, -4, 2, 3,
    -- layer=1 filter=153 channel=17
    -7, -6, 2, -8, -8, 4, 4, -3, 8,
    -- layer=1 filter=153 channel=18
    7, -8, 8, 5, 11, -5, -1, -5, -5,
    -- layer=1 filter=153 channel=19
    -5, 0, -4, -7, -1, -8, 9, -9, 7,
    -- layer=1 filter=153 channel=20
    -4, -9, -6, -3, 4, -6, -1, 2, 8,
    -- layer=1 filter=153 channel=21
    -4, -8, -8, 0, 7, 0, 6, 5, -11,
    -- layer=1 filter=153 channel=22
    -3, 4, 3, -11, 3, -3, -6, 3, -7,
    -- layer=1 filter=153 channel=23
    0, -7, 5, -4, 8, -6, 7, -8, 3,
    -- layer=1 filter=153 channel=24
    -9, 5, 7, 0, 6, 0, -5, 3, 1,
    -- layer=1 filter=153 channel=25
    3, 4, -6, 7, -5, 0, -12, -8, 4,
    -- layer=1 filter=153 channel=26
    3, -8, -7, -3, 10, 2, 3, 4, -5,
    -- layer=1 filter=153 channel=27
    7, -8, -1, 2, 4, -8, 0, 2, -2,
    -- layer=1 filter=153 channel=28
    1, -11, 6, -2, -4, 7, 1, -11, -11,
    -- layer=1 filter=153 channel=29
    -4, 4, -3, -5, -6, 6, 0, 0, 8,
    -- layer=1 filter=153 channel=30
    5, 2, -1, 6, 0, 1, 0, 8, -3,
    -- layer=1 filter=153 channel=31
    10, -8, -2, -4, 4, 3, 0, -4, 9,
    -- layer=1 filter=153 channel=32
    0, -4, 6, -6, 4, 7, -1, -11, -5,
    -- layer=1 filter=153 channel=33
    -6, -10, 9, -7, -2, -3, 10, -4, -9,
    -- layer=1 filter=153 channel=34
    6, -10, -5, -10, -11, 4, 8, 8, 4,
    -- layer=1 filter=153 channel=35
    5, -7, -5, -8, 6, 0, 3, -6, 3,
    -- layer=1 filter=153 channel=36
    -6, 5, 1, -4, -8, -1, -8, 3, 1,
    -- layer=1 filter=153 channel=37
    0, 3, -9, 2, -2, -7, -7, -2, 6,
    -- layer=1 filter=153 channel=38
    -8, -3, 1, -7, -11, 2, -3, 3, 5,
    -- layer=1 filter=153 channel=39
    -3, -4, 4, -6, 0, -11, -9, 1, -9,
    -- layer=1 filter=153 channel=40
    4, 3, 8, -3, -8, -4, 0, -4, 3,
    -- layer=1 filter=153 channel=41
    2, 2, -9, 7, -2, -7, -8, -3, -4,
    -- layer=1 filter=153 channel=42
    4, -12, 0, -3, 3, 3, 2, -10, 1,
    -- layer=1 filter=153 channel=43
    1, -3, 3, -10, -9, 5, 8, -7, -11,
    -- layer=1 filter=153 channel=44
    7, 6, 7, -9, 7, 1, 7, -4, -5,
    -- layer=1 filter=153 channel=45
    5, 8, -1, -1, -1, 6, -5, -12, 5,
    -- layer=1 filter=153 channel=46
    4, 7, -1, 7, -6, 5, -11, -5, 7,
    -- layer=1 filter=153 channel=47
    -11, 5, -8, 8, 5, -8, 3, 4, -3,
    -- layer=1 filter=153 channel=48
    1, -7, 1, 3, 6, -11, -6, -4, -6,
    -- layer=1 filter=153 channel=49
    -6, -5, 6, 1, -10, 1, -9, 0, 2,
    -- layer=1 filter=153 channel=50
    7, 5, 8, 4, 0, 0, 3, 2, 6,
    -- layer=1 filter=153 channel=51
    -10, 3, 2, 2, -4, 4, -6, 8, -7,
    -- layer=1 filter=153 channel=52
    10, -2, 6, 1, 7, -9, -2, 0, 1,
    -- layer=1 filter=153 channel=53
    5, -11, -4, 0, -2, -8, -11, -9, -2,
    -- layer=1 filter=153 channel=54
    -5, 0, -10, 4, 5, 6, -9, -2, 2,
    -- layer=1 filter=153 channel=55
    0, -6, 8, 4, -5, -12, -8, -11, 5,
    -- layer=1 filter=153 channel=56
    5, -7, 3, 8, -6, -1, 0, 0, -6,
    -- layer=1 filter=153 channel=57
    -7, 0, -2, 5, 6, -8, 7, -10, -1,
    -- layer=1 filter=153 channel=58
    4, 2, 2, 3, -4, 3, 5, 3, 5,
    -- layer=1 filter=153 channel=59
    -2, -4, 0, 1, -1, 0, 5, -8, -9,
    -- layer=1 filter=153 channel=60
    9, 0, 10, 4, 3, 8, 10, 1, 6,
    -- layer=1 filter=153 channel=61
    -3, 0, -6, -9, -7, 4, 9, 0, -4,
    -- layer=1 filter=153 channel=62
    -7, 2, 0, -7, 0, -9, -1, -6, -8,
    -- layer=1 filter=153 channel=63
    -9, -7, 4, 2, 5, 5, -2, 0, -10,
    -- layer=1 filter=153 channel=64
    2, -3, -1, -4, -11, -7, 1, 2, 0,
    -- layer=1 filter=153 channel=65
    -11, -2, 2, 7, 8, 6, 0, -2, -1,
    -- layer=1 filter=153 channel=66
    -2, -9, -7, -1, -1, 7, -11, 4, 0,
    -- layer=1 filter=153 channel=67
    4, -10, 0, 5, -2, 4, -9, 9, -4,
    -- layer=1 filter=153 channel=68
    8, 7, -2, -8, -8, 4, 6, -7, 8,
    -- layer=1 filter=153 channel=69
    1, 5, -5, 5, -10, -1, 6, 5, 0,
    -- layer=1 filter=153 channel=70
    7, 5, 8, -4, 3, -8, -7, -10, 3,
    -- layer=1 filter=153 channel=71
    -7, -9, 2, 5, 5, 3, -3, 6, 1,
    -- layer=1 filter=153 channel=72
    8, -6, 7, -2, 0, -10, -8, -9, -10,
    -- layer=1 filter=153 channel=73
    -2, 0, -10, -1, 0, -1, -11, -5, 2,
    -- layer=1 filter=153 channel=74
    4, -1, 8, -10, -8, 0, 0, 1, -6,
    -- layer=1 filter=153 channel=75
    -7, -10, 7, -10, 9, 2, 0, 0, -3,
    -- layer=1 filter=153 channel=76
    -6, 3, -2, -8, -8, -7, 3, -8, 0,
    -- layer=1 filter=153 channel=77
    7, -8, 8, -7, -5, 0, -1, 6, 2,
    -- layer=1 filter=153 channel=78
    -4, 8, 7, -10, -8, -7, 7, 0, 1,
    -- layer=1 filter=153 channel=79
    3, -6, -6, 8, -7, 0, -5, -11, -3,
    -- layer=1 filter=153 channel=80
    -6, 3, 7, 10, -5, -2, 0, 8, -2,
    -- layer=1 filter=153 channel=81
    6, -2, -3, -3, -5, 2, -3, -3, -6,
    -- layer=1 filter=153 channel=82
    -3, 8, 1, -9, -10, 7, -3, -4, 7,
    -- layer=1 filter=153 channel=83
    -7, -11, -1, 8, -5, 4, -9, 0, -1,
    -- layer=1 filter=153 channel=84
    -5, 2, 8, 3, -2, 0, -3, 0, -4,
    -- layer=1 filter=153 channel=85
    0, -1, -2, -1, 7, 4, 5, -10, 2,
    -- layer=1 filter=153 channel=86
    -6, -3, -7, -1, -4, -6, 4, 3, -6,
    -- layer=1 filter=153 channel=87
    3, 5, -3, 0, 5, -4, 8, 0, -11,
    -- layer=1 filter=153 channel=88
    -11, 2, 1, 7, -5, -12, -4, -11, 0,
    -- layer=1 filter=153 channel=89
    6, -1, -2, -8, -10, -1, 8, -9, 2,
    -- layer=1 filter=153 channel=90
    -9, 7, -7, -2, 8, 5, -3, -6, -8,
    -- layer=1 filter=153 channel=91
    4, 2, -1, -11, -8, -8, -6, 4, 6,
    -- layer=1 filter=153 channel=92
    1, -1, 8, 5, -7, -7, -6, 8, -7,
    -- layer=1 filter=153 channel=93
    5, 6, -11, -11, -6, 5, 1, 3, 1,
    -- layer=1 filter=153 channel=94
    -6, 4, 0, -2, 8, 6, -5, 6, -8,
    -- layer=1 filter=153 channel=95
    -10, 3, 0, -8, -9, 0, -8, 3, -7,
    -- layer=1 filter=153 channel=96
    4, 6, -4, -4, -1, -8, -4, -10, 0,
    -- layer=1 filter=153 channel=97
    2, -6, -11, 2, 7, 6, 3, 9, -10,
    -- layer=1 filter=153 channel=98
    -12, -1, 9, -7, -8, -3, -11, 4, 3,
    -- layer=1 filter=153 channel=99
    9, 8, 2, -1, -8, -3, -3, 5, 2,
    -- layer=1 filter=153 channel=100
    1, -7, 4, 0, 8, -4, 6, 4, 8,
    -- layer=1 filter=153 channel=101
    8, -6, -3, 4, 5, -11, 5, 0, 1,
    -- layer=1 filter=153 channel=102
    0, -7, -4, 5, -2, -2, 2, 8, 3,
    -- layer=1 filter=153 channel=103
    2, -7, 8, 0, 5, -2, 0, -7, -5,
    -- layer=1 filter=153 channel=104
    -1, -9, -10, -4, -5, -12, -8, 7, 3,
    -- layer=1 filter=153 channel=105
    -11, -3, -1, -2, 0, 0, -9, -9, -8,
    -- layer=1 filter=153 channel=106
    -9, -8, -8, -8, 5, -5, 8, 2, 8,
    -- layer=1 filter=153 channel=107
    -9, 0, 4, -7, -10, -2, -10, 7, -2,
    -- layer=1 filter=153 channel=108
    2, -8, 2, -1, -8, 1, -3, -11, -8,
    -- layer=1 filter=153 channel=109
    0, -6, -9, -7, 9, 1, 0, 2, 8,
    -- layer=1 filter=153 channel=110
    0, 8, -4, 8, -4, 2, 3, 3, -5,
    -- layer=1 filter=153 channel=111
    2, 3, -3, 7, 1, 3, -8, 11, 2,
    -- layer=1 filter=153 channel=112
    -8, 2, -3, 4, -6, 1, -9, -9, -8,
    -- layer=1 filter=153 channel=113
    -6, -1, 0, 2, -9, 0, -12, -9, 0,
    -- layer=1 filter=153 channel=114
    -2, -2, 0, -5, 0, 0, 1, -10, -5,
    -- layer=1 filter=153 channel=115
    0, 0, 1, 7, 3, -4, 1, 5, -10,
    -- layer=1 filter=153 channel=116
    -2, -1, -4, -3, -4, 5, 6, 9, 7,
    -- layer=1 filter=153 channel=117
    -10, 4, -11, -1, 6, -1, -3, 7, -2,
    -- layer=1 filter=153 channel=118
    8, -7, 5, -2, 0, 0, 0, -4, 5,
    -- layer=1 filter=153 channel=119
    -8, -3, -8, 7, 1, 2, 6, -5, 4,
    -- layer=1 filter=153 channel=120
    5, 4, -5, -4, 0, 4, -8, -8, 2,
    -- layer=1 filter=153 channel=121
    1, -2, -3, -7, 0, 5, 9, 5, -6,
    -- layer=1 filter=153 channel=122
    8, -9, 2, 7, 1, 0, -1, -2, -6,
    -- layer=1 filter=153 channel=123
    8, 8, -9, -4, -7, 8, 7, -6, -3,
    -- layer=1 filter=153 channel=124
    -6, 4, -6, 5, 12, 7, 2, -1, -3,
    -- layer=1 filter=153 channel=125
    -2, -4, 3, -3, 2, 2, -8, -8, -7,
    -- layer=1 filter=153 channel=126
    9, -4, 3, 8, -7, 1, 0, 0, 4,
    -- layer=1 filter=153 channel=127
    5, -7, -6, -10, -6, 4, 1, -9, 2,
    -- layer=1 filter=154 channel=0
    -25, -32, -26, -42, -50, -64, -23, -44, -49,
    -- layer=1 filter=154 channel=1
    -1, -12, -43, 0, -9, -5, -4, 0, 29,
    -- layer=1 filter=154 channel=2
    21, 33, 30, 36, 14, 13, 28, 29, 18,
    -- layer=1 filter=154 channel=3
    -9, 3, -3, 0, -2, -3, 0, 1, 6,
    -- layer=1 filter=154 channel=4
    -8, -24, -21, -8, -2, 4, -4, -10, -1,
    -- layer=1 filter=154 channel=5
    0, 4, -16, 25, 3, 0, 13, 24, 30,
    -- layer=1 filter=154 channel=6
    -10, -9, -33, 21, 32, -10, 21, 27, 3,
    -- layer=1 filter=154 channel=7
    -64, -38, 30, -29, -76, 26, -56, -34, 27,
    -- layer=1 filter=154 channel=8
    -4, 21, -22, 48, 17, 3, 3, 7, 18,
    -- layer=1 filter=154 channel=9
    8, 0, 22, -32, -11, -9, 16, 0, 40,
    -- layer=1 filter=154 channel=10
    -62, -72, 21, -28, -86, 3, -11, -21, 13,
    -- layer=1 filter=154 channel=11
    7, 13, 9, 10, -4, -4, 14, -2, -5,
    -- layer=1 filter=154 channel=12
    -2, 11, 6, 4, 13, -3, 46, 30, 42,
    -- layer=1 filter=154 channel=13
    8, 3, 8, 21, 48, 19, 9, 19, -11,
    -- layer=1 filter=154 channel=14
    -9, -39, 23, -40, -59, -10, 24, -35, -3,
    -- layer=1 filter=154 channel=15
    -8, 1, 7, 25, 52, 26, 34, 12, 26,
    -- layer=1 filter=154 channel=16
    10, 33, -8, 39, 29, 10, 23, 12, 6,
    -- layer=1 filter=154 channel=17
    0, 21, -5, 24, 35, 25, -8, 3, -11,
    -- layer=1 filter=154 channel=18
    29, 10, 25, 15, 22, 7, 36, 17, 9,
    -- layer=1 filter=154 channel=19
    23, 11, 7, 22, 29, 43, 33, -9, 1,
    -- layer=1 filter=154 channel=20
    1, 10, -18, 41, 29, 21, 29, 18, -4,
    -- layer=1 filter=154 channel=21
    -80, -46, -41, -28, -26, 0, 1, 8, 5,
    -- layer=1 filter=154 channel=22
    13, -1, -13, 44, 56, 35, 20, 27, 11,
    -- layer=1 filter=154 channel=23
    -28, -50, 16, -61, -79, 76, -72, -76, 67,
    -- layer=1 filter=154 channel=24
    -37, -19, -28, -29, -14, -34, -12, -1, 14,
    -- layer=1 filter=154 channel=25
    -42, -33, 24, 0, -29, 36, -7, -3, 51,
    -- layer=1 filter=154 channel=26
    3, 19, 12, 25, 43, 25, -11, 3, -13,
    -- layer=1 filter=154 channel=27
    25, 39, 12, 45, 45, 31, 40, 17, 29,
    -- layer=1 filter=154 channel=28
    -45, -26, 18, -32, -65, 12, -64, -61, 4,
    -- layer=1 filter=154 channel=29
    7, 7, 4, 40, 36, 27, 24, 1, 6,
    -- layer=1 filter=154 channel=30
    -12, -11, -6, -9, -2, -24, 40, 26, 22,
    -- layer=1 filter=154 channel=31
    42, 34, 25, 58, 66, 39, 70, 54, 34,
    -- layer=1 filter=154 channel=32
    -35, -4, -4, -42, -28, -12, -45, -33, -5,
    -- layer=1 filter=154 channel=33
    9, 0, -9, 11, 26, 2, 19, 14, -3,
    -- layer=1 filter=154 channel=34
    -17, -15, -28, 33, 38, -8, 18, 21, -18,
    -- layer=1 filter=154 channel=35
    -9, -18, -15, -21, -12, -20, 9, -9, -4,
    -- layer=1 filter=154 channel=36
    -2, 10, 9, -8, -25, -10, -4, -19, -22,
    -- layer=1 filter=154 channel=37
    -4, -7, -15, 22, 3, 9, 46, 26, 41,
    -- layer=1 filter=154 channel=38
    -11, -6, -37, 15, 20, 5, 6, 16, 5,
    -- layer=1 filter=154 channel=39
    14, 17, 2, -14, -8, -2, -25, -2, -12,
    -- layer=1 filter=154 channel=40
    37, 26, -1, 53, 69, 25, 67, 59, 6,
    -- layer=1 filter=154 channel=41
    -38, 4, 6, -77, -67, -23, -33, -35, 40,
    -- layer=1 filter=154 channel=42
    16, 37, 40, 42, 47, 60, 21, 30, 13,
    -- layer=1 filter=154 channel=43
    -6, 0, -7, 20, -2, 6, 7, 1, 14,
    -- layer=1 filter=154 channel=44
    -27, 2, 5, -18, -6, -1, -65, -48, -31,
    -- layer=1 filter=154 channel=45
    -56, -54, -64, -11, -5, -21, 5, 16, -14,
    -- layer=1 filter=154 channel=46
    -4, 7, -21, 27, 36, 15, 42, -6, 2,
    -- layer=1 filter=154 channel=47
    -30, -27, 42, -42, 8, 71, -8, 39, 68,
    -- layer=1 filter=154 channel=48
    -43, -44, -19, -49, -38, -32, -20, -20, -9,
    -- layer=1 filter=154 channel=49
    -23, -32, -17, 5, 10, -1, 33, 23, -4,
    -- layer=1 filter=154 channel=50
    17, -11, -1, 36, 43, 37, 10, 7, -3,
    -- layer=1 filter=154 channel=51
    -41, -57, -20, 6, -20, -9, 18, 10, 8,
    -- layer=1 filter=154 channel=52
    0, 17, 3, 11, 1, -12, -3, 11, 9,
    -- layer=1 filter=154 channel=53
    11, 10, 11, 13, 21, -3, 18, 20, 19,
    -- layer=1 filter=154 channel=54
    -30, -19, 28, 11, -2, 40, 14, 19, 29,
    -- layer=1 filter=154 channel=55
    29, 19, 24, 12, -4, -2, -9, -3, -1,
    -- layer=1 filter=154 channel=56
    0, -14, -1, -2, 11, -8, 3, 1, 2,
    -- layer=1 filter=154 channel=57
    11, -3, 22, 54, 27, 43, 45, 30, 40,
    -- layer=1 filter=154 channel=58
    -38, -79, 43, -76, -85, 62, -36, -34, 60,
    -- layer=1 filter=154 channel=59
    7, 5, -2, -15, -37, 4, -16, -14, -14,
    -- layer=1 filter=154 channel=60
    -29, -39, -38, 2, -18, 2, 8, -8, -4,
    -- layer=1 filter=154 channel=61
    -4, 13, 3, 3, 3, -1, -1, 3, -7,
    -- layer=1 filter=154 channel=62
    11, 8, -9, 14, 4, 0, 10, 1, 11,
    -- layer=1 filter=154 channel=63
    -4, 6, 0, -10, -16, -29, -12, -16, -30,
    -- layer=1 filter=154 channel=64
    -48, -34, -47, -22, -2, -22, -4, -9, -4,
    -- layer=1 filter=154 channel=65
    -42, -25, -40, -22, -32, -45, -19, -20, -46,
    -- layer=1 filter=154 channel=66
    -10, -5, -23, -37, -35, -43, -4, -11, -18,
    -- layer=1 filter=154 channel=67
    -21, -71, -90, -37, -34, -49, -3, -43, -39,
    -- layer=1 filter=154 channel=68
    -43, -13, -30, -55, -50, -29, -87, -61, -42,
    -- layer=1 filter=154 channel=69
    22, 14, -11, 24, 34, 2, 23, 17, 17,
    -- layer=1 filter=154 channel=70
    -9, -39, -48, 34, 29, -21, 52, 52, 2,
    -- layer=1 filter=154 channel=71
    -17, -12, -8, 1, -13, 6, -6, -34, -16,
    -- layer=1 filter=154 channel=72
    4, -2, -1, -5, 8, 3, 29, 18, 15,
    -- layer=1 filter=154 channel=73
    -10, -6, -11, 1, -3, 0, -8, -1, 4,
    -- layer=1 filter=154 channel=74
    -2, 4, -9, 9, 6, -8, 30, -10, 5,
    -- layer=1 filter=154 channel=75
    -9, 2, -1, -34, -12, -16, 26, 4, -5,
    -- layer=1 filter=154 channel=76
    -35, -38, -3, -50, -39, -40, -48, -80, -45,
    -- layer=1 filter=154 channel=77
    -56, -47, -39, -36, -31, -53, -6, 13, -1,
    -- layer=1 filter=154 channel=78
    2, 15, -17, 14, 4, 12, 11, 19, 20,
    -- layer=1 filter=154 channel=79
    12, 1, 7, 18, 23, 20, 11, 11, 7,
    -- layer=1 filter=154 channel=80
    -9, -10, -24, -18, -8, -4, -28, -13, -16,
    -- layer=1 filter=154 channel=81
    10, -16, 5, 2, -30, -8, 18, -11, 10,
    -- layer=1 filter=154 channel=82
    -76, -79, -59, -50, -52, -21, -23, -9, 4,
    -- layer=1 filter=154 channel=83
    -4, -24, -20, -27, -36, -33, -16, -4, 9,
    -- layer=1 filter=154 channel=84
    27, 40, 29, 26, 45, 35, 29, 16, -1,
    -- layer=1 filter=154 channel=85
    -7, -53, 49, -98, -73, 68, -38, -18, 27,
    -- layer=1 filter=154 channel=86
    53, 36, 39, 32, 29, 7, -9, 4, 9,
    -- layer=1 filter=154 channel=87
    34, 12, 27, 32, 48, 26, 72, 57, 43,
    -- layer=1 filter=154 channel=88
    -22, -32, -39, -31, -25, -33, 6, -2, -15,
    -- layer=1 filter=154 channel=89
    -57, -21, -47, -48, -32, -33, -8, 0, -33,
    -- layer=1 filter=154 channel=90
    -62, -27, -8, -74, -45, -38, -58, -41, -15,
    -- layer=1 filter=154 channel=91
    -16, -18, -23, 26, 22, 21, 25, 32, 20,
    -- layer=1 filter=154 channel=92
    -93, -19, -11, -66, -27, -15, -68, -58, 22,
    -- layer=1 filter=154 channel=93
    -64, -65, -32, -73, -84, -36, -32, -29, -6,
    -- layer=1 filter=154 channel=94
    -14, -5, -8, -6, 4, -22, -28, -29, -48,
    -- layer=1 filter=154 channel=95
    1, 2, 9, -9, -17, 0, 14, -6, -2,
    -- layer=1 filter=154 channel=96
    0, 6, -16, -20, -17, -31, -17, -12, -26,
    -- layer=1 filter=154 channel=97
    -15, -17, -8, -33, -29, -36, -41, -35, -34,
    -- layer=1 filter=154 channel=98
    -11, -30, -11, 19, -2, 5, 14, 8, 17,
    -- layer=1 filter=154 channel=99
    -55, -106, -47, -67, -124, -92, -52, -67, -36,
    -- layer=1 filter=154 channel=100
    -12, 6, 29, -13, 7, 0, 6, 13, 9,
    -- layer=1 filter=154 channel=101
    -24, -24, -33, 2, 13, -12, 7, 26, 4,
    -- layer=1 filter=154 channel=102
    -33, -19, -38, -12, 0, -35, -29, -35, -42,
    -- layer=1 filter=154 channel=103
    30, 20, 26, 11, 18, -2, 24, 22, 21,
    -- layer=1 filter=154 channel=104
    15, -15, 24, -5, -9, 50, -23, 12, 26,
    -- layer=1 filter=154 channel=105
    -7, -24, -4, -31, -43, -41, -40, -58, -29,
    -- layer=1 filter=154 channel=106
    -15, -16, -27, 0, 29, 3, 22, 20, 7,
    -- layer=1 filter=154 channel=107
    19, 0, -5, -11, -15, 1, -4, -6, 8,
    -- layer=1 filter=154 channel=108
    -41, -36, -23, -60, -44, -39, -48, -30, -11,
    -- layer=1 filter=154 channel=109
    3, -7, 6, -8, -7, 8, -3, -9, 0,
    -- layer=1 filter=154 channel=110
    -20, -11, -5, -15, -8, -15, -8, 2, -14,
    -- layer=1 filter=154 channel=111
    24, 0, 14, -10, -7, -33, 18, -12, -19,
    -- layer=1 filter=154 channel=112
    11, -14, 19, 27, 23, 16, 21, 17, 6,
    -- layer=1 filter=154 channel=113
    -9, -2, -5, 40, 36, 46, 60, 44, 8,
    -- layer=1 filter=154 channel=114
    62, 52, 19, 55, 31, 27, 21, 20, 26,
    -- layer=1 filter=154 channel=115
    23, 24, 24, 29, 10, 24, -10, -13, 11,
    -- layer=1 filter=154 channel=116
    1, -1, -5, 0, 4, 7, 8, -2, -10,
    -- layer=1 filter=154 channel=117
    33, 4, 10, 48, 23, 10, 36, 11, 7,
    -- layer=1 filter=154 channel=118
    5, 13, 15, 6, -4, -14, 9, 1, 13,
    -- layer=1 filter=154 channel=119
    -57, -42, -25, -88, -89, -76, -79, -69, -36,
    -- layer=1 filter=154 channel=120
    -63, -67, -19, -31, -30, 21, 0, 15, 34,
    -- layer=1 filter=154 channel=121
    26, 23, 8, 6, 13, 13, 22, -10, 4,
    -- layer=1 filter=154 channel=122
    9, -1, -1, 5, -2, -6, 9, -9, 2,
    -- layer=1 filter=154 channel=123
    0, 9, 14, 12, 2, 12, 31, -3, -1,
    -- layer=1 filter=154 channel=124
    6, 1, 6, -3, 8, 14, -2, 12, 11,
    -- layer=1 filter=154 channel=125
    -31, -41, -40, 16, 3, -3, 55, 53, 7,
    -- layer=1 filter=154 channel=126
    -24, -51, -40, 0, -23, -32, 6, 15, 31,
    -- layer=1 filter=154 channel=127
    8, 21, 5, 16, 18, 2, 29, 12, 30,
    -- layer=1 filter=155 channel=0
    3, -2, 1, -9, 6, 3, -11, -7, -8,
    -- layer=1 filter=155 channel=1
    -2, -13, 9, -2, 0, 4, 1, -17, -15,
    -- layer=1 filter=155 channel=2
    1, -13, -13, 0, -16, -3, 10, -2, 6,
    -- layer=1 filter=155 channel=3
    -3, -6, -6, 0, -7, -6, 8, 3, 5,
    -- layer=1 filter=155 channel=4
    -1, -1, 7, 2, -3, 7, -5, 0, 7,
    -- layer=1 filter=155 channel=5
    3, -2, -5, 3, -7, -10, -10, -9, -13,
    -- layer=1 filter=155 channel=6
    -8, -9, 0, -10, 5, -10, -7, -5, -8,
    -- layer=1 filter=155 channel=7
    6, -11, 0, 1, 8, -13, -12, 8, 5,
    -- layer=1 filter=155 channel=8
    -9, 11, 6, -8, -6, -5, -9, -7, -6,
    -- layer=1 filter=155 channel=9
    -3, -6, 3, -9, 0, -3, -3, -7, -12,
    -- layer=1 filter=155 channel=10
    -8, -18, -10, -10, -1, 9, -11, 7, -4,
    -- layer=1 filter=155 channel=11
    0, -7, -5, 6, 6, 7, 0, 0, 0,
    -- layer=1 filter=155 channel=12
    9, 5, -2, -4, -8, -4, 6, -8, 7,
    -- layer=1 filter=155 channel=13
    -6, -1, -16, -13, -9, 3, -13, -8, 1,
    -- layer=1 filter=155 channel=14
    -7, 2, -9, -7, 13, 0, -7, 0, 15,
    -- layer=1 filter=155 channel=15
    0, -5, -9, 5, 1, 5, 0, -3, -1,
    -- layer=1 filter=155 channel=16
    7, 0, 3, -1, -10, -11, -14, -13, 4,
    -- layer=1 filter=155 channel=17
    -6, -6, 4, -8, -12, -10, 4, -10, -14,
    -- layer=1 filter=155 channel=18
    1, -8, 4, 3, -2, 3, -3, 3, -6,
    -- layer=1 filter=155 channel=19
    -12, -13, -11, 2, 0, 3, 4, 9, -11,
    -- layer=1 filter=155 channel=20
    5, -6, -3, -5, -8, -6, -3, 1, -14,
    -- layer=1 filter=155 channel=21
    -3, 1, -12, 3, -5, 0, -15, -12, -6,
    -- layer=1 filter=155 channel=22
    0, 0, -2, -8, -3, -5, -3, -14, 8,
    -- layer=1 filter=155 channel=23
    7, -15, 8, 1, 0, -7, -2, -11, -4,
    -- layer=1 filter=155 channel=24
    2, -14, -2, -13, -15, 1, -15, -14, -13,
    -- layer=1 filter=155 channel=25
    -5, 6, 1, 2, -8, 0, -15, -3, 1,
    -- layer=1 filter=155 channel=26
    0, 3, 3, -5, -3, -12, 6, -9, 1,
    -- layer=1 filter=155 channel=27
    6, -4, 0, -9, 1, -6, 10, 0, -6,
    -- layer=1 filter=155 channel=28
    -6, -14, -4, 4, 0, -6, -8, 0, 5,
    -- layer=1 filter=155 channel=29
    5, -11, 7, -9, -2, 7, -5, 0, -5,
    -- layer=1 filter=155 channel=30
    -2, -2, 4, 6, 6, 3, 2, 0, 6,
    -- layer=1 filter=155 channel=31
    -8, -12, -8, -8, 0, 3, 1, -7, 0,
    -- layer=1 filter=155 channel=32
    -9, -17, 6, -4, -6, -7, 6, -1, -8,
    -- layer=1 filter=155 channel=33
    4, 4, 3, -3, -16, -10, -4, 6, 0,
    -- layer=1 filter=155 channel=34
    6, 8, 0, -2, -7, -6, 6, 3, -6,
    -- layer=1 filter=155 channel=35
    2, 6, 0, 3, 4, -4, -9, -8, 3,
    -- layer=1 filter=155 channel=36
    0, -1, -7, 6, 7, -6, -14, 4, -6,
    -- layer=1 filter=155 channel=37
    9, 10, -2, 0, 0, 4, -17, -12, -7,
    -- layer=1 filter=155 channel=38
    -13, -11, 2, -9, -7, -1, -4, 6, 7,
    -- layer=1 filter=155 channel=39
    8, -1, -8, 4, -4, 3, -2, -8, -1,
    -- layer=1 filter=155 channel=40
    0, -2, -4, 8, 8, -2, 7, 9, -7,
    -- layer=1 filter=155 channel=41
    -8, -7, 6, -3, 9, -4, 0, 0, -7,
    -- layer=1 filter=155 channel=42
    -11, -1, -12, -13, -3, -1, 2, 5, -5,
    -- layer=1 filter=155 channel=43
    2, -10, 1, -5, -16, -6, -6, -10, -2,
    -- layer=1 filter=155 channel=44
    -13, 0, 7, 0, -14, 4, -4, 2, 2,
    -- layer=1 filter=155 channel=45
    -6, -7, -6, -1, -9, 3, 2, -11, 0,
    -- layer=1 filter=155 channel=46
    -14, 9, -2, -13, -2, -8, -16, -9, -19,
    -- layer=1 filter=155 channel=47
    9, -9, -8, 5, -6, -2, 7, 7, -11,
    -- layer=1 filter=155 channel=48
    5, -11, 2, -12, -2, 0, -13, -3, -4,
    -- layer=1 filter=155 channel=49
    -4, -8, -3, 4, -8, -14, -1, -4, -6,
    -- layer=1 filter=155 channel=50
    -9, -13, -6, -8, -10, -1, -8, 5, -7,
    -- layer=1 filter=155 channel=51
    -11, 2, 3, 5, 1, -11, -5, -1, 5,
    -- layer=1 filter=155 channel=52
    2, -7, -9, 0, -4, 11, -8, 9, 8,
    -- layer=1 filter=155 channel=53
    -9, -2, 5, 5, -12, -8, 8, -4, -3,
    -- layer=1 filter=155 channel=54
    6, -1, 8, -19, 7, 0, 0, 0, -1,
    -- layer=1 filter=155 channel=55
    2, -9, 10, 6, 7, -11, -4, -6, -8,
    -- layer=1 filter=155 channel=56
    0, 6, 4, 4, -4, -1, 4, -7, -7,
    -- layer=1 filter=155 channel=57
    6, 2, 7, -9, -5, -8, -9, -9, 1,
    -- layer=1 filter=155 channel=58
    -3, -2, -12, -13, 0, -5, 2, 0, 5,
    -- layer=1 filter=155 channel=59
    -8, -6, -10, -11, -8, -7, -4, -10, 3,
    -- layer=1 filter=155 channel=60
    1, -10, -8, -4, -6, -4, 6, -4, -8,
    -- layer=1 filter=155 channel=61
    1, -9, 4, 0, 10, 6, -8, -2, 2,
    -- layer=1 filter=155 channel=62
    12, 4, 6, -4, -11, 9, 0, 3, -10,
    -- layer=1 filter=155 channel=63
    -9, -2, 3, 1, -9, -3, -10, -5, 0,
    -- layer=1 filter=155 channel=64
    -6, -7, 0, -13, -10, -15, -8, 2, 5,
    -- layer=1 filter=155 channel=65
    -2, -10, -2, -9, -6, -9, 4, -8, -10,
    -- layer=1 filter=155 channel=66
    1, 7, -4, 6, 0, -8, 1, 2, -14,
    -- layer=1 filter=155 channel=67
    -11, -5, -7, -6, 10, 6, -2, 1, 1,
    -- layer=1 filter=155 channel=68
    -11, 2, -10, 2, 4, 2, -8, -3, 3,
    -- layer=1 filter=155 channel=69
    0, 8, -6, 0, -15, -2, 0, 2, -11,
    -- layer=1 filter=155 channel=70
    -5, -10, -9, -4, 0, -11, 3, 0, 0,
    -- layer=1 filter=155 channel=71
    -3, 0, -7, -4, 7, -4, -11, -10, -8,
    -- layer=1 filter=155 channel=72
    4, -1, 6, 0, -9, -9, 6, 4, -1,
    -- layer=1 filter=155 channel=73
    -6, 7, 7, -2, 0, 1, -3, -2, 6,
    -- layer=1 filter=155 channel=74
    1, 4, 1, -4, -12, -11, 8, -9, -3,
    -- layer=1 filter=155 channel=75
    6, -11, 3, 22, 5, 12, 0, -3, 1,
    -- layer=1 filter=155 channel=76
    -6, -7, -11, 5, -11, -2, 2, 8, -4,
    -- layer=1 filter=155 channel=77
    5, -7, -10, -16, -5, -3, -10, -5, -7,
    -- layer=1 filter=155 channel=78
    0, -5, -2, -10, -7, -6, 0, -4, 1,
    -- layer=1 filter=155 channel=79
    -10, 0, 6, -10, -4, -6, 0, -7, 4,
    -- layer=1 filter=155 channel=80
    -2, 2, 0, -4, 3, -2, -10, -9, 0,
    -- layer=1 filter=155 channel=81
    -11, -8, -2, 0, -11, -13, -2, 0, 1,
    -- layer=1 filter=155 channel=82
    -10, 2, -11, -2, -10, -14, 1, -1, -6,
    -- layer=1 filter=155 channel=83
    -10, -8, 6, 5, -5, 0, -8, -14, 0,
    -- layer=1 filter=155 channel=84
    2, -18, -5, -4, 0, 10, 7, 5, 5,
    -- layer=1 filter=155 channel=85
    7, -6, -4, -4, -11, -4, -7, 0, 3,
    -- layer=1 filter=155 channel=86
    -1, 5, -5, 0, -5, 0, -13, 0, -4,
    -- layer=1 filter=155 channel=87
    7, -2, -3, 1, 9, 4, 2, 3, -3,
    -- layer=1 filter=155 channel=88
    -14, 2, 0, -12, -10, 0, -10, 5, -4,
    -- layer=1 filter=155 channel=89
    -9, -7, -3, 5, 4, -3, -6, -12, -12,
    -- layer=1 filter=155 channel=90
    -17, -17, -2, 2, -8, -4, -3, -10, 6,
    -- layer=1 filter=155 channel=91
    4, 7, -1, -4, 3, 5, 1, -9, -5,
    -- layer=1 filter=155 channel=92
    0, 4, 13, -5, 6, -11, -6, 0, 7,
    -- layer=1 filter=155 channel=93
    -1, -13, 4, -8, -13, -17, -2, 3, -11,
    -- layer=1 filter=155 channel=94
    -10, 0, -2, 0, 0, -9, -8, 5, 0,
    -- layer=1 filter=155 channel=95
    -11, -4, 3, 6, 4, -4, -8, -5, 1,
    -- layer=1 filter=155 channel=96
    5, -7, -8, 6, 0, -10, 0, 1, -10,
    -- layer=1 filter=155 channel=97
    -10, 3, -6, 2, 0, -6, 0, -15, 4,
    -- layer=1 filter=155 channel=98
    -1, 1, 9, -11, -10, -9, -5, -6, -5,
    -- layer=1 filter=155 channel=99
    4, 10, -3, -7, -2, -11, -5, -14, -5,
    -- layer=1 filter=155 channel=100
    -11, -8, 6, -3, 4, 1, -2, -12, -12,
    -- layer=1 filter=155 channel=101
    -4, -5, -10, 4, -9, -9, -8, 0, 4,
    -- layer=1 filter=155 channel=102
    -13, 2, -6, 3, -8, 0, 2, 0, 0,
    -- layer=1 filter=155 channel=103
    0, 9, -7, 7, -7, -3, 1, 3, 6,
    -- layer=1 filter=155 channel=104
    -7, -7, 4, -11, 7, 5, -9, -1, -6,
    -- layer=1 filter=155 channel=105
    -10, 1, 0, -2, -4, -6, -14, 4, 0,
    -- layer=1 filter=155 channel=106
    -10, -9, 0, -11, -6, -14, -14, 5, -3,
    -- layer=1 filter=155 channel=107
    9, 0, -1, 6, -9, 6, -4, 2, 12,
    -- layer=1 filter=155 channel=108
    -12, -12, 9, 2, -5, 4, 3, 0, 3,
    -- layer=1 filter=155 channel=109
    -7, -7, -3, -2, -4, 2, 3, -5, 9,
    -- layer=1 filter=155 channel=110
    -9, -7, 4, 5, 0, 0, -6, -5, -12,
    -- layer=1 filter=155 channel=111
    -5, -10, -8, -7, -1, -7, 3, 15, 3,
    -- layer=1 filter=155 channel=112
    -3, 8, -3, 0, 5, 0, -7, -4, 2,
    -- layer=1 filter=155 channel=113
    -10, -7, 6, 0, 0, -1, -4, -1, 3,
    -- layer=1 filter=155 channel=114
    -6, 5, 13, -3, -2, -15, -16, -12, -6,
    -- layer=1 filter=155 channel=115
    8, -11, -9, 2, -9, -13, -5, -9, -12,
    -- layer=1 filter=155 channel=116
    -7, -3, -9, 4, 11, 8, 4, 6, -1,
    -- layer=1 filter=155 channel=117
    -1, -3, 2, 1, 1, -7, 8, 6, -8,
    -- layer=1 filter=155 channel=118
    -13, -13, -9, 7, -12, 1, -3, -6, 0,
    -- layer=1 filter=155 channel=119
    -18, -6, -3, -2, -6, 5, -8, -7, -6,
    -- layer=1 filter=155 channel=120
    6, 1, 0, -6, -14, -1, 3, 2, -6,
    -- layer=1 filter=155 channel=121
    -3, -8, -8, -5, -8, 7, -8, 7, -8,
    -- layer=1 filter=155 channel=122
    0, -2, -5, -10, -3, 2, -4, 3, 0,
    -- layer=1 filter=155 channel=123
    4, -7, -7, -9, -4, 8, 2, -14, -9,
    -- layer=1 filter=155 channel=124
    0, -9, 1, 5, -10, 4, -2, 6, -11,
    -- layer=1 filter=155 channel=125
    -6, 6, -9, -17, 2, -7, 0, -5, -14,
    -- layer=1 filter=155 channel=126
    4, -5, 12, -4, 4, -11, -9, -16, 2,
    -- layer=1 filter=155 channel=127
    -4, -7, -8, 4, 5, 4, 0, -13, 3,
    -- layer=1 filter=156 channel=0
    -11, 12, 17, 8, 19, 13, 14, 23, 9,
    -- layer=1 filter=156 channel=1
    -11, -1, -17, -15, -8, 1, 13, 17, -13,
    -- layer=1 filter=156 channel=2
    3, -37, -23, 34, 20, 5, -8, 16, 29,
    -- layer=1 filter=156 channel=3
    1, 6, -8, -9, -6, 6, 6, 2, 1,
    -- layer=1 filter=156 channel=4
    -9, -6, 2, 6, -1, -4, 5, -1, 0,
    -- layer=1 filter=156 channel=5
    -19, 14, 0, -28, -26, -9, 21, 17, -21,
    -- layer=1 filter=156 channel=6
    23, 13, -8, -14, 6, 15, -34, -37, -35,
    -- layer=1 filter=156 channel=7
    49, 36, 10, 17, 17, 0, -2, -33, -4,
    -- layer=1 filter=156 channel=8
    -13, -6, -20, -16, -3, 8, 20, -1, -24,
    -- layer=1 filter=156 channel=9
    -9, 6, -23, -19, -10, 16, 20, -10, -47,
    -- layer=1 filter=156 channel=10
    53, 35, 19, 3, 7, 0, 14, -32, -7,
    -- layer=1 filter=156 channel=11
    -39, -18, 5, -6, -14, 11, -15, -24, -27,
    -- layer=1 filter=156 channel=12
    53, 14, 13, 9, 54, 60, -10, -27, 34,
    -- layer=1 filter=156 channel=13
    -46, -17, -23, -62, -46, -22, -28, -42, -16,
    -- layer=1 filter=156 channel=14
    43, 45, -8, 22, 27, 22, -1, -33, -13,
    -- layer=1 filter=156 channel=15
    -14, 4, -15, 4, -25, -21, 45, 41, 24,
    -- layer=1 filter=156 channel=16
    -1, -9, -32, -12, 0, 0, 26, 23, -5,
    -- layer=1 filter=156 channel=17
    -17, -10, 5, -30, -3, -9, -31, -11, 3,
    -- layer=1 filter=156 channel=18
    -21, -1, -6, -11, 37, 41, 4, -52, -41,
    -- layer=1 filter=156 channel=19
    8, -8, -35, -26, -16, -19, 7, -4, 9,
    -- layer=1 filter=156 channel=20
    -47, -10, -15, -55, -52, -3, -23, -26, -10,
    -- layer=1 filter=156 channel=21
    7, 1, -12, -9, -4, 1, 14, 0, -3,
    -- layer=1 filter=156 channel=22
    -10, -16, -12, -31, -25, 0, -4, -2, -9,
    -- layer=1 filter=156 channel=23
    46, 5, -9, 22, -15, -25, 2, 7, -30,
    -- layer=1 filter=156 channel=24
    -22, -45, -34, -17, -33, -1, 12, 1, 6,
    -- layer=1 filter=156 channel=25
    35, 41, 7, -3, -19, -12, 29, -14, -32,
    -- layer=1 filter=156 channel=26
    -36, -75, -24, -63, -62, -1, -20, -19, -17,
    -- layer=1 filter=156 channel=27
    -18, -26, -11, -24, -15, -36, -12, -31, -36,
    -- layer=1 filter=156 channel=28
    40, 26, -5, 4, 12, -4, 12, -12, -19,
    -- layer=1 filter=156 channel=29
    -31, -11, -7, -7, -8, -10, -9, -24, -25,
    -- layer=1 filter=156 channel=30
    1, 21, -7, -27, 12, 34, 13, -51, -9,
    -- layer=1 filter=156 channel=31
    19, 19, -17, -5, 32, 27, -1, 5, -2,
    -- layer=1 filter=156 channel=32
    -10, -28, -8, -32, -18, -20, -7, -22, -5,
    -- layer=1 filter=156 channel=33
    0, -11, -17, 0, 0, -7, 7, 9, -9,
    -- layer=1 filter=156 channel=34
    15, -2, 4, 2, 1, -9, -3, 5, -10,
    -- layer=1 filter=156 channel=35
    -10, -6, -8, -6, -2, 7, -2, -7, 0,
    -- layer=1 filter=156 channel=36
    -31, -17, 8, -17, 6, 1, -6, -18, -23,
    -- layer=1 filter=156 channel=37
    -6, 11, -24, 3, -13, -12, 18, 17, -16,
    -- layer=1 filter=156 channel=38
    -33, 7, -12, -50, -21, -13, -50, -27, -11,
    -- layer=1 filter=156 channel=39
    -7, 5, 13, -3, 2, 23, 5, 6, 0,
    -- layer=1 filter=156 channel=40
    12, 9, -23, -21, 5, 19, -29, -32, -12,
    -- layer=1 filter=156 channel=41
    5, -23, -43, -27, -3, -11, 19, -34, -21,
    -- layer=1 filter=156 channel=42
    30, -24, -25, 42, 24, -2, 0, 17, 24,
    -- layer=1 filter=156 channel=43
    24, 10, -8, -16, -3, -12, 20, 10, -11,
    -- layer=1 filter=156 channel=44
    -18, -41, -18, -14, -16, 3, 4, -16, 8,
    -- layer=1 filter=156 channel=45
    -32, 9, -40, -33, -16, -18, 8, 0, -11,
    -- layer=1 filter=156 channel=46
    15, -22, -34, 5, -12, -12, 2, 25, 18,
    -- layer=1 filter=156 channel=47
    19, -18, -3, 14, -41, -36, -14, -22, -31,
    -- layer=1 filter=156 channel=48
    30, 28, 15, -15, 6, 17, -14, -25, -8,
    -- layer=1 filter=156 channel=49
    0, -25, -26, 9, -14, -33, -3, -5, -11,
    -- layer=1 filter=156 channel=50
    -9, -5, 6, -7, 3, -8, 9, 1, -7,
    -- layer=1 filter=156 channel=51
    16, 9, -5, 3, 6, 1, -8, -39, -12,
    -- layer=1 filter=156 channel=52
    21, -30, -11, 25, 8, -17, -22, 0, -1,
    -- layer=1 filter=156 channel=53
    0, 1, 6, 5, 11, -2, -7, -5, 3,
    -- layer=1 filter=156 channel=54
    29, 37, -14, 12, -23, -22, 41, -24, -33,
    -- layer=1 filter=156 channel=55
    -26, -27, -18, -9, -27, -26, 5, -4, -41,
    -- layer=1 filter=156 channel=56
    1, 0, 0, -1, 1, 0, 0, -10, -2,
    -- layer=1 filter=156 channel=57
    44, 12, 5, 1, -8, -3, 13, -22, -35,
    -- layer=1 filter=156 channel=58
    56, 16, 8, -4, -32, -8, 23, -16, -39,
    -- layer=1 filter=156 channel=59
    -10, 3, 3, -9, -8, 0, -5, -4, 0,
    -- layer=1 filter=156 channel=60
    0, 5, 27, -1, 13, 14, -6, 33, 3,
    -- layer=1 filter=156 channel=61
    -3, -3, -2, -3, -5, -7, -3, -9, -2,
    -- layer=1 filter=156 channel=62
    -11, -4, -37, -24, 1, 0, 11, 20, -29,
    -- layer=1 filter=156 channel=63
    -30, 0, 11, -24, 3, 16, -14, -40, -41,
    -- layer=1 filter=156 channel=64
    13, 25, 34, -4, 0, -10, -9, 0, 5,
    -- layer=1 filter=156 channel=65
    12, 33, 5, -26, -15, 5, -27, -3, -17,
    -- layer=1 filter=156 channel=66
    -3, 4, 14, 6, 7, -4, -1, -17, -8,
    -- layer=1 filter=156 channel=67
    12, -17, -4, -16, -3, 2, 14, 6, -9,
    -- layer=1 filter=156 channel=68
    -40, -45, -27, -49, -40, -15, -18, -25, 10,
    -- layer=1 filter=156 channel=69
    -21, 0, -53, -35, -45, -31, 19, 9, -15,
    -- layer=1 filter=156 channel=70
    22, 15, 16, -1, 5, 7, 9, -22, 25,
    -- layer=1 filter=156 channel=71
    3, -6, -27, 0, -2, 0, -5, 9, -6,
    -- layer=1 filter=156 channel=72
    14, -6, -10, -22, 6, 17, 3, -12, -8,
    -- layer=1 filter=156 channel=73
    -1, 0, 5, -7, -7, -1, 7, 7, 6,
    -- layer=1 filter=156 channel=74
    5, -6, 13, 0, 19, 29, 8, -19, -5,
    -- layer=1 filter=156 channel=75
    13, -4, -29, 12, 26, 29, -43, -41, -2,
    -- layer=1 filter=156 channel=76
    -13, -9, 30, -25, -6, 32, -5, -21, -14,
    -- layer=1 filter=156 channel=77
    -25, 1, -1, -11, 4, 9, 3, -17, 0,
    -- layer=1 filter=156 channel=78
    2, 10, 29, 0, -4, 12, 30, -25, 19,
    -- layer=1 filter=156 channel=79
    0, -16, -37, -15, -15, -4, 21, 15, -17,
    -- layer=1 filter=156 channel=80
    14, 6, 24, 6, -8, -1, -9, -1, -10,
    -- layer=1 filter=156 channel=81
    -10, -12, 3, -19, -2, -13, 15, -4, -24,
    -- layer=1 filter=156 channel=82
    -7, 11, 20, -25, -7, 8, -31, -23, -9,
    -- layer=1 filter=156 channel=83
    -8, 9, -22, 0, -9, -16, 10, -7, -23,
    -- layer=1 filter=156 channel=84
    -28, -11, -6, -28, 24, 42, -3, -35, -37,
    -- layer=1 filter=156 channel=85
    45, -9, 0, 3, -11, -39, 8, -9, -26,
    -- layer=1 filter=156 channel=86
    -20, 2, -4, -13, 1, -21, 16, -12, -24,
    -- layer=1 filter=156 channel=87
    -5, -11, -30, -20, -27, -17, 20, -1, 31,
    -- layer=1 filter=156 channel=88
    18, 2, 10, 42, 20, 11, 22, 3, 4,
    -- layer=1 filter=156 channel=89
    -16, -2, 2, -7, -5, -3, -38, -16, 1,
    -- layer=1 filter=156 channel=90
    -16, -23, -8, -18, -50, 11, 3, -9, 6,
    -- layer=1 filter=156 channel=91
    7, 6, 18, -22, -10, 3, -27, -35, -34,
    -- layer=1 filter=156 channel=92
    -24, -15, -35, 0, -30, 3, 7, -5, 12,
    -- layer=1 filter=156 channel=93
    -8, -6, 2, -22, -8, -18, -7, 3, -8,
    -- layer=1 filter=156 channel=94
    -9, 4, 16, 0, 12, -2, 17, -1, -9,
    -- layer=1 filter=156 channel=95
    -22, 11, 1, -22, 27, 30, -2, -37, -44,
    -- layer=1 filter=156 channel=96
    -14, -9, -9, -4, -7, -16, 3, 0, 16,
    -- layer=1 filter=156 channel=97
    -28, -2, -5, -12, -16, -5, 4, -8, -5,
    -- layer=1 filter=156 channel=98
    -10, 4, -23, -14, 13, -1, 0, 10, -28,
    -- layer=1 filter=156 channel=99
    24, 4, -5, 26, 16, -1, -13, -11, -12,
    -- layer=1 filter=156 channel=100
    0, 1, 3, -27, 10, -1, 0, -24, -37,
    -- layer=1 filter=156 channel=101
    -7, 2, -5, -27, -4, -10, -67, -29, -7,
    -- layer=1 filter=156 channel=102
    -9, 10, 17, -1, 24, 1, -15, 0, -4,
    -- layer=1 filter=156 channel=103
    -27, -10, -19, -12, -26, 11, -22, -22, -42,
    -- layer=1 filter=156 channel=104
    19, 4, -7, 8, -18, -29, -3, 6, -23,
    -- layer=1 filter=156 channel=105
    -3, 4, -1, -5, -3, 4, -10, -5, -18,
    -- layer=1 filter=156 channel=106
    -44, -10, 5, -57, -41, -11, -41, -32, -7,
    -- layer=1 filter=156 channel=107
    -6, -11, 7, -3, 7, 0, 1, -3, -2,
    -- layer=1 filter=156 channel=108
    -11, -59, 9, -35, -48, -3, -11, -1, -11,
    -- layer=1 filter=156 channel=109
    10, -5, 7, -7, -5, 4, -8, 9, 1,
    -- layer=1 filter=156 channel=110
    4, -9, -16, -14, -9, -1, 10, 0, -11,
    -- layer=1 filter=156 channel=111
    -8, 9, -2, -17, 29, 29, 7, -57, -43,
    -- layer=1 filter=156 channel=112
    -19, -4, 0, -6, 37, 26, -37, -47, -3,
    -- layer=1 filter=156 channel=113
    42, -36, -6, 23, 0, -3, 30, 11, 13,
    -- layer=1 filter=156 channel=114
    6, 0, -30, -30, -16, -2, 9, 18, -20,
    -- layer=1 filter=156 channel=115
    13, 5, -9, 4, 5, -2, 13, -19, -24,
    -- layer=1 filter=156 channel=116
    -2, 5, -2, 9, -9, -1, 8, -6, 7,
    -- layer=1 filter=156 channel=117
    -15, 0, 0, -27, 27, 31, -19, -28, -31,
    -- layer=1 filter=156 channel=118
    -23, 1, -7, -31, 8, 19, -6, -37, -38,
    -- layer=1 filter=156 channel=119
    -6, -57, -14, -50, -35, -4, -8, -22, 0,
    -- layer=1 filter=156 channel=120
    31, 27, -4, -12, -32, -28, 8, -30, -55,
    -- layer=1 filter=156 channel=121
    0, 13, -30, -8, 16, 20, -50, -4, 29,
    -- layer=1 filter=156 channel=122
    9, -10, 6, -1, -5, 7, -8, -5, -3,
    -- layer=1 filter=156 channel=123
    1, -3, -22, -28, 5, -2, -22, -5, -17,
    -- layer=1 filter=156 channel=124
    6, -1, 3, 0, 8, -12, 1, 5, 2,
    -- layer=1 filter=156 channel=125
    29, 11, 14, 47, 8, 13, 2, -22, 7,
    -- layer=1 filter=156 channel=126
    -3, -8, -21, 1, 0, 9, 1, -4, -8,
    -- layer=1 filter=156 channel=127
    2, 0, -6, -23, 34, 33, 0, -45, -23,
    -- layer=1 filter=157 channel=0
    0, 2, 3, -2, -11, -6, -18, -12, -10,
    -- layer=1 filter=157 channel=1
    -1, 5, 2, -14, -12, -6, -15, -12, -10,
    -- layer=1 filter=157 channel=2
    0, -8, -15, 3, -8, -6, -3, 0, 1,
    -- layer=1 filter=157 channel=3
    -3, -6, -3, 4, 1, 6, -8, 9, 6,
    -- layer=1 filter=157 channel=4
    1, 4, -11, 8, 7, 8, -3, -4, 4,
    -- layer=1 filter=157 channel=5
    -1, 4, -8, 2, 4, -9, -7, -20, -9,
    -- layer=1 filter=157 channel=6
    -20, -5, 2, 7, 10, -3, 10, -3, 10,
    -- layer=1 filter=157 channel=7
    -6, 9, 0, 5, -11, -4, -1, -16, -19,
    -- layer=1 filter=157 channel=8
    -2, 8, 2, -12, -5, -4, 4, -7, 1,
    -- layer=1 filter=157 channel=9
    -6, 2, -18, -18, -9, 7, 2, 9, -8,
    -- layer=1 filter=157 channel=10
    -5, 3, 4, 0, -3, -7, -8, -4, -2,
    -- layer=1 filter=157 channel=11
    -14, -1, 8, 5, -9, -3, -2, -9, -3,
    -- layer=1 filter=157 channel=12
    -8, -7, 16, 0, -8, -16, -12, 6, -2,
    -- layer=1 filter=157 channel=13
    -6, -10, -10, -13, -3, 4, -13, 3, -5,
    -- layer=1 filter=157 channel=14
    -4, 9, 3, 15, -23, 7, -6, 5, 10,
    -- layer=1 filter=157 channel=15
    -8, 9, 7, -12, 4, 2, -7, 6, -12,
    -- layer=1 filter=157 channel=16
    6, -2, 2, -13, -6, 2, -15, -15, -16,
    -- layer=1 filter=157 channel=17
    -7, 3, 3, -17, -19, -6, -8, -9, -10,
    -- layer=1 filter=157 channel=18
    -3, -3, -1, 5, 1, 5, -6, -2, 11,
    -- layer=1 filter=157 channel=19
    5, 5, -1, -11, 4, -10, -4, -7, -9,
    -- layer=1 filter=157 channel=20
    -14, 2, -8, -2, -4, -5, 0, -8, -8,
    -- layer=1 filter=157 channel=21
    -18, -9, 1, -8, -13, -22, 0, -9, -17,
    -- layer=1 filter=157 channel=22
    -8, -7, -11, -16, -16, -7, -3, -1, -3,
    -- layer=1 filter=157 channel=23
    4, -4, -10, 4, -1, -8, -9, 2, 0,
    -- layer=1 filter=157 channel=24
    -2, -22, -2, -6, -2, -3, -7, 8, -12,
    -- layer=1 filter=157 channel=25
    3, -6, -5, -16, 3, -13, 0, -4, -20,
    -- layer=1 filter=157 channel=26
    -7, -4, -4, -26, 5, 15, -5, -9, 6,
    -- layer=1 filter=157 channel=27
    -7, 8, 7, -7, 6, -5, -4, 10, -10,
    -- layer=1 filter=157 channel=28
    -8, -11, 1, -10, 6, 4, -12, -7, -6,
    -- layer=1 filter=157 channel=29
    -9, -6, -15, -8, -6, -12, -14, 3, 3,
    -- layer=1 filter=157 channel=30
    6, -10, 4, 7, 3, 3, 0, 0, 3,
    -- layer=1 filter=157 channel=31
    7, 4, 3, 3, 9, 8, 0, 0, 15,
    -- layer=1 filter=157 channel=32
    -1, -18, -7, -29, -4, 18, -9, 2, -5,
    -- layer=1 filter=157 channel=33
    -1, 5, 7, 4, 3, 15, 11, -3, 5,
    -- layer=1 filter=157 channel=34
    -11, -6, 8, -1, 1, -11, -1, -3, 9,
    -- layer=1 filter=157 channel=35
    3, -10, -3, -8, -11, 3, 1, -6, -2,
    -- layer=1 filter=157 channel=36
    2, -2, -3, -3, -3, 0, -7, -9, -13,
    -- layer=1 filter=157 channel=37
    14, -3, 5, -2, -3, -20, -22, -14, -12,
    -- layer=1 filter=157 channel=38
    -14, -24, -23, -3, 6, 0, -17, -5, 0,
    -- layer=1 filter=157 channel=39
    -7, 2, -2, -9, 0, 1, -11, -6, -3,
    -- layer=1 filter=157 channel=40
    2, 0, 5, 9, 3, 11, 9, 9, 7,
    -- layer=1 filter=157 channel=41
    7, -11, -7, -12, 3, -1, -10, -9, -8,
    -- layer=1 filter=157 channel=42
    -11, -8, -10, 4, -18, -13, -2, -11, 2,
    -- layer=1 filter=157 channel=43
    7, 0, -7, -1, 4, -9, -10, -12, -7,
    -- layer=1 filter=157 channel=44
    -3, -14, -1, -10, 8, 0, -12, 1, -4,
    -- layer=1 filter=157 channel=45
    -1, -5, -3, -1, -4, -3, -13, -9, -5,
    -- layer=1 filter=157 channel=46
    4, -8, 1, -5, 1, 1, -5, -14, -14,
    -- layer=1 filter=157 channel=47
    -6, 0, -12, 0, -5, -11, -1, 0, -10,
    -- layer=1 filter=157 channel=48
    -9, -5, -15, -8, -9, -3, -13, 5, -3,
    -- layer=1 filter=157 channel=49
    -13, 0, -11, -2, -16, -7, -8, 10, -9,
    -- layer=1 filter=157 channel=50
    5, -7, 3, -10, 4, -9, 6, -3, 0,
    -- layer=1 filter=157 channel=51
    -14, 2, -7, 1, -1, -17, -3, 0, -1,
    -- layer=1 filter=157 channel=52
    -6, 5, 2, -3, -2, 7, 4, 3, 3,
    -- layer=1 filter=157 channel=53
    4, 2, -2, -9, -8, 1, -7, -6, -11,
    -- layer=1 filter=157 channel=54
    -9, -14, -10, -14, 0, -14, -21, 1, -8,
    -- layer=1 filter=157 channel=55
    -13, -14, 0, 0, -9, -2, 7, -14, -10,
    -- layer=1 filter=157 channel=56
    -6, 4, 8, 2, 0, -1, 8, 5, -11,
    -- layer=1 filter=157 channel=57
    7, -3, -5, -6, -6, 1, 0, -11, -6,
    -- layer=1 filter=157 channel=58
    -5, -10, -11, -11, -5, -3, -16, -16, -15,
    -- layer=1 filter=157 channel=59
    1, 3, -5, -4, -4, -2, 5, 8, 0,
    -- layer=1 filter=157 channel=60
    2, -1, 11, -1, -3, 10, -2, -5, -4,
    -- layer=1 filter=157 channel=61
    -10, 1, 0, 6, 8, 10, 6, -6, -3,
    -- layer=1 filter=157 channel=62
    14, 0, 15, 2, -11, -13, 1, 4, -15,
    -- layer=1 filter=157 channel=63
    -6, -4, 7, -1, -3, -8, -9, -4, -8,
    -- layer=1 filter=157 channel=64
    -14, 3, 2, -1, 0, -3, -4, -12, -6,
    -- layer=1 filter=157 channel=65
    -1, 1, -3, 4, -6, -3, -11, 0, 0,
    -- layer=1 filter=157 channel=66
    -13, -10, -10, 1, -9, -8, 0, -11, -16,
    -- layer=1 filter=157 channel=67
    6, -5, 2, -4, -7, -7, 5, 11, 0,
    -- layer=1 filter=157 channel=68
    -25, -5, 3, -6, 7, 1, -5, -1, -11,
    -- layer=1 filter=157 channel=69
    15, -4, -1, 6, -4, -10, -15, -2, 1,
    -- layer=1 filter=157 channel=70
    -6, 4, 18, 6, 12, 9, 11, 3, 10,
    -- layer=1 filter=157 channel=71
    -3, -14, -17, -18, -10, -10, -5, -4, -15,
    -- layer=1 filter=157 channel=72
    -2, -2, 2, -1, 0, 5, 0, 5, -3,
    -- layer=1 filter=157 channel=73
    -6, -8, -8, 2, -11, -10, -3, 5, -10,
    -- layer=1 filter=157 channel=74
    -2, -6, 7, -6, -7, -3, -4, 0, 7,
    -- layer=1 filter=157 channel=75
    8, 4, 14, -5, 0, -5, 5, 0, 13,
    -- layer=1 filter=157 channel=76
    -11, -14, -12, -2, -13, -3, -19, -6, -3,
    -- layer=1 filter=157 channel=77
    -10, 1, -6, 1, -13, -3, 2, 0, -5,
    -- layer=1 filter=157 channel=78
    0, -11, 0, -9, -2, -12, 3, -9, 6,
    -- layer=1 filter=157 channel=79
    9, -4, 5, -4, 0, -2, -14, 0, -5,
    -- layer=1 filter=157 channel=80
    7, 0, 4, 5, -11, -9, 9, 1, 1,
    -- layer=1 filter=157 channel=81
    -4, -5, 0, -8, -10, -15, -2, -10, -13,
    -- layer=1 filter=157 channel=82
    -20, -17, -3, -23, -21, -14, -6, 0, -3,
    -- layer=1 filter=157 channel=83
    -3, 3, -2, -8, -12, 3, -2, -8, -9,
    -- layer=1 filter=157 channel=84
    0, 6, 14, 9, -2, 3, 0, -6, 6,
    -- layer=1 filter=157 channel=85
    -8, 1, -4, -2, -8, 3, -3, 0, -9,
    -- layer=1 filter=157 channel=86
    4, -7, 5, -1, -14, 1, -8, -5, -20,
    -- layer=1 filter=157 channel=87
    4, -6, -12, -12, -3, -8, -1, -1, -5,
    -- layer=1 filter=157 channel=88
    -6, -5, 4, -13, -8, -20, 12, 4, -5,
    -- layer=1 filter=157 channel=89
    -6, -9, -4, -5, -11, -11, -4, -12, 0,
    -- layer=1 filter=157 channel=90
    0, -5, -5, -4, -10, 0, -13, -1, 1,
    -- layer=1 filter=157 channel=91
    -6, 1, -11, 7, -10, 2, -4, -2, -4,
    -- layer=1 filter=157 channel=92
    -5, -8, -8, -1, -6, 9, -15, 2, -9,
    -- layer=1 filter=157 channel=93
    -7, -15, 0, -20, -2, -18, -3, -17, -16,
    -- layer=1 filter=157 channel=94
    -1, -14, -6, -6, -13, 2, -12, -7, -19,
    -- layer=1 filter=157 channel=95
    -11, 1, 13, 10, -3, 1, -2, 6, -10,
    -- layer=1 filter=157 channel=96
    4, 3, -7, 2, 7, -3, 1, -6, 6,
    -- layer=1 filter=157 channel=97
    0, -6, 3, -18, -18, -11, -7, -14, 0,
    -- layer=1 filter=157 channel=98
    -13, -13, 2, -3, -2, -1, -11, -8, -10,
    -- layer=1 filter=157 channel=99
    -3, -9, -9, -4, -3, -10, -17, 1, 0,
    -- layer=1 filter=157 channel=100
    -9, 0, -1, -15, -9, -4, -3, -4, -13,
    -- layer=1 filter=157 channel=101
    -11, -12, 1, -7, -7, -10, -11, -12, -4,
    -- layer=1 filter=157 channel=102
    -17, -12, -7, -6, -8, -5, -11, -11, -4,
    -- layer=1 filter=157 channel=103
    -9, -4, 1, 2, 0, 0, -18, -13, -4,
    -- layer=1 filter=157 channel=104
    4, 3, -11, -9, -9, -9, -9, -3, -2,
    -- layer=1 filter=157 channel=105
    -9, 0, 1, 1, -6, -11, -6, -9, -8,
    -- layer=1 filter=157 channel=106
    -3, -11, 0, -5, 1, -8, -1, 2, 6,
    -- layer=1 filter=157 channel=107
    4, -2, 4, -10, 3, -1, 3, -6, -4,
    -- layer=1 filter=157 channel=108
    0, -13, -8, -15, 20, 9, 3, -2, -1,
    -- layer=1 filter=157 channel=109
    1, 11, 5, 9, -7, -3, -3, -3, -8,
    -- layer=1 filter=157 channel=110
    7, 4, 8, -12, 0, 1, -6, 0, -12,
    -- layer=1 filter=157 channel=111
    0, -6, 8, 7, 13, 7, 4, -4, -8,
    -- layer=1 filter=157 channel=112
    -1, -8, 3, -7, 1, -11, -7, -10, -13,
    -- layer=1 filter=157 channel=113
    0, -11, 7, 6, 0, -6, -5, 2, 5,
    -- layer=1 filter=157 channel=114
    14, -4, -9, 0, -16, -5, -11, 2, -9,
    -- layer=1 filter=157 channel=115
    -2, 3, -10, -2, -8, -17, -15, -3, -9,
    -- layer=1 filter=157 channel=116
    -6, -2, -3, 2, -7, 7, -10, -5, 0,
    -- layer=1 filter=157 channel=117
    -8, -4, 12, -3, 10, -4, -15, -4, 9,
    -- layer=1 filter=157 channel=118
    3, -2, -1, -7, 10, 5, -10, -2, -6,
    -- layer=1 filter=157 channel=119
    -16, -17, -14, -10, 5, 1, -12, 4, 5,
    -- layer=1 filter=157 channel=120
    -12, 0, -15, -8, -8, -23, -19, -13, 0,
    -- layer=1 filter=157 channel=121
    -3, -7, -10, 0, 0, 12, -2, 7, -3,
    -- layer=1 filter=157 channel=122
    -2, -8, -9, 0, -5, 0, -4, -6, -8,
    -- layer=1 filter=157 channel=123
    -4, 1, -9, -1, 0, 8, -5, -8, -13,
    -- layer=1 filter=157 channel=124
    -2, -11, 0, -4, 3, -4, 0, 12, 10,
    -- layer=1 filter=157 channel=125
    -15, 12, 2, -1, 9, 3, 5, -3, 5,
    -- layer=1 filter=157 channel=126
    4, 1, -10, 8, 3, -10, 8, -10, -8,
    -- layer=1 filter=157 channel=127
    -13, 1, 1, 0, 1, -2, -4, -7, -2,
    -- layer=1 filter=158 channel=0
    0, 3, 7, -3, -10, -9, -7, 7, 2,
    -- layer=1 filter=158 channel=1
    4, 0, 4, 4, -11, 0, -12, -9, 0,
    -- layer=1 filter=158 channel=2
    0, -11, 8, 0, -5, -5, -8, 4, 7,
    -- layer=1 filter=158 channel=3
    11, 8, 9, -8, 6, 8, -10, -9, 1,
    -- layer=1 filter=158 channel=4
    -1, -11, 0, -1, -12, 6, 3, -3, 7,
    -- layer=1 filter=158 channel=5
    -3, -8, -3, -1, -6, -9, 5, 0, -3,
    -- layer=1 filter=158 channel=6
    7, -3, 4, 2, 5, -10, -1, -6, -10,
    -- layer=1 filter=158 channel=7
    3, 7, 0, -8, -3, -7, -8, -4, -5,
    -- layer=1 filter=158 channel=8
    -6, 5, -2, -12, 5, 3, -8, 0, 0,
    -- layer=1 filter=158 channel=9
    7, -5, -2, 0, 6, 5, -9, -1, -8,
    -- layer=1 filter=158 channel=10
    -1, -2, 6, -7, -9, 9, 10, 9, -3,
    -- layer=1 filter=158 channel=11
    -3, -11, 6, 5, -9, -1, -6, 8, 2,
    -- layer=1 filter=158 channel=12
    4, 4, 5, 5, 4, 5, -4, -9, 7,
    -- layer=1 filter=158 channel=13
    3, -5, -1, 5, 3, 6, 7, 0, 1,
    -- layer=1 filter=158 channel=14
    -5, 0, 9, 7, 7, -5, 0, -6, 8,
    -- layer=1 filter=158 channel=15
    0, 3, 1, 8, 0, -4, -6, -7, -6,
    -- layer=1 filter=158 channel=16
    3, -3, 4, 1, -6, 5, -10, -12, -2,
    -- layer=1 filter=158 channel=17
    5, -1, -5, -7, -5, -5, -9, 1, 2,
    -- layer=1 filter=158 channel=18
    3, -7, -2, 4, 8, -11, -10, -4, -8,
    -- layer=1 filter=158 channel=19
    7, 1, -1, 6, 5, 0, -4, 2, 2,
    -- layer=1 filter=158 channel=20
    7, -11, -12, -1, 5, 4, 0, -2, -7,
    -- layer=1 filter=158 channel=21
    -4, 6, -2, 2, 2, -10, 2, 2, -6,
    -- layer=1 filter=158 channel=22
    1, 0, 5, 7, -8, -3, -1, 3, 0,
    -- layer=1 filter=158 channel=23
    -8, 2, 1, -3, -11, 1, -8, -6, 8,
    -- layer=1 filter=158 channel=24
    -3, -10, -9, -6, -5, -9, 0, 5, -4,
    -- layer=1 filter=158 channel=25
    -7, 0, -5, 10, -9, -1, 0, -2, 7,
    -- layer=1 filter=158 channel=26
    3, -4, 0, -2, 2, -2, 8, 0, 4,
    -- layer=1 filter=158 channel=27
    1, 6, -6, -2, -1, 0, 9, 4, -2,
    -- layer=1 filter=158 channel=28
    -11, -8, -4, 0, -2, -4, 1, -11, -5,
    -- layer=1 filter=158 channel=29
    -4, -7, 9, -8, -1, -3, 4, -5, 0,
    -- layer=1 filter=158 channel=30
    3, -5, -1, 0, 7, 9, -7, -2, -3,
    -- layer=1 filter=158 channel=31
    2, -9, 2, 8, 0, 8, 6, 0, 8,
    -- layer=1 filter=158 channel=32
    -6, 6, -2, -4, -7, 2, -6, -9, -4,
    -- layer=1 filter=158 channel=33
    -3, 1, -1, 2, 0, 3, -6, -5, -9,
    -- layer=1 filter=158 channel=34
    2, -12, -10, 6, -6, -3, -3, -12, -8,
    -- layer=1 filter=158 channel=35
    -11, 4, -10, 4, 6, -5, -4, 3, -4,
    -- layer=1 filter=158 channel=36
    -8, 6, -6, 6, -9, 3, 0, 6, 0,
    -- layer=1 filter=158 channel=37
    0, 3, -7, -4, -1, -6, 6, 4, -1,
    -- layer=1 filter=158 channel=38
    -10, 2, -5, -8, -4, -5, 1, 2, -8,
    -- layer=1 filter=158 channel=39
    2, -12, 0, -5, -5, -3, -10, 6, 6,
    -- layer=1 filter=158 channel=40
    0, -10, -2, -2, -3, 0, 4, 7, 6,
    -- layer=1 filter=158 channel=41
    -2, 1, -5, 3, -5, 6, 8, -4, -6,
    -- layer=1 filter=158 channel=42
    -8, -7, -5, 9, -7, 6, -5, -8, 7,
    -- layer=1 filter=158 channel=43
    -12, -11, -4, -8, 2, -10, -3, 3, 3,
    -- layer=1 filter=158 channel=44
    -3, -5, -5, -10, 7, -8, -1, -10, 2,
    -- layer=1 filter=158 channel=45
    3, 0, 0, 1, 0, -12, -5, 4, -4,
    -- layer=1 filter=158 channel=46
    1, 7, -10, -6, -7, 11, 9, -5, -1,
    -- layer=1 filter=158 channel=47
    -9, 0, -8, 3, -3, 4, -8, -11, -9,
    -- layer=1 filter=158 channel=48
    -6, 6, -7, -11, 2, -9, -3, 0, 7,
    -- layer=1 filter=158 channel=49
    6, -7, -9, 4, -8, 2, -10, -4, -3,
    -- layer=1 filter=158 channel=50
    -12, 0, 0, -1, 3, -6, -12, -5, 7,
    -- layer=1 filter=158 channel=51
    3, 0, 7, -5, -1, 6, -13, -12, 0,
    -- layer=1 filter=158 channel=52
    -2, -7, -2, 3, -2, -6, -7, -4, 0,
    -- layer=1 filter=158 channel=53
    0, 3, 3, -11, -11, -9, 2, 1, -8,
    -- layer=1 filter=158 channel=54
    0, -5, 2, 6, 2, 0, 7, -6, 3,
    -- layer=1 filter=158 channel=55
    -7, 7, 11, -7, 9, -1, 0, -9, 1,
    -- layer=1 filter=158 channel=56
    8, 6, -9, -10, 1, 8, 2, -10, 1,
    -- layer=1 filter=158 channel=57
    -12, 3, 0, -1, 0, 1, -10, 0, -10,
    -- layer=1 filter=158 channel=58
    4, -8, 2, -5, 5, -4, -4, 8, -7,
    -- layer=1 filter=158 channel=59
    -3, -8, 3, 2, 1, -6, 0, 2, 6,
    -- layer=1 filter=158 channel=60
    -1, -5, 2, -7, 8, -5, 7, -6, 1,
    -- layer=1 filter=158 channel=61
    -11, -1, 7, 0, -5, 7, 0, -4, -9,
    -- layer=1 filter=158 channel=62
    -6, 2, 0, -5, -3, 7, -1, -9, 2,
    -- layer=1 filter=158 channel=63
    0, -4, -5, 2, -4, -12, -5, -6, 2,
    -- layer=1 filter=158 channel=64
    0, -9, -7, 1, 3, -8, 7, 0, -3,
    -- layer=1 filter=158 channel=65
    -2, 0, 2, 8, -12, 6, -3, 6, -1,
    -- layer=1 filter=158 channel=66
    3, -1, -2, 1, 0, -11, -5, -4, 7,
    -- layer=1 filter=158 channel=67
    -4, 7, 5, -8, -2, 0, 0, 0, -1,
    -- layer=1 filter=158 channel=68
    -1, 0, 3, -12, 4, -2, 0, 2, 5,
    -- layer=1 filter=158 channel=69
    5, -3, 6, 5, 2, 8, -2, 0, 0,
    -- layer=1 filter=158 channel=70
    11, 9, 4, -3, -5, -7, -3, 4, -12,
    -- layer=1 filter=158 channel=71
    8, -10, 2, -11, -5, 2, -7, 2, -1,
    -- layer=1 filter=158 channel=72
    -4, -4, 2, -7, -4, -9, -1, -2, -9,
    -- layer=1 filter=158 channel=73
    -4, 4, -10, 5, -4, -11, -9, 6, 2,
    -- layer=1 filter=158 channel=74
    -1, 0, -7, -1, -2, -2, -6, -6, 3,
    -- layer=1 filter=158 channel=75
    3, 0, -6, -2, -10, 9, 4, 1, -2,
    -- layer=1 filter=158 channel=76
    7, -2, 4, -3, 1, -11, -8, -1, 0,
    -- layer=1 filter=158 channel=77
    -3, -5, -2, -5, 1, -9, -2, -7, -5,
    -- layer=1 filter=158 channel=78
    5, -8, 7, 0, -1, 0, 0, -2, 0,
    -- layer=1 filter=158 channel=79
    0, 3, 9, -1, 6, 1, -5, 0, 8,
    -- layer=1 filter=158 channel=80
    -6, -5, -4, 3, -4, 4, -3, 7, 4,
    -- layer=1 filter=158 channel=81
    -8, 0, -8, -4, 0, -11, -9, -11, 1,
    -- layer=1 filter=158 channel=82
    3, -6, 4, -11, -5, 1, -4, -1, -2,
    -- layer=1 filter=158 channel=83
    -10, 0, 6, 3, -7, 7, -1, -8, -9,
    -- layer=1 filter=158 channel=84
    1, -4, 0, 7, 0, -11, 0, 7, -8,
    -- layer=1 filter=158 channel=85
    -5, 2, -7, 0, 0, -6, 0, 1, 3,
    -- layer=1 filter=158 channel=86
    -5, 1, -2, 6, -8, 3, -7, -9, 0,
    -- layer=1 filter=158 channel=87
    -5, 6, -6, 5, 3, 3, 1, -5, 4,
    -- layer=1 filter=158 channel=88
    -11, 4, -3, 1, -10, -4, -2, 0, -1,
    -- layer=1 filter=158 channel=89
    -3, -12, -5, -6, -10, -9, 1, -9, 0,
    -- layer=1 filter=158 channel=90
    5, -2, -6, 6, 3, 4, 5, -12, -7,
    -- layer=1 filter=158 channel=91
    -3, -3, -12, 7, -1, -10, 7, -3, 7,
    -- layer=1 filter=158 channel=92
    7, -12, 5, 8, -10, 0, -11, 5, 1,
    -- layer=1 filter=158 channel=93
    7, -5, -10, 3, -11, 0, -7, -3, 6,
    -- layer=1 filter=158 channel=94
    -5, 0, -5, 8, 3, 1, 2, -9, 6,
    -- layer=1 filter=158 channel=95
    -8, 1, 3, -11, -3, 3, -5, 0, -12,
    -- layer=1 filter=158 channel=96
    -1, -4, 0, 8, 1, -7, -6, -7, 7,
    -- layer=1 filter=158 channel=97
    -9, -3, 4, -1, 7, 2, 7, 7, 6,
    -- layer=1 filter=158 channel=98
    -6, 6, -6, -8, 3, 0, -11, 5, -8,
    -- layer=1 filter=158 channel=99
    0, -9, -10, 3, 4, 6, 2, -5, -6,
    -- layer=1 filter=158 channel=100
    2, 0, -2, -5, -11, 6, -11, -7, 8,
    -- layer=1 filter=158 channel=101
    2, -5, -2, 6, 8, 4, -7, -7, 0,
    -- layer=1 filter=158 channel=102
    0, -8, -8, 0, -8, -7, -5, -8, -11,
    -- layer=1 filter=158 channel=103
    -2, -3, -3, -11, 6, -11, 0, -6, 5,
    -- layer=1 filter=158 channel=104
    -3, 6, 1, 5, 0, 7, 0, 3, 0,
    -- layer=1 filter=158 channel=105
    3, 5, 4, -2, 0, 0, 4, -5, -11,
    -- layer=1 filter=158 channel=106
    4, 3, -7, 7, 6, 4, -12, 1, 1,
    -- layer=1 filter=158 channel=107
    4, -8, 4, 7, 8, -10, 8, -6, 9,
    -- layer=1 filter=158 channel=108
    4, -9, 5, -6, -4, 8, 2, 4, -2,
    -- layer=1 filter=158 channel=109
    1, 0, 1, 1, -9, -9, -7, 8, 0,
    -- layer=1 filter=158 channel=110
    5, -8, -8, 3, 0, 0, 3, -10, 1,
    -- layer=1 filter=158 channel=111
    3, -1, -2, 5, 10, -4, 9, -8, 4,
    -- layer=1 filter=158 channel=112
    -10, -2, 0, 0, -9, -4, -8, -7, 3,
    -- layer=1 filter=158 channel=113
    6, 8, 8, -10, -12, 2, 4, -1, -3,
    -- layer=1 filter=158 channel=114
    0, 2, -1, 1, 6, 6, 3, -8, 2,
    -- layer=1 filter=158 channel=115
    1, -10, 3, -8, -11, -11, -1, -2, 1,
    -- layer=1 filter=158 channel=116
    2, 0, 8, -3, 5, 8, -4, 5, 3,
    -- layer=1 filter=158 channel=117
    -10, 3, -2, -3, 1, 0, 6, -8, 5,
    -- layer=1 filter=158 channel=118
    -10, 5, -7, 3, -9, 2, -9, 4, -10,
    -- layer=1 filter=158 channel=119
    -7, -2, -3, 1, 2, -6, 0, -5, 0,
    -- layer=1 filter=158 channel=120
    -11, 6, 0, -2, -11, -1, -11, 8, -6,
    -- layer=1 filter=158 channel=121
    4, 6, -6, 6, -6, -4, 2, 3, -2,
    -- layer=1 filter=158 channel=122
    -5, -4, -9, 10, -1, 0, -7, 5, 8,
    -- layer=1 filter=158 channel=123
    -12, 3, -8, -8, -6, -9, 0, -11, -7,
    -- layer=1 filter=158 channel=124
    6, 6, 1, 1, -1, -1, 3, 6, 9,
    -- layer=1 filter=158 channel=125
    -8, 8, 5, 2, 1, -11, 1, -3, 8,
    -- layer=1 filter=158 channel=126
    -3, 6, 4, -5, 7, -10, -9, -3, 8,
    -- layer=1 filter=158 channel=127
    -2, 8, 0, -8, -5, 2, 0, 6, -4,
    -- layer=1 filter=159 channel=0
    -1, -10, -4, -10, -3, -9, 0, -3, 3,
    -- layer=1 filter=159 channel=1
    -9, -10, 3, -1, -10, 0, 0, 3, 8,
    -- layer=1 filter=159 channel=2
    8, 8, -7, 0, -1, 1, -8, -13, -5,
    -- layer=1 filter=159 channel=3
    -1, 2, 7, -3, -3, 4, 1, 10, 7,
    -- layer=1 filter=159 channel=4
    -4, 0, 0, 6, -1, 4, -4, -10, -9,
    -- layer=1 filter=159 channel=5
    7, 3, 2, 0, 9, -2, 4, -6, -3,
    -- layer=1 filter=159 channel=6
    -7, -10, -7, -4, -3, -5, 6, -9, 5,
    -- layer=1 filter=159 channel=7
    -7, -10, 4, 6, -2, -8, -1, -3, -12,
    -- layer=1 filter=159 channel=8
    -5, -7, 8, 0, 2, -1, 0, 0, 4,
    -- layer=1 filter=159 channel=9
    3, -9, 3, 5, -11, 0, -1, -4, 4,
    -- layer=1 filter=159 channel=10
    2, 5, -4, 1, -5, -12, 0, 6, -11,
    -- layer=1 filter=159 channel=11
    5, 4, -8, -8, -17, 5, -12, 7, -7,
    -- layer=1 filter=159 channel=12
    -8, 0, 6, -6, 1, -5, 2, -6, 1,
    -- layer=1 filter=159 channel=13
    -2, -8, 2, -7, -8, 4, -1, 3, -8,
    -- layer=1 filter=159 channel=14
    -3, 5, 6, 3, -3, 10, -1, -3, 4,
    -- layer=1 filter=159 channel=15
    -2, 0, 5, 10, 3, -4, 6, -5, 6,
    -- layer=1 filter=159 channel=16
    5, 10, 1, 4, 0, 5, -4, -1, -9,
    -- layer=1 filter=159 channel=17
    -9, -11, -6, 8, -10, -6, 0, 2, 3,
    -- layer=1 filter=159 channel=18
    -12, -3, 2, 3, -1, -15, 4, -10, 3,
    -- layer=1 filter=159 channel=19
    -7, -8, -2, 3, -9, 6, 6, 3, -5,
    -- layer=1 filter=159 channel=20
    7, 3, 2, -4, -4, -2, -8, -8, -2,
    -- layer=1 filter=159 channel=21
    -7, 5, 6, 2, -1, 2, -5, 0, -3,
    -- layer=1 filter=159 channel=22
    2, 0, 3, 3, -11, 6, 3, -6, -8,
    -- layer=1 filter=159 channel=23
    -2, 6, 2, 4, -10, -2, -8, -7, 3,
    -- layer=1 filter=159 channel=24
    -8, 6, -4, 3, -11, -9, 0, -10, -14,
    -- layer=1 filter=159 channel=25
    -13, -1, 3, 0, -6, -2, -8, 3, 0,
    -- layer=1 filter=159 channel=26
    -8, -7, 0, -5, 0, 4, 0, -14, -1,
    -- layer=1 filter=159 channel=27
    -4, -10, 4, 3, -9, 5, -6, 7, 4,
    -- layer=1 filter=159 channel=28
    5, -7, -10, 0, -9, -7, 1, -2, -4,
    -- layer=1 filter=159 channel=29
    5, -6, 10, -6, -10, -9, -2, 8, -7,
    -- layer=1 filter=159 channel=30
    5, -1, -7, -10, -8, -13, -3, -8, -2,
    -- layer=1 filter=159 channel=31
    2, 8, -15, -12, -2, -9, -4, -15, 0,
    -- layer=1 filter=159 channel=32
    -7, 1, 6, -5, -5, 5, -1, -5, 7,
    -- layer=1 filter=159 channel=33
    -7, -4, 0, -3, -8, 7, -6, -10, -6,
    -- layer=1 filter=159 channel=34
    -8, -4, -4, 1, 4, -3, -7, -8, -7,
    -- layer=1 filter=159 channel=35
    -3, 0, -8, -4, -9, -3, 1, -4, -8,
    -- layer=1 filter=159 channel=36
    -2, -11, 8, 6, -2, 1, 0, 7, 0,
    -- layer=1 filter=159 channel=37
    -1, 7, -7, -11, -1, 7, 4, 6, -8,
    -- layer=1 filter=159 channel=38
    3, -3, -8, -13, -8, 0, -1, 5, -7,
    -- layer=1 filter=159 channel=39
    3, -5, -8, -9, 1, 0, -8, -10, -9,
    -- layer=1 filter=159 channel=40
    6, -7, -10, -12, -3, -9, -7, -7, 4,
    -- layer=1 filter=159 channel=41
    -5, -2, -5, -4, 4, -7, 7, -14, -5,
    -- layer=1 filter=159 channel=42
    1, 8, -2, 0, -9, 4, -1, -11, 1,
    -- layer=1 filter=159 channel=43
    -9, -11, -7, -2, 1, -4, 5, 5, 4,
    -- layer=1 filter=159 channel=44
    6, -10, 7, -1, -4, -11, -3, 4, -9,
    -- layer=1 filter=159 channel=45
    -5, -3, 7, -5, -5, 0, -13, 3, 5,
    -- layer=1 filter=159 channel=46
    4, -8, 3, 5, -6, -7, 0, 4, -5,
    -- layer=1 filter=159 channel=47
    0, -4, -1, -3, -6, -11, -1, -11, 5,
    -- layer=1 filter=159 channel=48
    -5, -9, -12, 0, -4, 0, -1, 5, 5,
    -- layer=1 filter=159 channel=49
    4, 8, 2, 3, 1, 2, 2, 2, 3,
    -- layer=1 filter=159 channel=50
    0, 0, 6, 5, -8, -9, -10, -3, -2,
    -- layer=1 filter=159 channel=51
    -8, -11, -7, -4, 4, -4, -3, 7, 4,
    -- layer=1 filter=159 channel=52
    5, -8, -7, -9, 7, 2, 7, -10, -3,
    -- layer=1 filter=159 channel=53
    -8, -6, 5, 0, -6, 0, 2, 4, -3,
    -- layer=1 filter=159 channel=54
    0, -7, 7, 0, -6, -7, 5, -8, 0,
    -- layer=1 filter=159 channel=55
    8, 6, 4, -6, -4, 4, 7, 4, -11,
    -- layer=1 filter=159 channel=56
    -8, -10, -9, 2, -11, 0, -6, 3, 3,
    -- layer=1 filter=159 channel=57
    2, -10, 7, -11, 7, -5, -10, -3, 5,
    -- layer=1 filter=159 channel=58
    0, 3, -5, -5, -1, -10, -7, -10, 5,
    -- layer=1 filter=159 channel=59
    0, 4, -5, 7, 6, 1, 1, -10, 8,
    -- layer=1 filter=159 channel=60
    0, -5, 7, -9, 7, 8, 10, -4, 7,
    -- layer=1 filter=159 channel=61
    -4, -8, 6, 3, 8, -8, 0, 6, -6,
    -- layer=1 filter=159 channel=62
    -2, 4, 1, -3, -3, 4, -4, -8, 0,
    -- layer=1 filter=159 channel=63
    -8, -5, -10, -7, 1, 2, 3, -11, 0,
    -- layer=1 filter=159 channel=64
    -1, 0, 6, 2, -7, 8, 0, -3, 6,
    -- layer=1 filter=159 channel=65
    -2, -6, 0, -12, 1, 1, 0, -11, -8,
    -- layer=1 filter=159 channel=66
    3, -2, -6, 1, -5, -11, 2, -7, -6,
    -- layer=1 filter=159 channel=67
    -6, -1, -9, -9, -5, -2, -6, 4, -7,
    -- layer=1 filter=159 channel=68
    2, -10, -7, 5, 6, 2, -1, -1, 4,
    -- layer=1 filter=159 channel=69
    0, -4, 12, -4, -9, 0, -6, 7, -8,
    -- layer=1 filter=159 channel=70
    -8, 9, 0, 1, 0, -9, 5, -7, -4,
    -- layer=1 filter=159 channel=71
    -13, -2, 0, -9, -3, -3, -1, -6, -9,
    -- layer=1 filter=159 channel=72
    -5, 7, -2, 2, 2, -3, 3, 1, -1,
    -- layer=1 filter=159 channel=73
    -10, -5, -3, 7, 0, -2, 3, 3, -9,
    -- layer=1 filter=159 channel=74
    0, 4, -2, 5, 4, -11, 7, 5, -7,
    -- layer=1 filter=159 channel=75
    0, -8, -6, -2, -13, -12, 0, -9, 15,
    -- layer=1 filter=159 channel=76
    -5, 2, -4, 4, -5, -6, -5, 0, 0,
    -- layer=1 filter=159 channel=77
    -11, -4, 0, -8, -2, -4, -8, -4, -4,
    -- layer=1 filter=159 channel=78
    -4, -1, -3, -2, -4, -10, -7, -3, 5,
    -- layer=1 filter=159 channel=79
    0, 8, -11, -7, 4, 4, 1, -6, -9,
    -- layer=1 filter=159 channel=80
    9, -4, 0, 6, 1, 7, 0, -8, 1,
    -- layer=1 filter=159 channel=81
    1, 8, 8, -3, -11, 4, 0, -11, 1,
    -- layer=1 filter=159 channel=82
    8, 4, 4, 4, -5, -7, -2, 0, -4,
    -- layer=1 filter=159 channel=83
    7, -11, -11, 0, -8, -6, -1, 2, 4,
    -- layer=1 filter=159 channel=84
    -6, -4, -11, -4, 0, 6, -4, 2, 0,
    -- layer=1 filter=159 channel=85
    1, 5, -9, 5, 5, 4, 6, -5, 6,
    -- layer=1 filter=159 channel=86
    -7, -17, -4, 3, -4, -12, -1, -8, 5,
    -- layer=1 filter=159 channel=87
    0, 1, -3, 4, -10, 0, 6, -5, 8,
    -- layer=1 filter=159 channel=88
    -6, 2, 7, -6, -9, 3, -6, -9, -6,
    -- layer=1 filter=159 channel=89
    6, 7, -3, 4, -1, -10, -7, -7, -1,
    -- layer=1 filter=159 channel=90
    2, 1, -8, 1, -12, -8, -8, -8, -4,
    -- layer=1 filter=159 channel=91
    -8, -10, -4, -1, 0, 1, 5, 1, 2,
    -- layer=1 filter=159 channel=92
    5, -6, 4, 0, 6, 3, 4, -8, -11,
    -- layer=1 filter=159 channel=93
    -12, -7, 3, -5, 0, 0, -7, -11, -5,
    -- layer=1 filter=159 channel=94
    -11, 1, 5, -2, -10, 4, 0, -4, 2,
    -- layer=1 filter=159 channel=95
    1, -1, -10, -4, 7, 0, 0, 0, 2,
    -- layer=1 filter=159 channel=96
    6, -1, -5, -5, -5, -11, -4, -7, -1,
    -- layer=1 filter=159 channel=97
    -11, -9, 6, 3, 1, 4, 4, 8, 1,
    -- layer=1 filter=159 channel=98
    0, -1, -11, -9, -4, -6, 7, -11, -5,
    -- layer=1 filter=159 channel=99
    2, 0, 7, -10, 5, 6, 0, -9, -4,
    -- layer=1 filter=159 channel=100
    -1, -8, 7, -3, -13, -6, 3, -11, -5,
    -- layer=1 filter=159 channel=101
    5, 5, -8, 5, -5, 7, 5, 8, 2,
    -- layer=1 filter=159 channel=102
    6, -4, 1, 1, -10, -7, -11, 5, 7,
    -- layer=1 filter=159 channel=103
    -1, -6, 5, -7, -5, 0, -8, -5, -1,
    -- layer=1 filter=159 channel=104
    5, -5, -5, 7, 4, 6, -9, -11, 0,
    -- layer=1 filter=159 channel=105
    -1, -2, -4, -7, -7, 8, -4, -3, 1,
    -- layer=1 filter=159 channel=106
    6, -3, 0, -9, 3, 0, 0, -5, -1,
    -- layer=1 filter=159 channel=107
    -3, -3, 8, -2, 0, 5, 1, -1, 10,
    -- layer=1 filter=159 channel=108
    -5, 0, 7, 0, -3, -2, -13, -10, 6,
    -- layer=1 filter=159 channel=109
    -8, 0, -1, -2, 9, 1, 0, 0, 7,
    -- layer=1 filter=159 channel=110
    -8, -7, 0, -7, 4, 0, -2, 4, -5,
    -- layer=1 filter=159 channel=111
    -7, 1, -13, 3, 4, 2, -7, 6, 3,
    -- layer=1 filter=159 channel=112
    -8, -7, 6, 0, 5, -4, -10, 8, -10,
    -- layer=1 filter=159 channel=113
    0, -1, -8, 1, -6, -13, -12, 0, -4,
    -- layer=1 filter=159 channel=114
    2, -1, -5, -2, 0, 8, -7, -9, -4,
    -- layer=1 filter=159 channel=115
    -17, -3, 5, -8, -3, -7, 3, -1, -1,
    -- layer=1 filter=159 channel=116
    6, -7, 0, 1, 3, 1, 8, 0, 4,
    -- layer=1 filter=159 channel=117
    8, -8, -3, 0, 8, -2, -7, 7, 9,
    -- layer=1 filter=159 channel=118
    2, -16, -8, 0, -5, -1, 3, -8, -9,
    -- layer=1 filter=159 channel=119
    0, -9, 6, 6, -6, 4, -10, 0, -3,
    -- layer=1 filter=159 channel=120
    4, 0, 8, 0, 6, -4, 2, -12, -2,
    -- layer=1 filter=159 channel=121
    -8, -1, -1, -7, -9, -1, -1, 2, 14,
    -- layer=1 filter=159 channel=122
    -5, 5, 5, 2, -1, 3, -5, 6, -9,
    -- layer=1 filter=159 channel=123
    0, -1, -9, -12, -2, -6, 5, 5, 7,
    -- layer=1 filter=159 channel=124
    -1, 2, 7, 10, -9, 4, -1, 3, -8,
    -- layer=1 filter=159 channel=125
    3, -11, 9, 3, -5, 7, 0, -10, -2,
    -- layer=1 filter=159 channel=126
    -2, -2, -7, 5, -2, 2, -12, -11, -2,
    -- layer=1 filter=159 channel=127
    -12, -5, 0, -9, 0, 0, 0, -10, 8,
    -- layer=1 filter=160 channel=0
    5, 5, 1, 6, 1, 0, -3, 6, -5,
    -- layer=1 filter=160 channel=1
    0, -10, -4, 3, 1, -6, 6, -9, 0,
    -- layer=1 filter=160 channel=2
    0, 0, -8, 3, -6, 5, -4, -8, -1,
    -- layer=1 filter=160 channel=3
    -6, 7, 3, 9, 8, 4, 8, 9, 3,
    -- layer=1 filter=160 channel=4
    -6, 0, -3, 0, 8, -6, 0, -9, -2,
    -- layer=1 filter=160 channel=5
    -3, -7, -3, -4, 3, -1, 0, 8, -6,
    -- layer=1 filter=160 channel=6
    -1, -6, -8, 0, -7, 7, 6, -9, -7,
    -- layer=1 filter=160 channel=7
    -3, -4, 0, -1, -12, 7, -1, 0, 7,
    -- layer=1 filter=160 channel=8
    -3, 5, -6, -8, 4, -10, 0, 6, 5,
    -- layer=1 filter=160 channel=9
    0, 0, -1, -5, -5, 4, 0, -5, -5,
    -- layer=1 filter=160 channel=10
    -4, 0, -3, -9, -2, 5, -1, 5, -6,
    -- layer=1 filter=160 channel=11
    8, -1, 7, -7, 7, -5, 2, -2, -11,
    -- layer=1 filter=160 channel=12
    1, -7, -5, -10, -9, 4, -9, 9, -5,
    -- layer=1 filter=160 channel=13
    3, 9, 0, -12, 5, -9, 2, -1, -6,
    -- layer=1 filter=160 channel=14
    -6, 11, 7, 2, -1, -6, 10, 11, -3,
    -- layer=1 filter=160 channel=15
    4, 4, -1, 7, 4, -4, -2, 1, -11,
    -- layer=1 filter=160 channel=16
    -8, -11, 0, -4, -7, 1, 7, -7, -13,
    -- layer=1 filter=160 channel=17
    5, 4, -8, -9, -5, -11, -10, -8, -2,
    -- layer=1 filter=160 channel=18
    -9, -8, -10, 2, 1, 2, 7, -5, -5,
    -- layer=1 filter=160 channel=19
    -9, 0, -11, -6, -11, 0, -1, -1, -1,
    -- layer=1 filter=160 channel=20
    -7, -5, -3, -11, 0, 0, 0, -2, -4,
    -- layer=1 filter=160 channel=21
    -4, -1, 2, -4, 0, 2, -5, -10, 5,
    -- layer=1 filter=160 channel=22
    9, -1, 0, 8, 2, 0, -2, -3, -10,
    -- layer=1 filter=160 channel=23
    6, -4, 7, 5, 8, -2, 0, 1, -10,
    -- layer=1 filter=160 channel=24
    4, 9, -1, -1, -9, 2, 0, -1, -7,
    -- layer=1 filter=160 channel=25
    3, 9, -6, 6, 0, -7, 3, -4, -6,
    -- layer=1 filter=160 channel=26
    -4, 2, -2, -5, 5, -5, 6, -4, -2,
    -- layer=1 filter=160 channel=27
    -3, -10, 5, 4, 0, -3, -4, -5, -1,
    -- layer=1 filter=160 channel=28
    -8, -2, 0, 2, 3, 0, 5, -12, 1,
    -- layer=1 filter=160 channel=29
    -9, 0, -6, 4, 8, 4, 5, -10, 0,
    -- layer=1 filter=160 channel=30
    2, 9, 10, -6, 2, -10, 5, 8, -4,
    -- layer=1 filter=160 channel=31
    -3, 5, 0, -9, -3, -4, -7, -7, -2,
    -- layer=1 filter=160 channel=32
    -4, 3, -3, -11, -11, -9, -8, 4, -7,
    -- layer=1 filter=160 channel=33
    -4, 0, -8, -2, -1, -7, 1, -3, -6,
    -- layer=1 filter=160 channel=34
    0, 5, -10, -8, -2, 2, 4, 4, -10,
    -- layer=1 filter=160 channel=35
    9, -10, 1, 3, -9, -6, -8, 6, 0,
    -- layer=1 filter=160 channel=36
    0, 0, -6, 7, -6, 3, 3, 0, -11,
    -- layer=1 filter=160 channel=37
    -5, -4, -11, 0, 10, 10, -4, -6, -5,
    -- layer=1 filter=160 channel=38
    -9, -5, 3, -7, 2, -11, 0, -1, -4,
    -- layer=1 filter=160 channel=39
    -9, 5, -7, 1, -7, 2, -2, 6, -1,
    -- layer=1 filter=160 channel=40
    4, -3, 6, 8, 5, -5, -15, -8, 0,
    -- layer=1 filter=160 channel=41
    -7, 7, 5, 7, -2, 3, -3, -8, -11,
    -- layer=1 filter=160 channel=42
    9, -2, -7, 6, -10, 9, 1, -8, -4,
    -- layer=1 filter=160 channel=43
    -2, 6, 6, 5, -2, 8, 8, -7, -4,
    -- layer=1 filter=160 channel=44
    4, 4, -11, -9, -7, 3, -8, 3, 6,
    -- layer=1 filter=160 channel=45
    0, 3, -7, 4, -11, -10, -11, -3, -4,
    -- layer=1 filter=160 channel=46
    -7, 8, 0, 6, 7, 3, -2, 0, -8,
    -- layer=1 filter=160 channel=47
    -7, -7, 7, 0, 6, -12, 3, -10, -12,
    -- layer=1 filter=160 channel=48
    5, -12, 0, -10, 6, -7, 6, -1, -8,
    -- layer=1 filter=160 channel=49
    0, -6, 3, -2, -11, 7, 6, 2, -6,
    -- layer=1 filter=160 channel=50
    6, 0, -3, 0, -9, 7, 1, 4, 3,
    -- layer=1 filter=160 channel=51
    9, 4, -11, -6, -3, -5, 5, -14, 1,
    -- layer=1 filter=160 channel=52
    -5, 10, -5, 0, 3, 5, -6, -3, -6,
    -- layer=1 filter=160 channel=53
    0, 7, 8, -4, 7, -11, 0, -8, -3,
    -- layer=1 filter=160 channel=54
    5, 7, -3, -2, -4, 10, -2, -2, -5,
    -- layer=1 filter=160 channel=55
    -12, -9, 4, -6, -4, -7, -1, -4, -2,
    -- layer=1 filter=160 channel=56
    5, 6, -7, 4, 3, -4, 4, 0, -9,
    -- layer=1 filter=160 channel=57
    7, 0, -10, -5, -6, 1, -11, -8, 0,
    -- layer=1 filter=160 channel=58
    -2, 7, -7, 0, 0, 2, 1, 5, -4,
    -- layer=1 filter=160 channel=59
    5, -2, 2, -7, 2, -2, 6, -7, -3,
    -- layer=1 filter=160 channel=60
    -7, 0, -9, -6, -1, 4, 2, -8, 6,
    -- layer=1 filter=160 channel=61
    1, 6, -4, 3, -11, 2, -1, -2, -5,
    -- layer=1 filter=160 channel=62
    5, 7, -6, 4, 0, -8, 7, 0, -10,
    -- layer=1 filter=160 channel=63
    -2, -6, -2, -1, -11, 0, -8, 0, -3,
    -- layer=1 filter=160 channel=64
    2, -2, -9, 5, 8, -10, -10, 6, 6,
    -- layer=1 filter=160 channel=65
    2, 2, 0, -11, -4, 3, 0, 2, -2,
    -- layer=1 filter=160 channel=66
    -7, -9, 1, -8, 0, -2, 0, -8, -7,
    -- layer=1 filter=160 channel=67
    -1, 7, -2, 8, -3, 8, 1, -5, 4,
    -- layer=1 filter=160 channel=68
    12, 1, -11, 0, -4, 7, -11, -10, -5,
    -- layer=1 filter=160 channel=69
    9, -7, 3, -6, -5, 3, -6, 3, 2,
    -- layer=1 filter=160 channel=70
    -9, 8, 7, -3, 3, 4, 1, 1, 6,
    -- layer=1 filter=160 channel=71
    -10, -6, 0, -1, -2, -7, -12, 4, -6,
    -- layer=1 filter=160 channel=72
    3, -8, -10, -4, 0, -1, 6, -3, -10,
    -- layer=1 filter=160 channel=73
    0, 7, 5, -7, 1, 5, 2, 5, 6,
    -- layer=1 filter=160 channel=74
    4, 0, -1, 5, 0, -4, -3, -7, 2,
    -- layer=1 filter=160 channel=75
    -13, 5, -7, -1, 0, 8, -11, -10, 0,
    -- layer=1 filter=160 channel=76
    -1, 2, -9, 7, -8, -5, -6, -11, 0,
    -- layer=1 filter=160 channel=77
    7, -3, -2, 1, -8, 2, -8, 4, -6,
    -- layer=1 filter=160 channel=78
    -5, -10, 6, 4, -2, 6, 2, -10, 7,
    -- layer=1 filter=160 channel=79
    4, -6, 5, 6, -8, -3, 8, 0, 5,
    -- layer=1 filter=160 channel=80
    0, -10, -5, 9, 1, 0, 5, 5, 4,
    -- layer=1 filter=160 channel=81
    -10, -8, 2, 3, -12, -10, -10, 1, 3,
    -- layer=1 filter=160 channel=82
    2, 5, -11, -8, -6, -2, -5, -2, -6,
    -- layer=1 filter=160 channel=83
    -8, -8, 8, 8, -1, -6, 0, 1, -10,
    -- layer=1 filter=160 channel=84
    -5, 8, -9, -3, -1, -3, 3, -9, -6,
    -- layer=1 filter=160 channel=85
    -6, 8, -10, 4, 0, 4, 5, -4, -6,
    -- layer=1 filter=160 channel=86
    6, 2, 6, 8, -11, 2, 1, -10, -5,
    -- layer=1 filter=160 channel=87
    6, -1, -8, -8, -7, -3, 4, -12, -3,
    -- layer=1 filter=160 channel=88
    0, 1, -12, -9, -10, 1, -7, -4, -2,
    -- layer=1 filter=160 channel=89
    -2, 7, 8, 5, 5, 5, -9, -5, 0,
    -- layer=1 filter=160 channel=90
    1, -12, 6, -2, 0, 6, 8, -2, 8,
    -- layer=1 filter=160 channel=91
    9, -7, -5, -1, 0, -13, 8, -5, -7,
    -- layer=1 filter=160 channel=92
    -4, -12, -8, 5, 0, 0, -10, -6, -5,
    -- layer=1 filter=160 channel=93
    4, -6, -10, 0, 5, -5, -2, -3, -2,
    -- layer=1 filter=160 channel=94
    7, -9, 4, -8, -2, 2, -9, -1, 0,
    -- layer=1 filter=160 channel=95
    -6, -4, 7, -7, -7, -3, -3, 4, 3,
    -- layer=1 filter=160 channel=96
    6, 5, 2, -6, -7, -3, -3, -3, -5,
    -- layer=1 filter=160 channel=97
    -8, 8, 0, -9, 0, -2, 8, -10, 0,
    -- layer=1 filter=160 channel=98
    7, -2, 3, 4, -6, 10, -10, -10, -7,
    -- layer=1 filter=160 channel=99
    -1, 3, -2, 0, -7, 5, -8, -7, -7,
    -- layer=1 filter=160 channel=100
    7, 0, -2, -6, 8, -5, -4, -7, -6,
    -- layer=1 filter=160 channel=101
    -9, -5, 0, -5, -1, -3, -8, 1, -1,
    -- layer=1 filter=160 channel=102
    -4, 6, -8, 5, 8, -1, -5, 8, -7,
    -- layer=1 filter=160 channel=103
    0, 6, -2, 3, -11, -5, -2, 1, -3,
    -- layer=1 filter=160 channel=104
    3, -5, -5, -7, -5, -5, -12, 8, 0,
    -- layer=1 filter=160 channel=105
    6, -2, -2, 3, -3, 7, -2, -5, -11,
    -- layer=1 filter=160 channel=106
    -7, -3, 4, -7, 0, 7, -1, -1, -1,
    -- layer=1 filter=160 channel=107
    -2, 7, -10, 4, 11, 1, 1, 3, 0,
    -- layer=1 filter=160 channel=108
    7, 4, 5, 1, -10, 0, -1, -8, 5,
    -- layer=1 filter=160 channel=109
    6, -10, 5, -3, -9, 2, 1, 2, -6,
    -- layer=1 filter=160 channel=110
    0, -4, 4, -11, 0, -2, 5, 1, -6,
    -- layer=1 filter=160 channel=111
    -8, 9, 5, -10, 1, 0, 4, 5, -3,
    -- layer=1 filter=160 channel=112
    5, -11, 0, -5, 3, -4, 1, 8, -11,
    -- layer=1 filter=160 channel=113
    -5, 3, 5, 5, -1, 3, -4, 0, 7,
    -- layer=1 filter=160 channel=114
    -4, 6, -8, -7, 7, -10, -3, -9, 0,
    -- layer=1 filter=160 channel=115
    0, 1, 5, -8, -11, -2, -4, 9, 2,
    -- layer=1 filter=160 channel=116
    7, 10, 10, -10, -2, -9, 8, 11, 7,
    -- layer=1 filter=160 channel=117
    -2, -7, 1, 5, -1, 3, 3, 1, 4,
    -- layer=1 filter=160 channel=118
    6, -3, -8, -1, -2, 0, -5, -3, -7,
    -- layer=1 filter=160 channel=119
    -11, -5, -8, 0, -10, -7, 0, -5, -3,
    -- layer=1 filter=160 channel=120
    -13, -10, 3, 6, -1, -4, -10, 7, -3,
    -- layer=1 filter=160 channel=121
    1, -7, 6, -4, 2, -4, 3, 8, -3,
    -- layer=1 filter=160 channel=122
    1, -7, -8, 7, 6, 0, 10, -6, 7,
    -- layer=1 filter=160 channel=123
    6, -6, -5, -9, -10, 0, -3, -4, 4,
    -- layer=1 filter=160 channel=124
    -4, -8, -11, 6, 0, 8, -4, -10, -4,
    -- layer=1 filter=160 channel=125
    -10, 6, 0, -2, 6, -8, -2, 0, -8,
    -- layer=1 filter=160 channel=126
    6, -9, -1, 3, 9, -4, 4, 1, -7,
    -- layer=1 filter=160 channel=127
    -8, 6, -5, -9, 1, 5, -1, 0, -3,
    -- layer=1 filter=161 channel=0
    3, 5, -4, 24, 19, -14, 9, 2, -19,
    -- layer=1 filter=161 channel=1
    16, 50, -9, 11, -23, -6, 6, -68, -26,
    -- layer=1 filter=161 channel=2
    38, -27, 3, -17, -50, 12, -33, -51, -4,
    -- layer=1 filter=161 channel=3
    -1, 0, 12, 10, 8, 10, 0, 4, -12,
    -- layer=1 filter=161 channel=4
    1, -2, 8, -6, 1, 3, 0, -5, -6,
    -- layer=1 filter=161 channel=5
    36, 39, -14, -22, -63, 12, 0, -64, -23,
    -- layer=1 filter=161 channel=6
    -28, -40, 33, -31, -18, 60, 29, 31, 84,
    -- layer=1 filter=161 channel=7
    20, 42, -62, 34, -21, -59, 7, -43, -53,
    -- layer=1 filter=161 channel=8
    37, 54, 11, 24, 4, 3, 13, -72, -6,
    -- layer=1 filter=161 channel=9
    0, 12, 18, 6, -6, 32, 3, 30, 32,
    -- layer=1 filter=161 channel=10
    30, 38, -77, 14, -4, -52, 0, -24, -64,
    -- layer=1 filter=161 channel=11
    5, 20, 9, 18, 25, 0, 19, 17, 3,
    -- layer=1 filter=161 channel=12
    -15, 33, 20, 3, -84, -70, -12, -32, 9,
    -- layer=1 filter=161 channel=13
    -41, -7, 29, -30, -1, 41, -16, 27, 31,
    -- layer=1 filter=161 channel=14
    -17, 23, -68, 15, -31, -43, -23, -22, -42,
    -- layer=1 filter=161 channel=15
    -36, 20, -32, -27, -91, 9, -27, -35, -24,
    -- layer=1 filter=161 channel=16
    42, 41, -11, 6, -53, -26, 10, -66, -44,
    -- layer=1 filter=161 channel=17
    9, 12, -5, 1, 12, -5, -4, -8, -3,
    -- layer=1 filter=161 channel=18
    -4, -16, 19, -22, -4, -15, 12, -14, 1,
    -- layer=1 filter=161 channel=19
    39, -29, -3, -100, -32, -27, -17, -14, -38,
    -- layer=1 filter=161 channel=20
    -18, 5, 19, -25, -5, 8, -2, 10, 20,
    -- layer=1 filter=161 channel=21
    -29, -18, -12, -4, -17, 0, 11, -2, 21,
    -- layer=1 filter=161 channel=22
    -12, 0, 17, -18, 0, 21, -24, -12, 8,
    -- layer=1 filter=161 channel=23
    -28, -33, -55, -13, -40, -75, -5, -61, -14,
    -- layer=1 filter=161 channel=24
    -20, -29, 12, -45, -4, -7, -26, -18, 13,
    -- layer=1 filter=161 channel=25
    42, 28, -53, 33, -54, -30, 5, -65, -78,
    -- layer=1 filter=161 channel=26
    -55, 7, 52, -47, 29, 47, -5, 6, 27,
    -- layer=1 filter=161 channel=27
    12, 15, -21, 5, -7, -7, 6, 12, 10,
    -- layer=1 filter=161 channel=28
    15, 34, -64, 22, -18, -60, 1, -19, -49,
    -- layer=1 filter=161 channel=29
    -9, -1, -27, 7, -10, -15, 1, 2, -7,
    -- layer=1 filter=161 channel=30
    7, -42, 0, -31, -12, 0, 19, -16, 17,
    -- layer=1 filter=161 channel=31
    -27, -25, -6, -10, -48, -37, 3, -32, -9,
    -- layer=1 filter=161 channel=32
    -88, 1, 24, 0, 17, 41, 11, 20, 29,
    -- layer=1 filter=161 channel=33
    1, 9, 6, 8, 19, 7, 6, 16, -4,
    -- layer=1 filter=161 channel=34
    30, -21, 16, 16, -2, 30, 15, 20, 21,
    -- layer=1 filter=161 channel=35
    -4, -8, -12, -4, -16, -8, -15, -6, -2,
    -- layer=1 filter=161 channel=36
    36, 30, 15, 25, 24, -2, 25, 20, 10,
    -- layer=1 filter=161 channel=37
    39, 17, -44, -10, -72, -20, -9, -62, -43,
    -- layer=1 filter=161 channel=38
    -33, -24, 19, -43, 0, 38, -9, 31, 36,
    -- layer=1 filter=161 channel=39
    25, 22, -18, 13, 5, -22, 10, -20, -13,
    -- layer=1 filter=161 channel=40
    -35, -16, -11, -37, -45, 10, -8, -5, 30,
    -- layer=1 filter=161 channel=41
    35, -12, 24, -2, 7, 21, 20, -1, 21,
    -- layer=1 filter=161 channel=42
    21, 6, -5, 16, -17, -7, -32, -98, -44,
    -- layer=1 filter=161 channel=43
    16, 34, -29, 38, -34, -31, 4, -60, -58,
    -- layer=1 filter=161 channel=44
    -55, 33, 54, 8, 40, 50, 4, 31, 31,
    -- layer=1 filter=161 channel=45
    -22, -12, 7, -26, -5, 26, -13, 10, 0,
    -- layer=1 filter=161 channel=46
    15, -45, -31, -75, -79, -51, -57, -73, -47,
    -- layer=1 filter=161 channel=47
    -25, -72, -83, -40, -59, -28, -18, -27, 18,
    -- layer=1 filter=161 channel=48
    -6, -29, -5, -14, -7, 3, 12, 0, 21,
    -- layer=1 filter=161 channel=49
    -15, -42, -21, -33, -19, 18, -20, 15, 46,
    -- layer=1 filter=161 channel=50
    -15, -4, 17, -22, 13, 13, -7, 19, -2,
    -- layer=1 filter=161 channel=51
    -10, 3, -10, -7, 12, 18, -3, 13, 19,
    -- layer=1 filter=161 channel=52
    10, 14, -6, -3, 11, 2, 13, 18, 6,
    -- layer=1 filter=161 channel=53
    -4, -4, 1, -2, 6, -8, 2, -8, -9,
    -- layer=1 filter=161 channel=54
    26, 19, -53, 3, -68, 4, -19, -52, -65,
    -- layer=1 filter=161 channel=55
    22, 0, -12, 24, 16, -8, 11, 2, -6,
    -- layer=1 filter=161 channel=56
    4, 3, -6, 0, -10, -11, -2, 1, -4,
    -- layer=1 filter=161 channel=57
    12, 0, -70, 11, -19, -10, -6, -17, -24,
    -- layer=1 filter=161 channel=58
    24, -63, -143, -5, -82, -139, 17, -90, -40,
    -- layer=1 filter=161 channel=59
    11, 2, -11, 13, -2, -8, -1, -8, -1,
    -- layer=1 filter=161 channel=60
    4, 16, 11, 12, 16, 18, 6, 7, 2,
    -- layer=1 filter=161 channel=61
    2, 7, 7, 5, -3, 6, -3, 9, 5,
    -- layer=1 filter=161 channel=62
    39, 30, -11, -8, -23, -27, -20, -78, -28,
    -- layer=1 filter=161 channel=63
    5, 19, -1, 32, 9, 1, 29, 19, -10,
    -- layer=1 filter=161 channel=64
    -8, -10, 0, 0, 0, 9, 0, -9, 4,
    -- layer=1 filter=161 channel=65
    -23, -5, 19, -3, 1, 5, 16, 14, 16,
    -- layer=1 filter=161 channel=66
    9, 20, -18, 33, 14, -3, 2, 5, -7,
    -- layer=1 filter=161 channel=67
    -32, -40, -2, -16, -14, 18, -16, 2, 26,
    -- layer=1 filter=161 channel=68
    -52, 27, 58, 0, 41, 52, 19, 27, 14,
    -- layer=1 filter=161 channel=69
    -4, 7, -4, -44, -35, -6, -35, -36, -43,
    -- layer=1 filter=161 channel=70
    -37, -38, 17, -35, -45, -7, -37, -16, 34,
    -- layer=1 filter=161 channel=71
    -1, 0, -37, 14, -11, -29, 4, -33, -40,
    -- layer=1 filter=161 channel=72
    19, -57, 28, -43, -15, -1, 5, 5, 1,
    -- layer=1 filter=161 channel=73
    7, 5, -10, -5, -1, 0, 8, -9, -7,
    -- layer=1 filter=161 channel=74
    -47, 18, 57, -32, 26, 7, 22, 17, -12,
    -- layer=1 filter=161 channel=75
    -16, -1, -37, -6, -57, -72, 6, -37, 15,
    -- layer=1 filter=161 channel=76
    -33, -3, 27, -8, 27, 40, 15, 24, 15,
    -- layer=1 filter=161 channel=77
    -12, -27, -13, 11, -29, -10, 4, 0, -3,
    -- layer=1 filter=161 channel=78
    13, 9, -12, 4, 10, -8, -1, 7, 2,
    -- layer=1 filter=161 channel=79
    33, 23, 0, 1, -32, -24, -2, -39, -26,
    -- layer=1 filter=161 channel=80
    -8, -6, 1, 10, -10, 0, 6, -9, -10,
    -- layer=1 filter=161 channel=81
    20, -24, -32, 10, -23, -37, 6, -39, -25,
    -- layer=1 filter=161 channel=82
    -24, -23, 7, 4, -13, 12, 9, 9, 34,
    -- layer=1 filter=161 channel=83
    6, 26, 5, -20, -9, 7, -33, -36, 0,
    -- layer=1 filter=161 channel=84
    -19, 13, 68, -24, 30, 47, 32, 12, 16,
    -- layer=1 filter=161 channel=85
    27, -65, -50, -1, -23, -75, 25, -27, 0,
    -- layer=1 filter=161 channel=86
    17, 26, -26, 26, 5, -14, 0, -10, -26,
    -- layer=1 filter=161 channel=87
    29, -37, 9, -58, 19, -1, 9, 22, 7,
    -- layer=1 filter=161 channel=88
    -10, -17, -1, -2, 3, 8, 12, 22, 18,
    -- layer=1 filter=161 channel=89
    -17, -20, 23, -9, -14, 19, 1, 21, 18,
    -- layer=1 filter=161 channel=90
    -28, 10, 48, -33, 21, 45, -26, 0, 11,
    -- layer=1 filter=161 channel=91
    -17, -13, 4, -21, -12, 8, -9, -2, 27,
    -- layer=1 filter=161 channel=92
    -51, 33, -48, 0, -11, 17, -17, -11, -35,
    -- layer=1 filter=161 channel=93
    -12, 12, 0, 5, 1, -4, -3, 0, -6,
    -- layer=1 filter=161 channel=94
    7, 15, -21, 31, 25, -12, 15, 14, -27,
    -- layer=1 filter=161 channel=95
    -22, 7, 47, -16, 11, 38, 2, 32, 5,
    -- layer=1 filter=161 channel=96
    3, -4, 0, 5, 0, 7, 4, 11, 6,
    -- layer=1 filter=161 channel=97
    16, 11, 0, 8, 13, -19, 10, -2, -20,
    -- layer=1 filter=161 channel=98
    44, 33, -4, 17, -19, -15, -27, -58, -38,
    -- layer=1 filter=161 channel=99
    -35, 17, -40, -14, -8, -81, -51, 14, -81,
    -- layer=1 filter=161 channel=100
    -6, 4, 20, 13, 21, -4, 12, 6, 15,
    -- layer=1 filter=161 channel=101
    -30, -7, 16, -14, 0, 30, -8, 15, 19,
    -- layer=1 filter=161 channel=102
    2, 1, -12, 7, 12, 0, 8, 8, -17,
    -- layer=1 filter=161 channel=103
    1, 16, 7, 0, 4, -12, 20, -4, 12,
    -- layer=1 filter=161 channel=104
    -18, -33, -44, -28, 23, -37, 6, 15, -8,
    -- layer=1 filter=161 channel=105
    22, 6, -20, 28, 13, -16, 1, -1, -15,
    -- layer=1 filter=161 channel=106
    -53, -10, 37, -46, 11, 47, -3, 22, 25,
    -- layer=1 filter=161 channel=107
    10, 5, -1, 4, 6, -5, 1, -2, 12,
    -- layer=1 filter=161 channel=108
    -60, 20, 39, -40, 30, 57, -33, 14, 9,
    -- layer=1 filter=161 channel=109
    -4, 0, 7, 2, -10, 0, -9, -3, -4,
    -- layer=1 filter=161 channel=110
    8, -6, -11, -4, -4, -6, 0, 0, 4,
    -- layer=1 filter=161 channel=111
    -3, 0, 35, -21, 13, 21, 25, 18, 16,
    -- layer=1 filter=161 channel=112
    -17, 35, 35, -6, 1, 11, -6, 4, 3,
    -- layer=1 filter=161 channel=113
    -46, -15, -2, -21, -18, 31, -8, -28, 15,
    -- layer=1 filter=161 channel=114
    40, 20, -36, -11, -39, 23, 9, -26, -28,
    -- layer=1 filter=161 channel=115
    33, 18, -38, 28, 11, -24, 0, -15, -44,
    -- layer=1 filter=161 channel=116
    0, 2, 0, 5, -8, -6, -1, -11, 0,
    -- layer=1 filter=161 channel=117
    -21, 2, 7, -34, -42, -12, -40, -35, -19,
    -- layer=1 filter=161 channel=118
    -27, -11, 55, -48, 22, 33, 27, 6, 22,
    -- layer=1 filter=161 channel=119
    -39, -4, 42, -15, 31, 54, 10, 9, 24,
    -- layer=1 filter=161 channel=120
    10, -11, -27, -3, -15, -8, 8, -16, 0,
    -- layer=1 filter=161 channel=121
    -7, -22, -55, -7, -9, -25, -19, -32, -19,
    -- layer=1 filter=161 channel=122
    6, -6, 6, 6, 10, 8, 4, 10, -1,
    -- layer=1 filter=161 channel=123
    31, 3, -19, 20, 4, -4, 27, -27, 6,
    -- layer=1 filter=161 channel=124
    0, -19, -2, -15, 2, -14, -1, -7, -15,
    -- layer=1 filter=161 channel=125
    -50, -26, 9, -51, -57, 31, -39, -13, 54,
    -- layer=1 filter=161 channel=126
    23, 21, -29, 6, -19, -27, -40, -74, 12,
    -- layer=1 filter=161 channel=127
    -17, 11, 48, -17, 14, 10, 13, 3, 9,
    -- layer=1 filter=162 channel=0
    36, -23, -39, 15, -22, -33, -24, -36, -23,
    -- layer=1 filter=162 channel=1
    24, -69, -65, -49, -80, -64, -54, -86, -14,
    -- layer=1 filter=162 channel=2
    0, 16, 35, 13, 31, 30, 31, 24, 33,
    -- layer=1 filter=162 channel=3
    -6, 7, 6, -10, 3, 4, -5, 9, -4,
    -- layer=1 filter=162 channel=4
    8, -16, -9, 3, 1, -2, -8, 3, 3,
    -- layer=1 filter=162 channel=5
    -27, -125, -87, -66, -92, -76, -113, -83, -43,
    -- layer=1 filter=162 channel=6
    -10, -53, -31, -33, -61, -17, -23, -9, -4,
    -- layer=1 filter=162 channel=7
    0, -60, -7, -45, 1, 1, 28, -16, 31,
    -- layer=1 filter=162 channel=8
    -9, -127, -59, -68, -91, -66, -89, -64, -18,
    -- layer=1 filter=162 channel=9
    75, 97, -5, 92, 42, -6, -15, -15, -2,
    -- layer=1 filter=162 channel=10
    -9, -52, -7, -31, 2, 13, 16, -22, 29,
    -- layer=1 filter=162 channel=11
    58, 17, -32, 36, -7, -6, 38, -6, -1,
    -- layer=1 filter=162 channel=12
    -14, -43, -13, 4, -59, -62, -7, 8, 22,
    -- layer=1 filter=162 channel=13
    35, 34, 8, 34, 2, 4, 36, 5, 16,
    -- layer=1 filter=162 channel=14
    7, -94, -20, -27, -6, -20, -15, -26, 0,
    -- layer=1 filter=162 channel=15
    -34, 29, -29, 9, -10, 10, 4, 23, 1,
    -- layer=1 filter=162 channel=16
    -70, -120, -28, -83, -93, -49, -83, -75, -44,
    -- layer=1 filter=162 channel=17
    32, 4, -37, 8, -25, -15, 15, -32, -27,
    -- layer=1 filter=162 channel=18
    70, -11, -79, 27, -52, -102, -44, -52, -13,
    -- layer=1 filter=162 channel=19
    30, 47, -38, 67, 14, -67, -11, -32, -48,
    -- layer=1 filter=162 channel=20
    -15, -30, 28, -18, -17, -3, -5, -25, 4,
    -- layer=1 filter=162 channel=21
    -21, -25, 35, -27, 14, 25, 6, -13, 7,
    -- layer=1 filter=162 channel=22
    6, -76, -12, -34, -66, -13, 6, -18, 14,
    -- layer=1 filter=162 channel=23
    -4, 8, -33, -32, -19, -12, -9, 42, -5,
    -- layer=1 filter=162 channel=24
    -4, 63, 26, 33, 19, 8, 17, -7, -14,
    -- layer=1 filter=162 channel=25
    51, -28, 4, -10, -24, 17, 4, -19, 36,
    -- layer=1 filter=162 channel=26
    61, 91, 0, 63, -6, -54, 49, -47, -53,
    -- layer=1 filter=162 channel=27
    11, 6, 35, -1, 11, 18, 2, 14, 7,
    -- layer=1 filter=162 channel=28
    27, -66, -13, -8, -1, -10, -2, -65, 13,
    -- layer=1 filter=162 channel=29
    -40, -76, -37, -47, -46, -56, -45, -51, -45,
    -- layer=1 filter=162 channel=30
    51, 32, -128, 71, -26, -147, -37, -105, -67,
    -- layer=1 filter=162 channel=31
    32, -52, -24, 35, -6, -18, 0, 4, 33,
    -- layer=1 filter=162 channel=32
    69, 89, -19, 67, 0, -77, 42, -48, -55,
    -- layer=1 filter=162 channel=33
    -9, 0, 23, 7, -20, -4, -27, -36, -21,
    -- layer=1 filter=162 channel=34
    10, -2, -5, 3, 0, 15, -18, -23, 6,
    -- layer=1 filter=162 channel=35
    7, 3, -15, 6, -2, -7, 10, 3, 6,
    -- layer=1 filter=162 channel=36
    48, 14, -10, 27, 3, 4, 14, 0, 1,
    -- layer=1 filter=162 channel=37
    -59, -72, -38, -42, -76, -45, -80, -52, -56,
    -- layer=1 filter=162 channel=38
    -11, -8, 18, 19, -1, 15, 4, 1, 17,
    -- layer=1 filter=162 channel=39
    -17, -22, -26, -28, -9, -33, -16, -18, -16,
    -- layer=1 filter=162 channel=40
    -8, -74, -80, -31, -64, -38, -42, -26, 21,
    -- layer=1 filter=162 channel=41
    96, 145, -55, 108, 35, -25, 70, -20, -52,
    -- layer=1 filter=162 channel=42
    -13, 12, 33, 30, 31, 43, 19, 28, 32,
    -- layer=1 filter=162 channel=43
    8, -48, -34, -88, -93, -15, -40, -39, 0,
    -- layer=1 filter=162 channel=44
    62, 55, -22, 52, -31, -81, 49, -43, -27,
    -- layer=1 filter=162 channel=45
    -37, 9, 5, -5, -13, -2, -5, -19, -3,
    -- layer=1 filter=162 channel=46
    2, -34, -40, 35, -23, -48, -36, 2, -44,
    -- layer=1 filter=162 channel=47
    36, 62, -15, 44, -11, 17, 28, 2, -2,
    -- layer=1 filter=162 channel=48
    -64, -17, -12, -55, -9, 16, -40, -17, 5,
    -- layer=1 filter=162 channel=49
    -13, 16, 10, 4, 15, 27, -14, 20, 23,
    -- layer=1 filter=162 channel=50
    0, -5, 2, 22, -28, -7, -25, -9, 2,
    -- layer=1 filter=162 channel=51
    -13, -25, 2, -22, -1, 16, 32, -13, 41,
    -- layer=1 filter=162 channel=52
    -13, 13, -3, -10, -31, -45, 1, 0, -12,
    -- layer=1 filter=162 channel=53
    11, 4, 2, -2, -20, -10, -8, -15, -5,
    -- layer=1 filter=162 channel=54
    40, 23, 4, 25, -14, 33, 0, -7, 37,
    -- layer=1 filter=162 channel=55
    30, 26, 17, 34, 11, 24, 35, 16, -1,
    -- layer=1 filter=162 channel=56
    3, 7, 3, -2, -9, 1, -8, -5, 8,
    -- layer=1 filter=162 channel=57
    8, -56, 8, -6, -5, 24, -5, -19, 45,
    -- layer=1 filter=162 channel=58
    -27, -7, -5, -19, 17, 46, -58, 26, 36,
    -- layer=1 filter=162 channel=59
    -2, -2, -6, 3, 8, -12, -1, -3, 4,
    -- layer=1 filter=162 channel=60
    15, -23, 17, -26, 13, -4, -23, 9, -9,
    -- layer=1 filter=162 channel=61
    0, -10, -8, 6, -12, -6, 0, -5, -6,
    -- layer=1 filter=162 channel=62
    -55, -126, -47, -128, -91, -57, -107, -55, -35,
    -- layer=1 filter=162 channel=63
    51, 13, -43, 45, -17, -23, 29, -4, -23,
    -- layer=1 filter=162 channel=64
    35, -54, -27, -20, -26, -1, -35, -68, 13,
    -- layer=1 filter=162 channel=65
    -45, -26, -9, -45, 6, -6, -19, -24, -8,
    -- layer=1 filter=162 channel=66
    26, -11, -21, -2, 13, -16, -4, -9, -10,
    -- layer=1 filter=162 channel=67
    -14, -56, -46, -43, -26, -32, -31, -36, -19,
    -- layer=1 filter=162 channel=68
    60, 46, -57, 52, -64, -79, 41, -47, -45,
    -- layer=1 filter=162 channel=69
    -29, -8, -22, -14, -38, -61, -15, -34, -56,
    -- layer=1 filter=162 channel=70
    -6, -28, -16, -42, -76, -25, -87, -52, 23,
    -- layer=1 filter=162 channel=71
    -58, -1, 8, -30, 19, -7, -20, 6, 9,
    -- layer=1 filter=162 channel=72
    52, 49, -57, 67, -10, -103, -40, -58, -78,
    -- layer=1 filter=162 channel=73
    -11, -5, 0, -12, -11, 0, -2, -10, -7,
    -- layer=1 filter=162 channel=74
    66, -16, -88, 49, -93, -89, 5, -35, -32,
    -- layer=1 filter=162 channel=75
    4, -75, -69, -10, -55, -98, -52, 1, 33,
    -- layer=1 filter=162 channel=76
    63, 62, -32, 57, -7, -16, 47, -43, -53,
    -- layer=1 filter=162 channel=77
    -56, -20, -24, -31, -11, -5, -23, -22, -23,
    -- layer=1 filter=162 channel=78
    4, -21, -24, -32, -21, -39, 2, -27, -8,
    -- layer=1 filter=162 channel=79
    -61, -104, -28, -80, -74, -36, -102, -42, -30,
    -- layer=1 filter=162 channel=80
    9, -32, 0, -6, 5, 16, 26, -10, -3,
    -- layer=1 filter=162 channel=81
    -66, -1, 19, -30, 7, 8, -23, 3, -10,
    -- layer=1 filter=162 channel=82
    -36, -8, 5, -32, 6, 14, 0, 15, 9,
    -- layer=1 filter=162 channel=83
    -19, -5, -61, -3, -77, -35, -9, -60, -26,
    -- layer=1 filter=162 channel=84
    104, 65, -115, 56, -59, -116, 34, -46, -84,
    -- layer=1 filter=162 channel=85
    40, 51, -39, 38, 2, 4, -16, 11, 19,
    -- layer=1 filter=162 channel=86
    28, -25, -25, 21, -4, -7, 22, -9, 6,
    -- layer=1 filter=162 channel=87
    71, 32, -18, 88, 44, -32, -49, -27, -45,
    -- layer=1 filter=162 channel=88
    -30, -8, 20, -16, -9, 5, -16, 1, -13,
    -- layer=1 filter=162 channel=89
    4, -12, -10, -22, 1, -24, -17, 2, -11,
    -- layer=1 filter=162 channel=90
    28, 54, -14, 56, -27, -69, 41, -45, -36,
    -- layer=1 filter=162 channel=91
    9, -32, -18, -28, -13, 23, -4, -1, 28,
    -- layer=1 filter=162 channel=92
    27, 57, -9, 36, -17, -9, 53, -39, 30,
    -- layer=1 filter=162 channel=93
    -12, -15, 8, -17, 0, 21, -23, -3, 8,
    -- layer=1 filter=162 channel=94
    54, -37, -68, 2, -9, -35, -12, -33, -9,
    -- layer=1 filter=162 channel=95
    82, 7, -120, 43, -75, -150, -13, -50, -70,
    -- layer=1 filter=162 channel=96
    18, 21, 45, 1, -27, -2, 7, -6, -6,
    -- layer=1 filter=162 channel=97
    30, -26, -16, -7, -11, -15, -13, -40, -4,
    -- layer=1 filter=162 channel=98
    -4, -101, -20, -108, -78, 0, -67, -47, -13,
    -- layer=1 filter=162 channel=99
    -9, -86, -45, -75, -60, -40, -24, -118, -22,
    -- layer=1 filter=162 channel=100
    65, 12, -18, 50, -23, -9, 15, -4, -13,
    -- layer=1 filter=162 channel=101
    10, -20, -2, -19, -14, 11, 7, 9, 31,
    -- layer=1 filter=162 channel=102
    45, -14, -69, 22, -52, -27, 3, -43, -2,
    -- layer=1 filter=162 channel=103
    37, 27, -8, 31, 29, -8, 23, -8, -4,
    -- layer=1 filter=162 channel=104
    34, 73, -27, 30, 31, -34, 27, 15, 12,
    -- layer=1 filter=162 channel=105
    14, -42, -43, -32, -5, 8, -32, -29, 10,
    -- layer=1 filter=162 channel=106
    42, 66, -13, 26, -18, -16, 40, -8, -2,
    -- layer=1 filter=162 channel=107
    10, -11, -12, -2, -4, 4, 8, -4, 5,
    -- layer=1 filter=162 channel=108
    44, 92, -17, 57, 14, -72, 34, -25, -50,
    -- layer=1 filter=162 channel=109
    7, -2, 0, 1, -8, 0, -4, 4, 10,
    -- layer=1 filter=162 channel=110
    -1, -9, -28, -8, 13, -18, -3, 9, -23,
    -- layer=1 filter=162 channel=111
    55, -14, -137, 16, -84, -144, -44, -76, -61,
    -- layer=1 filter=162 channel=112
    61, -3, -87, -46, -83, -66, -12, 5, -30,
    -- layer=1 filter=162 channel=113
    -1, -16, 60, 35, -1, 41, 30, 5, 39,
    -- layer=1 filter=162 channel=114
    -73, -61, -47, -44, -57, -35, -89, -59, -34,
    -- layer=1 filter=162 channel=115
    -2, -33, -38, -44, -13, -2, -51, -6, 18,
    -- layer=1 filter=162 channel=116
    0, -8, 2, -7, 8, 4, 7, -8, 8,
    -- layer=1 filter=162 channel=117
    22, -56, -81, -99, -47, -63, -21, -31, -14,
    -- layer=1 filter=162 channel=118
    67, 45, -102, 59, -37, -126, 4, -75, -37,
    -- layer=1 filter=162 channel=119
    45, 101, -38, 49, -13, -72, 41, -52, -80,
    -- layer=1 filter=162 channel=120
    -27, -26, 29, -23, 15, 52, 5, 6, 35,
    -- layer=1 filter=162 channel=121
    9, -27, -43, 51, 10, -32, -25, 3, -1,
    -- layer=1 filter=162 channel=122
    0, -7, 9, -6, 3, 6, 2, 1, -5,
    -- layer=1 filter=162 channel=123
    8, -8, -25, 7, 17, -15, -24, 14, -12,
    -- layer=1 filter=162 channel=124
    2, 5, 0, 2, -9, -1, -12, -19, -12,
    -- layer=1 filter=162 channel=125
    39, -25, 24, 21, -68, 27, 29, -45, 10,
    -- layer=1 filter=162 channel=126
    -38, -117, -103, -110, -148, -54, -66, -58, -64,
    -- layer=1 filter=162 channel=127
    74, 11, -131, 50, -73, -163, -14, -72, -55,
    -- layer=1 filter=163 channel=0
    5, 1, 2, -10, 0, 7, -9, -10, -10,
    -- layer=1 filter=163 channel=1
    6, -4, -5, 3, -9, 8, 0, -9, 0,
    -- layer=1 filter=163 channel=2
    -15, 0, -4, -1, -14, -9, -13, 6, -10,
    -- layer=1 filter=163 channel=3
    5, 4, 8, -9, 2, 1, -4, 9, -8,
    -- layer=1 filter=163 channel=4
    8, 7, 7, -5, -7, -7, 1, 4, 1,
    -- layer=1 filter=163 channel=5
    3, 3, -9, -11, 3, -10, -10, -8, -8,
    -- layer=1 filter=163 channel=6
    2, 3, 0, 8, 0, -11, 1, 4, 7,
    -- layer=1 filter=163 channel=7
    -7, 0, 0, 0, 5, -8, -11, 0, -6,
    -- layer=1 filter=163 channel=8
    -4, -2, -3, 1, -4, -8, -10, -1, -8,
    -- layer=1 filter=163 channel=9
    -3, 8, 2, -1, -11, 7, 9, -4, 0,
    -- layer=1 filter=163 channel=10
    2, 0, -5, -1, 3, -6, 0, 2, -7,
    -- layer=1 filter=163 channel=11
    -11, 0, 1, -4, 5, -1, 3, 3, -7,
    -- layer=1 filter=163 channel=12
    -9, 0, 0, 9, -1, 0, -4, -8, 5,
    -- layer=1 filter=163 channel=13
    -9, -4, -2, -1, 7, 1, -1, 4, 6,
    -- layer=1 filter=163 channel=14
    -7, -9, 1, -6, -12, 4, -10, 4, -9,
    -- layer=1 filter=163 channel=15
    -6, -10, 1, -5, -4, -2, -11, 1, 12,
    -- layer=1 filter=163 channel=16
    1, -5, -5, -7, -7, -5, -7, -9, 0,
    -- layer=1 filter=163 channel=17
    8, -5, -10, 6, 8, -9, -5, -7, 1,
    -- layer=1 filter=163 channel=18
    10, -5, 4, 4, -5, -10, 2, 0, 4,
    -- layer=1 filter=163 channel=19
    3, 3, -11, -3, -6, -10, 9, -1, -9,
    -- layer=1 filter=163 channel=20
    -7, -6, -7, 0, 1, -5, 4, -1, 5,
    -- layer=1 filter=163 channel=21
    3, -7, 5, -11, 3, -7, -6, 6, 11,
    -- layer=1 filter=163 channel=22
    0, 1, -5, 2, 4, -3, -10, -1, 9,
    -- layer=1 filter=163 channel=23
    -6, 8, 7, 0, -1, -10, -1, -3, -11,
    -- layer=1 filter=163 channel=24
    -8, 7, -1, 3, 0, -7, -3, 2, -4,
    -- layer=1 filter=163 channel=25
    -5, 1, -11, 0, 7, 5, 3, -2, 2,
    -- layer=1 filter=163 channel=26
    -6, 3, -7, 5, 4, 4, -5, -6, -7,
    -- layer=1 filter=163 channel=27
    5, 9, 0, 0, -2, 7, -9, -2, -8,
    -- layer=1 filter=163 channel=28
    1, 7, -4, 3, 7, -7, -4, -12, 0,
    -- layer=1 filter=163 channel=29
    11, 0, 4, -6, -10, 0, 4, 7, -4,
    -- layer=1 filter=163 channel=30
    -7, 4, -12, 4, -5, -7, 0, -4, 5,
    -- layer=1 filter=163 channel=31
    0, 0, 3, -1, 8, -2, 6, 4, -7,
    -- layer=1 filter=163 channel=32
    -10, 3, -8, 7, 5, -3, 6, 7, 6,
    -- layer=1 filter=163 channel=33
    7, 8, 4, 6, -5, -2, 1, 9, -8,
    -- layer=1 filter=163 channel=34
    2, -8, -4, -2, 4, -3, 0, 1, -8,
    -- layer=1 filter=163 channel=35
    -9, -2, -11, 0, 10, -5, 7, 9, 6,
    -- layer=1 filter=163 channel=36
    -4, 0, -4, 6, 3, -3, -8, -5, -3,
    -- layer=1 filter=163 channel=37
    -5, -5, -1, 5, 4, -9, -8, -1, -13,
    -- layer=1 filter=163 channel=38
    6, -3, 0, -10, -3, 1, 3, -8, 3,
    -- layer=1 filter=163 channel=39
    -11, -3, 1, -5, 6, -2, -7, 3, 0,
    -- layer=1 filter=163 channel=40
    -4, -4, -1, 8, 0, 0, 5, 6, -4,
    -- layer=1 filter=163 channel=41
    7, -4, -5, -7, -1, -3, -8, -3, -11,
    -- layer=1 filter=163 channel=42
    -10, -8, 0, -10, 5, -13, -2, -3, -7,
    -- layer=1 filter=163 channel=43
    -10, -2, -9, -10, -6, -10, 2, -1, -9,
    -- layer=1 filter=163 channel=44
    -3, 3, 8, -8, 8, -11, -10, 1, 4,
    -- layer=1 filter=163 channel=45
    -6, 5, -2, 0, -9, -4, -6, 2, -10,
    -- layer=1 filter=163 channel=46
    7, -6, 3, 2, -5, -7, -11, -6, 2,
    -- layer=1 filter=163 channel=47
    -3, -8, 3, 8, -4, -11, -1, 10, 1,
    -- layer=1 filter=163 channel=48
    -6, -7, 6, -8, -8, -7, -3, 8, 6,
    -- layer=1 filter=163 channel=49
    0, -11, 7, -6, 7, -3, 6, -1, 0,
    -- layer=1 filter=163 channel=50
    4, -9, -3, 2, 8, 4, 2, 2, -1,
    -- layer=1 filter=163 channel=51
    0, -8, -3, 4, 3, 7, 0, 0, 5,
    -- layer=1 filter=163 channel=52
    -5, 0, -2, -1, -8, 1, 4, 0, 3,
    -- layer=1 filter=163 channel=53
    5, 7, -6, 4, 0, 3, -1, -6, 4,
    -- layer=1 filter=163 channel=54
    -9, 1, -4, 4, 1, 8, -9, 0, -2,
    -- layer=1 filter=163 channel=55
    0, 0, -10, -10, 7, 5, -7, -3, -13,
    -- layer=1 filter=163 channel=56
    7, -5, -5, 3, -5, -9, 7, 1, 4,
    -- layer=1 filter=163 channel=57
    -11, -1, 3, -11, -1, 8, -7, 5, -9,
    -- layer=1 filter=163 channel=58
    0, -2, -4, 0, -11, 10, -10, 8, -9,
    -- layer=1 filter=163 channel=59
    0, 8, -9, 3, 0, -9, -11, 3, -6,
    -- layer=1 filter=163 channel=60
    -4, -8, 0, 2, 1, 4, 0, 0, -5,
    -- layer=1 filter=163 channel=61
    9, -2, 7, -7, -4, -9, -7, -4, -3,
    -- layer=1 filter=163 channel=62
    7, -1, 7, -11, 3, 7, -11, 1, 2,
    -- layer=1 filter=163 channel=63
    4, -9, -8, -10, -2, -7, -1, -2, -8,
    -- layer=1 filter=163 channel=64
    -9, -5, 3, -5, -1, -11, 6, 7, 1,
    -- layer=1 filter=163 channel=65
    -9, 2, 6, -8, 6, 8, 9, -10, -5,
    -- layer=1 filter=163 channel=66
    2, -8, 6, 8, 5, 5, -12, -9, -12,
    -- layer=1 filter=163 channel=67
    1, -1, -1, -3, -6, -10, -4, -1, -2,
    -- layer=1 filter=163 channel=68
    -10, -1, 0, 5, 6, -1, -1, -11, 12,
    -- layer=1 filter=163 channel=69
    -6, -7, -6, -12, 0, -3, -1, -6, -7,
    -- layer=1 filter=163 channel=70
    0, 4, 5, 6, 3, -9, -3, -2, 6,
    -- layer=1 filter=163 channel=71
    3, -9, 5, -2, -2, 2, -9, -11, 6,
    -- layer=1 filter=163 channel=72
    -12, 7, -6, 4, 8, -4, -10, 0, 9,
    -- layer=1 filter=163 channel=73
    1, -8, -8, 8, 5, -3, 2, -3, 7,
    -- layer=1 filter=163 channel=74
    -5, -8, 0, 0, 0, 3, 1, 0, 4,
    -- layer=1 filter=163 channel=75
    -1, -5, -2, 4, -3, 5, 3, 10, 0,
    -- layer=1 filter=163 channel=76
    1, 1, 3, 2, 1, 8, -9, -1, 0,
    -- layer=1 filter=163 channel=77
    -1, -11, 0, 4, -5, 7, -4, -8, -11,
    -- layer=1 filter=163 channel=78
    -3, -8, 0, 3, -4, 8, 4, -9, -1,
    -- layer=1 filter=163 channel=79
    -5, 8, 0, 8, -7, 2, -12, 2, -16,
    -- layer=1 filter=163 channel=80
    9, 4, 1, -5, 8, -9, -3, -4, -6,
    -- layer=1 filter=163 channel=81
    -4, -10, -9, -11, 4, 0, 0, 7, 0,
    -- layer=1 filter=163 channel=82
    0, -6, 4, -10, 3, -5, 5, 0, -7,
    -- layer=1 filter=163 channel=83
    5, -10, -4, 6, -2, -4, 4, -4, 6,
    -- layer=1 filter=163 channel=84
    -8, -10, 0, -9, -8, -5, 2, -10, -4,
    -- layer=1 filter=163 channel=85
    -5, -4, -11, -10, 3, -8, -2, -2, -9,
    -- layer=1 filter=163 channel=86
    4, -1, 7, 0, 7, 5, -3, 6, -8,
    -- layer=1 filter=163 channel=87
    -3, -7, -1, -4, 6, 0, -11, 9, 0,
    -- layer=1 filter=163 channel=88
    4, 0, -4, -2, -4, 0, -9, 2, -7,
    -- layer=1 filter=163 channel=89
    -2, 2, -11, -10, -4, -5, 6, -5, -4,
    -- layer=1 filter=163 channel=90
    -4, -2, -7, 4, -11, 1, -1, 7, -9,
    -- layer=1 filter=163 channel=91
    4, -12, 6, 2, 0, 0, -10, -9, -7,
    -- layer=1 filter=163 channel=92
    0, 8, 5, -1, 4, 0, 0, -10, -2,
    -- layer=1 filter=163 channel=93
    -10, -1, 3, -2, 0, 2, -9, 7, -11,
    -- layer=1 filter=163 channel=94
    -8, 0, -10, -3, -10, -5, 5, 4, -4,
    -- layer=1 filter=163 channel=95
    -4, 2, -3, -7, 2, 6, -5, 1, -11,
    -- layer=1 filter=163 channel=96
    6, 6, -9, 0, 7, -4, -8, 8, 6,
    -- layer=1 filter=163 channel=97
    1, -3, 6, -10, 5, 0, 0, -3, 8,
    -- layer=1 filter=163 channel=98
    -12, -11, 3, -6, -13, -4, 6, -4, -6,
    -- layer=1 filter=163 channel=99
    4, -7, 0, 0, 2, 4, 3, 6, 6,
    -- layer=1 filter=163 channel=100
    7, 0, 3, -10, 0, -6, 4, -5, -9,
    -- layer=1 filter=163 channel=101
    5, -10, -5, 6, -11, 6, -2, -9, -10,
    -- layer=1 filter=163 channel=102
    3, 3, -1, -4, 7, 0, 7, -2, 5,
    -- layer=1 filter=163 channel=103
    -6, -8, -3, 6, -2, 3, 4, -7, -6,
    -- layer=1 filter=163 channel=104
    -4, -9, 4, -1, -8, 6, 1, -3, 0,
    -- layer=1 filter=163 channel=105
    4, -5, 2, -6, -8, -6, -10, -9, -6,
    -- layer=1 filter=163 channel=106
    0, -7, 3, -4, -6, 2, -4, -10, -5,
    -- layer=1 filter=163 channel=107
    5, -1, -7, -7, -8, -8, 4, -8, 9,
    -- layer=1 filter=163 channel=108
    4, -9, 3, -11, -1, -7, 0, 7, -2,
    -- layer=1 filter=163 channel=109
    -3, 0, 9, -1, 5, 0, 6, 0, -6,
    -- layer=1 filter=163 channel=110
    -1, -1, -2, 0, -10, 5, -7, -10, 7,
    -- layer=1 filter=163 channel=111
    -5, 7, 7, -6, 0, 7, -3, 8, 1,
    -- layer=1 filter=163 channel=112
    0, -11, 0, 0, 4, -11, -11, -6, -6,
    -- layer=1 filter=163 channel=113
    3, 5, -6, -5, 9, -4, 7, 3, -5,
    -- layer=1 filter=163 channel=114
    1, 4, 5, 0, 4, -3, -7, -4, 0,
    -- layer=1 filter=163 channel=115
    -4, 5, -2, 3, -12, 0, 8, -6, -5,
    -- layer=1 filter=163 channel=116
    3, 6, -6, -4, -2, -7, 8, -1, 10,
    -- layer=1 filter=163 channel=117
    -2, 9, 1, -4, -3, 5, -8, 0, -2,
    -- layer=1 filter=163 channel=118
    -9, 4, -7, -4, -7, -11, -6, 3, -6,
    -- layer=1 filter=163 channel=119
    -2, 4, 4, 8, -10, -8, -1, 4, 4,
    -- layer=1 filter=163 channel=120
    -4, 2, -1, -10, -5, -12, -11, 4, 5,
    -- layer=1 filter=163 channel=121
    6, -2, 5, 5, 0, 0, -8, -6, -9,
    -- layer=1 filter=163 channel=122
    -7, -4, 0, -8, -1, 4, 0, -3, 9,
    -- layer=1 filter=163 channel=123
    -9, -6, 0, 2, -1, -1, -8, -7, -1,
    -- layer=1 filter=163 channel=124
    1, 5, 8, 0, 9, 1, -4, 7, -5,
    -- layer=1 filter=163 channel=125
    6, -5, 4, -10, 9, 4, -1, 0, 0,
    -- layer=1 filter=163 channel=126
    5, 2, 6, 1, 3, 7, 1, 2, -10,
    -- layer=1 filter=163 channel=127
    11, 10, -1, 0, -9, 1, -10, 7, 0,
    -- layer=1 filter=164 channel=0
    -7, 6, -4, 6, 1, -3, -11, 3, 6,
    -- layer=1 filter=164 channel=1
    -10, -3, -6, 7, 1, 8, 1, 5, 2,
    -- layer=1 filter=164 channel=2
    -1, -5, -5, -3, 0, 6, 3, 10, 11,
    -- layer=1 filter=164 channel=3
    9, -10, -2, 5, 0, 9, -6, -2, 5,
    -- layer=1 filter=164 channel=4
    -1, -1, -6, 4, 5, 0, -7, 5, 6,
    -- layer=1 filter=164 channel=5
    -2, 0, 0, -11, 7, 1, 2, 2, 2,
    -- layer=1 filter=164 channel=6
    2, -4, 0, -6, 7, 4, 0, -2, 0,
    -- layer=1 filter=164 channel=7
    -5, 4, -3, -1, -21, -7, -15, 5, -7,
    -- layer=1 filter=164 channel=8
    -3, -5, 6, -6, 3, 8, -6, -11, 8,
    -- layer=1 filter=164 channel=9
    -3, -9, -13, -2, 6, 8, -8, 10, 0,
    -- layer=1 filter=164 channel=10
    5, -7, -7, -12, -14, 0, -5, 3, -15,
    -- layer=1 filter=164 channel=11
    -8, -3, 5, -5, 2, 0, 8, 3, -6,
    -- layer=1 filter=164 channel=12
    -8, -2, 4, -10, -8, 9, -2, -5, 1,
    -- layer=1 filter=164 channel=13
    0, 4, 5, -3, -9, 0, -1, -2, 6,
    -- layer=1 filter=164 channel=14
    2, -8, 4, -7, 1, -10, -8, -11, 0,
    -- layer=1 filter=164 channel=15
    -9, 0, 0, -8, -11, 0, 2, 1, 3,
    -- layer=1 filter=164 channel=16
    3, 0, -1, -1, -8, 0, 1, -12, -2,
    -- layer=1 filter=164 channel=17
    2, -3, -5, 3, 9, 3, -7, 8, -1,
    -- layer=1 filter=164 channel=18
    0, -5, 2, 6, 5, -5, -5, -6, -5,
    -- layer=1 filter=164 channel=19
    0, -2, -2, -10, 6, 6, -1, -7, -7,
    -- layer=1 filter=164 channel=20
    -1, -8, 2, -5, 3, -7, 3, -12, 0,
    -- layer=1 filter=164 channel=21
    2, -10, -3, -4, -3, -10, -1, -5, -4,
    -- layer=1 filter=164 channel=22
    -3, -6, -10, 0, 0, -3, -10, 6, 1,
    -- layer=1 filter=164 channel=23
    -10, 0, 6, 5, -11, 0, -2, -10, -1,
    -- layer=1 filter=164 channel=24
    -9, 0, -1, 0, -6, 7, 3, -12, 0,
    -- layer=1 filter=164 channel=25
    -3, -8, 3, 0, -11, 3, 2, -4, -7,
    -- layer=1 filter=164 channel=26
    0, -6, -13, 3, 1, 10, 7, 1, 0,
    -- layer=1 filter=164 channel=27
    3, -10, 4, 2, -7, 2, 0, 6, -2,
    -- layer=1 filter=164 channel=28
    -5, -10, 8, -6, -10, 6, -8, 3, 6,
    -- layer=1 filter=164 channel=29
    1, 4, -4, -8, 0, 5, -1, -5, 0,
    -- layer=1 filter=164 channel=30
    -11, -10, 1, -14, -6, 6, 0, -3, 1,
    -- layer=1 filter=164 channel=31
    -10, -4, 0, -7, -8, -1, 10, 0, -7,
    -- layer=1 filter=164 channel=32
    -2, -9, -5, -8, 4, -2, -7, -1, -11,
    -- layer=1 filter=164 channel=33
    -5, 0, -12, 6, 5, 2, -1, 3, -7,
    -- layer=1 filter=164 channel=34
    4, -9, -8, -2, -3, 1, 3, 8, -10,
    -- layer=1 filter=164 channel=35
    2, -2, 8, 7, 6, -11, 8, -9, -12,
    -- layer=1 filter=164 channel=36
    -8, -4, 6, 3, 1, -10, -11, -2, 3,
    -- layer=1 filter=164 channel=37
    4, -1, -11, -1, -8, -3, -8, -11, 1,
    -- layer=1 filter=164 channel=38
    0, 2, 6, -2, -3, -1, -8, -7, 0,
    -- layer=1 filter=164 channel=39
    -9, 4, 3, 1, -6, 6, -2, 5, -7,
    -- layer=1 filter=164 channel=40
    -10, 1, 2, -10, -4, -9, 1, 3, -5,
    -- layer=1 filter=164 channel=41
    -2, -1, 4, -3, -2, 5, -10, -7, -1,
    -- layer=1 filter=164 channel=42
    3, -10, -10, -2, 8, -5, 0, -6, -4,
    -- layer=1 filter=164 channel=43
    4, 4, 4, -2, 6, 4, 0, 0, 9,
    -- layer=1 filter=164 channel=44
    0, 9, 3, -5, -11, -10, -4, -2, 2,
    -- layer=1 filter=164 channel=45
    1, 4, 0, 0, 4, -3, 5, 4, 5,
    -- layer=1 filter=164 channel=46
    -7, -8, -7, -2, 3, 1, -11, 4, 7,
    -- layer=1 filter=164 channel=47
    -12, -9, 0, -6, -13, 2, -2, -6, 0,
    -- layer=1 filter=164 channel=48
    6, -1, -7, 2, -2, 4, -1, 2, -7,
    -- layer=1 filter=164 channel=49
    -9, -1, -3, -7, 2, 4, -3, -6, -8,
    -- layer=1 filter=164 channel=50
    -1, 0, -12, 4, -6, 5, 0, -10, 2,
    -- layer=1 filter=164 channel=51
    4, -6, 4, 0, 2, 5, 4, 1, -13,
    -- layer=1 filter=164 channel=52
    8, 10, 10, 8, 3, -7, 1, -10, 7,
    -- layer=1 filter=164 channel=53
    2, 5, 4, -10, 0, -10, 5, 7, -10,
    -- layer=1 filter=164 channel=54
    0, 2, 6, -9, -4, -4, -5, -10, -6,
    -- layer=1 filter=164 channel=55
    -1, 0, 1, 0, -6, -7, 8, 0, -12,
    -- layer=1 filter=164 channel=56
    2, 4, 0, -3, -3, -10, -1, 2, -2,
    -- layer=1 filter=164 channel=57
    4, -1, 1, -8, 7, 0, 9, 4, 6,
    -- layer=1 filter=164 channel=58
    0, -7, -5, -4, -3, 0, -12, -4, 6,
    -- layer=1 filter=164 channel=59
    -5, -6, -6, 7, -7, -7, 0, -8, -8,
    -- layer=1 filter=164 channel=60
    6, -8, 0, -1, -7, -3, 2, 7, -3,
    -- layer=1 filter=164 channel=61
    8, -9, 7, 0, 6, 9, -3, 11, 9,
    -- layer=1 filter=164 channel=62
    2, -7, 7, 4, 0, 3, -3, -12, -5,
    -- layer=1 filter=164 channel=63
    -6, -7, -3, -8, 5, 7, 5, -3, 4,
    -- layer=1 filter=164 channel=64
    8, -7, 1, 6, -8, 0, -6, 6, 0,
    -- layer=1 filter=164 channel=65
    0, -8, -8, -5, -6, -3, -1, -2, 0,
    -- layer=1 filter=164 channel=66
    -9, 2, -12, -9, 1, -3, -9, 8, -9,
    -- layer=1 filter=164 channel=67
    -7, 9, 4, -9, -4, -9, 10, 6, -3,
    -- layer=1 filter=164 channel=68
    -7, -8, 1, 7, -9, -3, 0, 0, 2,
    -- layer=1 filter=164 channel=69
    -9, -6, -6, -4, 0, 1, 13, -11, 8,
    -- layer=1 filter=164 channel=70
    -3, 2, -12, -2, -14, -19, -9, 2, -1,
    -- layer=1 filter=164 channel=71
    4, -9, 3, -1, 4, 1, 0, 5, -1,
    -- layer=1 filter=164 channel=72
    4, -9, 0, -12, 2, 3, -3, -9, 8,
    -- layer=1 filter=164 channel=73
    9, -5, -5, 6, 4, -4, -1, -11, 5,
    -- layer=1 filter=164 channel=74
    -5, -12, -4, -3, 4, 8, -7, -2, 1,
    -- layer=1 filter=164 channel=75
    -15, 5, -1, 7, 2, 6, -3, -5, -13,
    -- layer=1 filter=164 channel=76
    -9, 6, 4, -11, 0, 6, 8, -10, -11,
    -- layer=1 filter=164 channel=77
    -5, -11, -6, -6, -8, -6, 7, -5, -11,
    -- layer=1 filter=164 channel=78
    -6, -7, -3, 0, 3, 2, -7, 1, -3,
    -- layer=1 filter=164 channel=79
    -2, -9, -5, -5, 0, 3, 6, 3, 5,
    -- layer=1 filter=164 channel=80
    0, 2, 4, 7, -6, 4, -7, -4, -6,
    -- layer=1 filter=164 channel=81
    -1, -6, -2, 8, 8, -9, 0, -3, -5,
    -- layer=1 filter=164 channel=82
    -12, -3, 7, 7, -7, -11, -5, -12, 1,
    -- layer=1 filter=164 channel=83
    -7, 2, 2, 6, 4, -11, -11, -2, -10,
    -- layer=1 filter=164 channel=84
    -11, -8, 1, -9, 0, 2, 0, 11, 4,
    -- layer=1 filter=164 channel=85
    7, -6, -7, 1, 6, 5, -10, 3, 0,
    -- layer=1 filter=164 channel=86
    -7, 3, 2, -2, 3, -11, -12, -2, -4,
    -- layer=1 filter=164 channel=87
    4, 6, -11, 6, 3, -10, -6, 9, 8,
    -- layer=1 filter=164 channel=88
    -10, 2, -11, 3, -2, -13, -12, -12, 2,
    -- layer=1 filter=164 channel=89
    -9, -4, 6, -1, -6, 7, 6, 0, -5,
    -- layer=1 filter=164 channel=90
    2, -6, 2, 8, 0, -8, 0, 0, 2,
    -- layer=1 filter=164 channel=91
    -2, 6, 1, -8, 3, -4, -5, -6, -1,
    -- layer=1 filter=164 channel=92
    3, -6, 4, 0, -9, 0, 8, 1, -12,
    -- layer=1 filter=164 channel=93
    -8, 0, 2, -11, -2, -1, 6, -5, 0,
    -- layer=1 filter=164 channel=94
    -10, -11, 5, -7, -5, -3, 1, -4, 6,
    -- layer=1 filter=164 channel=95
    2, 1, -5, -5, -12, 3, 3, -6, 2,
    -- layer=1 filter=164 channel=96
    8, -4, 7, -3, -4, 0, 4, -9, 4,
    -- layer=1 filter=164 channel=97
    -6, 8, 7, 6, -6, 5, -4, -11, 6,
    -- layer=1 filter=164 channel=98
    -9, 2, 3, 4, -7, -9, 0, 1, 0,
    -- layer=1 filter=164 channel=99
    2, -8, -3, -9, -12, 3, -3, 6, 1,
    -- layer=1 filter=164 channel=100
    7, 6, 6, 8, 0, -4, 3, 6, 6,
    -- layer=1 filter=164 channel=101
    -2, -4, -10, 2, -9, 6, -9, 6, 7,
    -- layer=1 filter=164 channel=102
    -8, -7, -1, 0, -7, 6, -5, -8, -6,
    -- layer=1 filter=164 channel=103
    7, 2, -8, 8, 9, -12, 4, 0, 3,
    -- layer=1 filter=164 channel=104
    0, -6, -10, 8, 8, -3, 4, -6, -2,
    -- layer=1 filter=164 channel=105
    2, -5, 6, -4, 6, -6, 7, -6, -2,
    -- layer=1 filter=164 channel=106
    4, 2, 1, 4, -10, -2, 7, -6, 1,
    -- layer=1 filter=164 channel=107
    -2, 10, -5, -6, -8, -9, 0, 8, 0,
    -- layer=1 filter=164 channel=108
    5, -5, -7, -12, -10, 8, 11, 7, -7,
    -- layer=1 filter=164 channel=109
    6, 0, 0, 0, 1, 8, -5, 3, -1,
    -- layer=1 filter=164 channel=110
    -9, 6, -6, -9, 7, -10, -9, 7, 6,
    -- layer=1 filter=164 channel=111
    -12, -1, -9, -2, -1, -13, -8, 1, -6,
    -- layer=1 filter=164 channel=112
    -2, 5, 0, 1, 0, -9, 6, -7, -10,
    -- layer=1 filter=164 channel=113
    -7, 1, 2, -7, -7, -8, 7, 8, 2,
    -- layer=1 filter=164 channel=114
    -6, -10, 3, -10, -15, -17, -10, -8, -14,
    -- layer=1 filter=164 channel=115
    -4, -2, -10, 8, 7, -1, 2, -1, 3,
    -- layer=1 filter=164 channel=116
    -11, -1, -2, -1, -4, -3, 4, 10, 1,
    -- layer=1 filter=164 channel=117
    10, 5, 0, -7, -4, -1, 2, 0, -1,
    -- layer=1 filter=164 channel=118
    -6, -7, -8, 5, 3, 6, -3, -2, -3,
    -- layer=1 filter=164 channel=119
    -9, 7, 7, -5, -3, 6, -2, -4, 5,
    -- layer=1 filter=164 channel=120
    -5, -1, 0, -6, -7, -3, -4, 2, -10,
    -- layer=1 filter=164 channel=121
    7, 0, -4, 3, 6, 1, -6, -11, 2,
    -- layer=1 filter=164 channel=122
    -4, 0, 1, 4, -3, 4, -1, -6, 10,
    -- layer=1 filter=164 channel=123
    -11, -9, 3, 4, 3, 4, 8, 1, -8,
    -- layer=1 filter=164 channel=124
    5, 4, -10, 1, 0, -7, -4, 3, 0,
    -- layer=1 filter=164 channel=125
    -2, -9, -2, 4, 2, -5, -3, -3, -14,
    -- layer=1 filter=164 channel=126
    -1, 2, 2, -9, -5, 6, -7, 2, -11,
    -- layer=1 filter=164 channel=127
    -12, -2, 8, 0, 2, -6, 3, -4, -3,
    -- layer=1 filter=165 channel=0
    -2, 0, 0, -9, 0, -3, -18, -5, 6,
    -- layer=1 filter=165 channel=1
    4, 2, 6, 5, 3, 5, 7, -6, -7,
    -- layer=1 filter=165 channel=2
    -22, 15, -19, -29, -8, -6, -12, 13, -3,
    -- layer=1 filter=165 channel=3
    11, 0, 11, 5, -7, -6, 0, 6, 1,
    -- layer=1 filter=165 channel=4
    -6, -6, -5, 1, 8, -1, -1, -1, -2,
    -- layer=1 filter=165 channel=5
    21, 13, 39, -21, 19, 7, 43, 6, 14,
    -- layer=1 filter=165 channel=6
    -45, -53, -34, -58, -58, -70, -60, -97, -50,
    -- layer=1 filter=165 channel=7
    -11, -8, -23, 33, 12, -18, 39, 30, 0,
    -- layer=1 filter=165 channel=8
    17, 3, 2, -3, 1, -14, 15, 7, 16,
    -- layer=1 filter=165 channel=9
    -22, -53, -45, -2, -18, 6, -27, -71, -31,
    -- layer=1 filter=165 channel=10
    -4, -13, -4, 25, 17, -24, 40, 46, 15,
    -- layer=1 filter=165 channel=11
    -6, -20, -12, 1, 1, 18, 5, 6, 26,
    -- layer=1 filter=165 channel=12
    -74, -55, -40, 26, -1, 0, -57, -52, -70,
    -- layer=1 filter=165 channel=13
    6, 23, -18, 3, -27, -13, -11, -33, -24,
    -- layer=1 filter=165 channel=14
    -50, -15, -34, 30, 24, -27, -31, 31, -13,
    -- layer=1 filter=165 channel=15
    -32, -33, -14, -25, -27, -52, -10, -38, -8,
    -- layer=1 filter=165 channel=16
    -11, -23, -2, -22, -11, -22, 23, -12, -4,
    -- layer=1 filter=165 channel=17
    12, 2, -7, -8, -16, -15, -7, -16, -5,
    -- layer=1 filter=165 channel=18
    11, -11, -2, 13, 13, -19, -13, -7, -15,
    -- layer=1 filter=165 channel=19
    28, 10, 38, 15, 45, -10, 11, -28, 31,
    -- layer=1 filter=165 channel=20
    0, 10, -12, -14, -25, -34, -27, -36, -43,
    -- layer=1 filter=165 channel=21
    -1, -5, -4, -11, 0, -22, -10, -6, -45,
    -- layer=1 filter=165 channel=22
    -1, 4, 7, -9, -1, -15, -35, -37, -28,
    -- layer=1 filter=165 channel=23
    -23, 6, -18, 6, 10, -71, 55, 2, 15,
    -- layer=1 filter=165 channel=24
    -3, 19, 19, -2, 18, 40, 12, -3, 26,
    -- layer=1 filter=165 channel=25
    -5, -24, -39, -14, -20, -35, 22, 14, -3,
    -- layer=1 filter=165 channel=26
    12, -4, 1, -19, 15, -12, 0, -33, 12,
    -- layer=1 filter=165 channel=27
    -79, -66, -60, -34, -60, -23, 3, -13, -6,
    -- layer=1 filter=165 channel=28
    -30, -12, -15, 29, 18, -27, 21, 46, 1,
    -- layer=1 filter=165 channel=29
    -49, -37, -35, -25, -20, -5, -10, -7, -11,
    -- layer=1 filter=165 channel=30
    52, 22, 25, 44, 32, -1, 15, 7, -3,
    -- layer=1 filter=165 channel=31
    -34, -30, -10, 31, -4, -17, -53, -42, -53,
    -- layer=1 filter=165 channel=32
    -8, 15, 0, 10, 2, -20, 9, 12, 12,
    -- layer=1 filter=165 channel=33
    -4, 6, -2, -10, -1, 4, 9, -1, 13,
    -- layer=1 filter=165 channel=34
    -23, -3, -15, -13, -5, -11, 1, -14, -10,
    -- layer=1 filter=165 channel=35
    -13, -1, -3, -10, -16, -4, -6, -1, -3,
    -- layer=1 filter=165 channel=36
    3, -10, 14, 13, 19, 29, 6, 25, 34,
    -- layer=1 filter=165 channel=37
    21, 17, 24, -4, 15, -11, 31, 2, 17,
    -- layer=1 filter=165 channel=38
    14, 0, 6, -9, -22, -28, -8, -39, -54,
    -- layer=1 filter=165 channel=39
    -16, -30, -6, -9, 4, -18, 0, -3, 7,
    -- layer=1 filter=165 channel=40
    -19, -44, -45, 1, -43, -90, -64, -32, -57,
    -- layer=1 filter=165 channel=41
    -2, 43, -19, -2, 14, -6, 3, -10, -4,
    -- layer=1 filter=165 channel=42
    -34, -29, 0, -53, -29, -25, -32, -22, -32,
    -- layer=1 filter=165 channel=43
    -14, -16, -5, -38, 3, -38, 12, -18, -8,
    -- layer=1 filter=165 channel=44
    -1, -6, 9, 19, 8, 0, 14, 20, 12,
    -- layer=1 filter=165 channel=45
    -11, -29, 10, -9, 5, -26, -7, -40, -11,
    -- layer=1 filter=165 channel=46
    4, -28, 51, -58, -22, -3, -34, -53, -34,
    -- layer=1 filter=165 channel=47
    -52, 58, -41, 9, 17, -34, 23, 19, -5,
    -- layer=1 filter=165 channel=48
    -2, 6, -6, 4, 7, -11, -19, -18, -29,
    -- layer=1 filter=165 channel=49
    -41, -5, -27, -56, -30, -33, -40, -49, -40,
    -- layer=1 filter=165 channel=50
    -5, -5, -4, -7, -19, 0, -9, -17, 4,
    -- layer=1 filter=165 channel=51
    -14, 11, -25, 0, 2, -47, -21, -22, -43,
    -- layer=1 filter=165 channel=52
    11, 8, 15, 8, -10, 6, 27, 13, 7,
    -- layer=1 filter=165 channel=53
    7, 11, 2, -2, -5, -17, 0, -10, -6,
    -- layer=1 filter=165 channel=54
    -7, -12, -16, -13, -10, -34, 21, 5, 30,
    -- layer=1 filter=165 channel=55
    -7, -6, 4, 8, 20, 22, 32, 27, 54,
    -- layer=1 filter=165 channel=56
    -1, 6, -8, 5, 9, 6, 10, 6, 4,
    -- layer=1 filter=165 channel=57
    -18, -32, -46, 6, -16, -71, 5, -2, -14,
    -- layer=1 filter=165 channel=58
    -11, -8, -44, 36, -27, -71, 43, 18, 18,
    -- layer=1 filter=165 channel=59
    -15, -5, -8, -1, -2, -12, -14, -4, -12,
    -- layer=1 filter=165 channel=60
    -12, -8, -11, -12, -22, -2, 1, -6, -4,
    -- layer=1 filter=165 channel=61
    -8, -7, 1, 4, 2, -4, 1, -4, 9,
    -- layer=1 filter=165 channel=62
    7, -6, 3, -28, 4, -26, 24, -12, 4,
    -- layer=1 filter=165 channel=63
    7, -4, 6, -3, 6, 16, -2, 24, 33,
    -- layer=1 filter=165 channel=64
    9, 11, 23, 4, 14, -3, -5, 0, 1,
    -- layer=1 filter=165 channel=65
    7, 14, 10, 7, -6, -15, -24, 0, -36,
    -- layer=1 filter=165 channel=66
    4, -8, 0, 8, 0, 11, 10, 13, 23,
    -- layer=1 filter=165 channel=67
    -22, -20, -22, -1, -23, 5, -52, -48, -37,
    -- layer=1 filter=165 channel=68
    21, -7, 8, 22, 5, 6, 49, 6, 29,
    -- layer=1 filter=165 channel=69
    -6, 1, 9, 0, 18, -19, 19, -5, 14,
    -- layer=1 filter=165 channel=70
    -36, -13, -19, -25, 2, -20, -54, -73, -61,
    -- layer=1 filter=165 channel=71
    -8, -10, 9, -1, 9, 8, 21, 29, 3,
    -- layer=1 filter=165 channel=72
    9, -4, 27, 21, 7, -21, 6, -50, -7,
    -- layer=1 filter=165 channel=73
    3, 0, 4, 0, 9, 9, 2, 11, 11,
    -- layer=1 filter=165 channel=74
    8, -19, 15, -4, -20, -2, -15, -48, -41,
    -- layer=1 filter=165 channel=75
    -17, -33, -3, 25, -33, -61, -20, -1, -40,
    -- layer=1 filter=165 channel=76
    8, -7, -1, -12, -4, -11, 0, -5, -9,
    -- layer=1 filter=165 channel=77
    -22, 0, -2, -10, 11, 2, -13, 5, -22,
    -- layer=1 filter=165 channel=78
    -5, 5, -7, 8, 0, -2, -24, 18, 3,
    -- layer=1 filter=165 channel=79
    -8, -10, -1, -2, -4, -29, 1, -24, -9,
    -- layer=1 filter=165 channel=80
    2, 1, 1, 2, 0, 0, 1, 8, -4,
    -- layer=1 filter=165 channel=81
    -26, -4, -6, -2, 22, 13, 14, 3, 22,
    -- layer=1 filter=165 channel=82
    -8, 11, 18, -4, 18, -7, -13, -18, -24,
    -- layer=1 filter=165 channel=83
    -11, -13, -13, 3, 10, -37, 2, -9, 16,
    -- layer=1 filter=165 channel=84
    34, 11, 6, -2, -22, -3, 0, -20, 9,
    -- layer=1 filter=165 channel=85
    -28, 21, -2, 1, 17, -71, 2, -17, 25,
    -- layer=1 filter=165 channel=86
    0, 2, -5, -4, -5, 8, -3, 19, 12,
    -- layer=1 filter=165 channel=87
    7, 6, 47, -2, -8, -9, -23, -66, -10,
    -- layer=1 filter=165 channel=88
    -10, -8, -9, -24, 1, 10, -46, -24, -24,
    -- layer=1 filter=165 channel=89
    2, -12, 5, -10, -10, -15, -3, -2, -32,
    -- layer=1 filter=165 channel=90
    -4, -14, 1, 8, 6, 0, 34, -16, 9,
    -- layer=1 filter=165 channel=91
    2, 1, 2, -2, -24, -46, -10, -41, -45,
    -- layer=1 filter=165 channel=92
    -27, 0, -34, -15, -37, -36, 6, -5, -38,
    -- layer=1 filter=165 channel=93
    13, 21, 6, 3, 22, 2, 13, 11, 1,
    -- layer=1 filter=165 channel=94
    4, -10, -5, 0, 3, 1, -16, -8, -8,
    -- layer=1 filter=165 channel=95
    32, 7, 20, 12, 1, 3, -1, 14, 1,
    -- layer=1 filter=165 channel=96
    -3, -2, 12, -3, 4, 1, 10, 20, 10,
    -- layer=1 filter=165 channel=97
    0, 16, 2, 13, 21, 11, -1, 3, 4,
    -- layer=1 filter=165 channel=98
    -14, 3, -4, -36, 5, -36, -2, -33, -7,
    -- layer=1 filter=165 channel=99
    -5, 3, -17, 49, 39, -3, 31, 70, 15,
    -- layer=1 filter=165 channel=100
    -15, -14, -4, 2, 6, 19, 10, 17, 13,
    -- layer=1 filter=165 channel=101
    4, 14, 2, 0, -23, -19, -10, -24, -52,
    -- layer=1 filter=165 channel=102
    8, 1, -12, 0, -15, -8, -13, -10, -16,
    -- layer=1 filter=165 channel=103
    -24, -24, -6, -8, -7, -11, -17, -14, 4,
    -- layer=1 filter=165 channel=104
    -16, 33, 4, -8, 30, -25, 2, -8, 17,
    -- layer=1 filter=165 channel=105
    9, 3, 6, 12, 0, 16, 6, 26, 21,
    -- layer=1 filter=165 channel=106
    2, -1, -3, -17, -30, -3, -21, -16, -39,
    -- layer=1 filter=165 channel=107
    1, -5, -8, 0, -18, -18, 14, 0, 9,
    -- layer=1 filter=165 channel=108
    -8, 16, -5, 18, 20, 21, 16, -8, 15,
    -- layer=1 filter=165 channel=109
    -5, 0, 9, -5, 10, 9, 7, -6, -1,
    -- layer=1 filter=165 channel=110
    0, 0, 1, -10, 6, -10, -11, 3, 1,
    -- layer=1 filter=165 channel=111
    58, 3, 15, 25, 4, -14, 0, 6, 0,
    -- layer=1 filter=165 channel=112
    -4, -13, -3, 0, -21, 0, -33, -46, 21,
    -- layer=1 filter=165 channel=113
    -44, -30, -30, -30, -71, -62, -44, -58, -7,
    -- layer=1 filter=165 channel=114
    -19, -23, -14, -41, 0, -26, 31, 12, 10,
    -- layer=1 filter=165 channel=115
    -2, -20, -25, -5, -4, -25, -10, -6, 0,
    -- layer=1 filter=165 channel=116
    1, -2, 4, 2, 9, -11, -11, 3, 6,
    -- layer=1 filter=165 channel=117
    19, -36, -38, 13, -43, -20, -58, -41, -12,
    -- layer=1 filter=165 channel=118
    29, 9, 7, -3, -2, 0, -8, -29, -27,
    -- layer=1 filter=165 channel=119
    -2, 17, 7, -6, 26, 19, 20, 1, 42,
    -- layer=1 filter=165 channel=120
    -9, 9, -20, 5, 0, -35, -8, -11, -32,
    -- layer=1 filter=165 channel=121
    7, -24, -26, 23, -15, 9, 8, 27, 10,
    -- layer=1 filter=165 channel=122
    0, 4, 4, 0, 9, -5, 0, -6, -5,
    -- layer=1 filter=165 channel=123
    -15, -34, -35, 8, -15, 11, 34, 13, 28,
    -- layer=1 filter=165 channel=124
    -9, -18, -15, -6, -12, -16, -10, -21, -10,
    -- layer=1 filter=165 channel=125
    -16, -18, -16, -48, -21, 20, -76, -81, -60,
    -- layer=1 filter=165 channel=126
    6, 20, 13, 0, 22, -38, 0, -6, 12,
    -- layer=1 filter=165 channel=127
    31, 3, 26, 13, 16, -8, 1, -13, -13,
    -- layer=1 filter=166 channel=0
    6, 10, 0, 15, 0, 2, 7, 9, -3,
    -- layer=1 filter=166 channel=1
    18, 32, 25, -18, -9, -20, -8, -28, -28,
    -- layer=1 filter=166 channel=2
    -9, -29, -69, 8, -24, -22, 2, -35, -4,
    -- layer=1 filter=166 channel=3
    -5, 0, 11, -11, 7, 14, -2, 4, 7,
    -- layer=1 filter=166 channel=4
    -8, 0, -2, -3, 4, -5, 3, 6, 2,
    -- layer=1 filter=166 channel=5
    -1, 12, 17, -72, -80, -55, -38, -87, -93,
    -- layer=1 filter=166 channel=6
    -12, 17, 25, 3, 13, 21, 4, 7, 6,
    -- layer=1 filter=166 channel=7
    24, -4, -64, 37, -28, -119, 33, -33, -78,
    -- layer=1 filter=166 channel=8
    13, 38, 40, -75, -79, -82, -56, -120, -102,
    -- layer=1 filter=166 channel=9
    -44, -38, -22, -8, 1, 8, -12, -31, -4,
    -- layer=1 filter=166 channel=10
    34, -22, -98, 37, -44, -94, 35, -29, -84,
    -- layer=1 filter=166 channel=11
    0, 2, 3, -28, -3, 8, -23, -2, -4,
    -- layer=1 filter=166 channel=12
    6, -48, 18, 20, 6, 21, 3, -3, 30,
    -- layer=1 filter=166 channel=13
    2, 14, 35, 0, 3, 14, -22, 9, 5,
    -- layer=1 filter=166 channel=14
    -21, -39, -20, 50, -45, -85, 2, 3, -80,
    -- layer=1 filter=166 channel=15
    -19, 14, 4, -36, -39, 12, -16, -15, -17,
    -- layer=1 filter=166 channel=16
    10, 9, 10, -50, -91, -95, -39, -82, -80,
    -- layer=1 filter=166 channel=17
    1, 8, 19, -4, 12, 24, -2, 14, 21,
    -- layer=1 filter=166 channel=18
    -5, -6, 4, -24, -39, -27, 0, -10, -18,
    -- layer=1 filter=166 channel=19
    -16, -79, -49, -58, -113, -94, -81, -144, -124,
    -- layer=1 filter=166 channel=20
    8, 27, 13, 5, 23, 9, 15, 22, 22,
    -- layer=1 filter=166 channel=21
    3, -1, 7, 1, 7, 1, 21, 7, 0,
    -- layer=1 filter=166 channel=22
    -2, 21, 30, 3, 5, 1, -7, 4, 12,
    -- layer=1 filter=166 channel=23
    -26, -37, -35, -25, -75, -27, -15, -68, -40,
    -- layer=1 filter=166 channel=24
    -17, -3, 24, -20, -16, 5, -27, -19, -1,
    -- layer=1 filter=166 channel=25
    32, -3, -56, 27, -43, -110, 27, -65, -86,
    -- layer=1 filter=166 channel=26
    -32, 3, 35, -28, -25, 37, -46, -21, 13,
    -- layer=1 filter=166 channel=27
    -9, 6, 0, -5, 11, 0, 1, 18, 3,
    -- layer=1 filter=166 channel=28
    22, 7, -23, 36, -6, -58, 27, -18, -30,
    -- layer=1 filter=166 channel=29
    -8, 0, -11, -1, -10, -4, -4, 1, 0,
    -- layer=1 filter=166 channel=30
    -40, -77, -84, -54, -71, -55, -36, -83, -99,
    -- layer=1 filter=166 channel=31
    1, -12, -4, 12, 6, 28, 25, 29, 9,
    -- layer=1 filter=166 channel=32
    -100, -43, 3, -61, -64, 0, -70, -55, 0,
    -- layer=1 filter=166 channel=33
    12, -4, -3, 10, -7, -2, 10, 6, -4,
    -- layer=1 filter=166 channel=34
    23, -14, 0, 2, -5, 9, -3, 6, 0,
    -- layer=1 filter=166 channel=35
    -5, 2, 1, -3, -3, 2, -11, -7, -2,
    -- layer=1 filter=166 channel=36
    2, 9, 17, 2, 0, 15, -13, -1, -7,
    -- layer=1 filter=166 channel=37
    10, 13, 2, -68, -123, -87, -51, -103, -94,
    -- layer=1 filter=166 channel=38
    4, 3, 26, 14, 20, 13, 2, 17, 17,
    -- layer=1 filter=166 channel=39
    6, 7, 15, -15, 5, 1, -15, -5, -1,
    -- layer=1 filter=166 channel=40
    -8, 3, 17, 10, 8, 6, 25, 20, 10,
    -- layer=1 filter=166 channel=41
    -56, -63, 7, 19, -79, -44, -26, -47, -32,
    -- layer=1 filter=166 channel=42
    -28, -54, -39, 33, -47, -12, 38, -44, -3,
    -- layer=1 filter=166 channel=43
    -4, 9, 6, -16, -50, -93, -6, -68, -74,
    -- layer=1 filter=166 channel=44
    -70, -9, 29, -61, -46, 20, -59, -37, -3,
    -- layer=1 filter=166 channel=45
    1, 20, 35, -26, -9, 7, -11, 0, 6,
    -- layer=1 filter=166 channel=46
    -48, -44, -6, -63, -90, -47, -71, -103, -65,
    -- layer=1 filter=166 channel=47
    -27, -50, -32, -27, -71, -4, 5, -51, -29,
    -- layer=1 filter=166 channel=48
    16, 11, 1, 10, 11, 2, 12, 5, 6,
    -- layer=1 filter=166 channel=49
    4, 5, -1, -8, 0, -6, 9, -5, -6,
    -- layer=1 filter=166 channel=50
    4, 5, 19, 6, 14, 11, 23, 11, 19,
    -- layer=1 filter=166 channel=51
    23, 8, -8, 26, 18, -12, 12, 9, -8,
    -- layer=1 filter=166 channel=52
    8, -13, -9, 0, -9, -1, -4, -16, -15,
    -- layer=1 filter=166 channel=53
    19, 12, 2, 10, 8, 21, 2, 5, 0,
    -- layer=1 filter=166 channel=54
    37, -22, -71, -2, -65, -151, 3, -51, -120,
    -- layer=1 filter=166 channel=55
    -19, -23, 5, -41, -24, -12, -33, -13, -9,
    -- layer=1 filter=166 channel=56
    -10, -4, -11, 4, 5, 5, 2, -7, 6,
    -- layer=1 filter=166 channel=57
    26, -1, -50, 30, -3, -40, 23, -13, -29,
    -- layer=1 filter=166 channel=58
    10, -54, -95, -27, -135, -134, -14, -69, -102,
    -- layer=1 filter=166 channel=59
    9, 9, -5, -10, -11, -7, -7, -1, 6,
    -- layer=1 filter=166 channel=60
    17, -6, 1, 17, 11, 9, 2, 13, 16,
    -- layer=1 filter=166 channel=61
    -12, -5, 0, 0, -5, -5, -2, -11, 0,
    -- layer=1 filter=166 channel=62
    2, 17, 18, -71, -125, -75, -77, -138, -109,
    -- layer=1 filter=166 channel=63
    -13, 1, 6, -14, -12, -13, -7, 2, -10,
    -- layer=1 filter=166 channel=64
    -3, 12, 11, -5, 1, -5, 1, -1, -12,
    -- layer=1 filter=166 channel=65
    5, 17, 3, 10, 16, 0, 3, 2, -5,
    -- layer=1 filter=166 channel=66
    -4, 4, 0, -6, 9, 0, 7, -4, 3,
    -- layer=1 filter=166 channel=67
    -11, 2, -6, -22, -15, -11, -17, -13, -8,
    -- layer=1 filter=166 channel=68
    -92, -18, 45, -65, -53, 19, -81, -25, -4,
    -- layer=1 filter=166 channel=69
    -5, 18, 30, -84, -69, -6, -64, -61, -33,
    -- layer=1 filter=166 channel=70
    27, 18, 16, 17, 13, 18, 18, 27, 9,
    -- layer=1 filter=166 channel=71
    3, -3, 0, 13, -3, 0, 18, 6, 4,
    -- layer=1 filter=166 channel=72
    -39, -101, -45, -49, -70, -66, -43, -115, -69,
    -- layer=1 filter=166 channel=73
    5, -11, 3, -10, -8, -10, -3, 6, 0,
    -- layer=1 filter=166 channel=74
    -61, -21, 41, -13, -4, 8, -30, 11, -36,
    -- layer=1 filter=166 channel=75
    -39, -29, -25, 15, -79, -58, -51, -89, -80,
    -- layer=1 filter=166 channel=76
    -11, 17, 14, -6, 4, 14, -6, 18, -13,
    -- layer=1 filter=166 channel=77
    7, 9, 8, 8, 8, -3, -5, 9, 4,
    -- layer=1 filter=166 channel=78
    -3, 2, -10, -12, -1, 7, -3, 2, -14,
    -- layer=1 filter=166 channel=79
    5, 25, 22, -62, -85, -58, -36, -77, -75,
    -- layer=1 filter=166 channel=80
    -7, 1, -6, 10, -4, 6, -6, 0, 6,
    -- layer=1 filter=166 channel=81
    1, -1, 9, -3, -10, -6, 12, -7, 4,
    -- layer=1 filter=166 channel=82
    15, 10, 11, 11, 18, 18, 12, 7, 12,
    -- layer=1 filter=166 channel=83
    0, 33, 23, -15, -39, 11, -26, -38, -11,
    -- layer=1 filter=166 channel=84
    -93, -88, -7, -82, -66, -37, -44, -41, -50,
    -- layer=1 filter=166 channel=85
    7, -7, -20, -18, -87, -31, 10, -12, -24,
    -- layer=1 filter=166 channel=86
    -13, 12, 0, -7, 4, -8, 2, 2, 1,
    -- layer=1 filter=166 channel=87
    -38, -26, -14, -21, -32, -2, 18, -69, -13,
    -- layer=1 filter=166 channel=88
    7, 4, -8, 1, 8, 5, 4, 12, 4,
    -- layer=1 filter=166 channel=89
    12, 10, 23, 6, 5, 25, 8, 15, 2,
    -- layer=1 filter=166 channel=90
    -74, 13, 59, -100, -75, 11, -111, -57, -14,
    -- layer=1 filter=166 channel=91
    6, 16, 2, 12, 8, 20, 23, 19, 24,
    -- layer=1 filter=166 channel=92
    -30, -48, -18, -49, -36, -1, -17, 0, -48,
    -- layer=1 filter=166 channel=93
    16, 22, 16, 3, 17, -2, 2, 13, 6,
    -- layer=1 filter=166 channel=94
    8, 22, 12, 12, 10, -4, 11, 19, 13,
    -- layer=1 filter=166 channel=95
    -81, -76, -8, -88, -94, -51, -75, -75, -87,
    -- layer=1 filter=166 channel=96
    -8, -18, -17, -14, 0, -15, -7, -10, -7,
    -- layer=1 filter=166 channel=97
    12, 15, 8, 6, 6, 4, 15, -2, 13,
    -- layer=1 filter=166 channel=98
    24, 53, 27, -19, -51, -41, -20, -59, -61,
    -- layer=1 filter=166 channel=99
    -4, -27, -28, 32, -12, -45, 32, 0, -26,
    -- layer=1 filter=166 channel=100
    0, -2, 15, -12, -8, -16, -38, -20, -3,
    -- layer=1 filter=166 channel=101
    5, 20, 25, 9, 12, 15, 15, 15, 21,
    -- layer=1 filter=166 channel=102
    10, 9, 14, 20, 28, 13, 11, 16, 12,
    -- layer=1 filter=166 channel=103
    14, 19, 20, -7, 6, 10, 0, 10, 8,
    -- layer=1 filter=166 channel=104
    20, -9, -21, -1, -19, -3, 1, -4, -8,
    -- layer=1 filter=166 channel=105
    15, 23, 0, 25, 16, 6, 10, 16, -1,
    -- layer=1 filter=166 channel=106
    3, 6, 29, -2, 4, 20, -8, 13, 13,
    -- layer=1 filter=166 channel=107
    6, 7, 12, 8, 19, 16, 3, 17, 8,
    -- layer=1 filter=166 channel=108
    -92, 0, 30, -75, -87, -9, -90, -70, -25,
    -- layer=1 filter=166 channel=109
    -2, -11, -4, 4, 4, 8, -5, -3, 6,
    -- layer=1 filter=166 channel=110
    1, -5, 1, 5, 0, 4, -8, 4, 2,
    -- layer=1 filter=166 channel=111
    -35, -31, -20, -30, -44, -41, 0, -5, -62,
    -- layer=1 filter=166 channel=112
    -49, -54, -15, -15, -57, -52, -10, -14, -63,
    -- layer=1 filter=166 channel=113
    8, 5, -13, 18, -12, -13, 9, 14, 6,
    -- layer=1 filter=166 channel=114
    -24, -1, 12, -30, 8, 2, -21, -18, -23,
    -- layer=1 filter=166 channel=115
    14, 7, -25, 12, 8, -18, 13, 5, -8,
    -- layer=1 filter=166 channel=116
    7, 0, 4, 6, -9, 10, 3, -3, -3,
    -- layer=1 filter=166 channel=117
    -76, -81, -47, -75, -92, -95, -31, -45, -82,
    -- layer=1 filter=166 channel=118
    -62, -27, 0, -49, -9, -6, -18, -9, -13,
    -- layer=1 filter=166 channel=119
    -73, -25, 12, -68, -67, -1, -88, -72, -7,
    -- layer=1 filter=166 channel=120
    28, 18, -5, 10, -1, -13, 9, 7, -1,
    -- layer=1 filter=166 channel=121
    -5, 4, -16, -6, -24, -22, -34, -61, -29,
    -- layer=1 filter=166 channel=122
    0, -4, 7, -1, -7, 7, 5, 10, 2,
    -- layer=1 filter=166 channel=123
    1, -8, -11, -17, -14, -15, -29, -36, -23,
    -- layer=1 filter=166 channel=124
    8, -11, 2, -3, 6, 8, -2, 0, 0,
    -- layer=1 filter=166 channel=125
    7, 1, 4, 3, -13, 5, 5, 6, 6,
    -- layer=1 filter=166 channel=126
    11, 42, 11, -61, -58, -44, -67, -83, -64,
    -- layer=1 filter=166 channel=127
    -87, -86, -24, -72, -45, -55, -43, -58, -74,
    -- layer=1 filter=167 channel=0
    5, 11, 2, -1, 4, -13, -2, -19, -17,
    -- layer=1 filter=167 channel=1
    12, 8, 3, 0, 15, 8, -29, -22, 17,
    -- layer=1 filter=167 channel=2
    -23, 1, -17, -43, -25, -36, -17, -20, -22,
    -- layer=1 filter=167 channel=3
    2, -4, 14, 3, -7, -15, 18, 8, 0,
    -- layer=1 filter=167 channel=4
    8, -8, -8, 2, -3, 4, 10, -1, -3,
    -- layer=1 filter=167 channel=5
    8, -5, -25, -24, -16, -14, -60, -9, 4,
    -- layer=1 filter=167 channel=6
    -35, -13, -14, 6, 16, 4, 26, 29, 16,
    -- layer=1 filter=167 channel=7
    -53, -69, -34, -38, -87, -23, -41, -79, -39,
    -- layer=1 filter=167 channel=8
    25, 8, 16, -5, 18, 0, -77, -44, -31,
    -- layer=1 filter=167 channel=9
    -22, 27, 17, -10, -32, -30, 0, -33, -57,
    -- layer=1 filter=167 channel=10
    -37, -92, -53, -28, -87, -18, -21, -38, -23,
    -- layer=1 filter=167 channel=11
    33, 23, 19, 7, 2, 5, -12, 5, -9,
    -- layer=1 filter=167 channel=12
    -19, 3, -13, -9, 11, 23, -88, -76, -57,
    -- layer=1 filter=167 channel=13
    9, 9, 7, 7, 22, -2, 1, 7, -11,
    -- layer=1 filter=167 channel=14
    -37, -45, -36, -34, -53, -19, -38, -68, -36,
    -- layer=1 filter=167 channel=15
    -18, -10, -27, -25, -24, -5, -21, 1, -24,
    -- layer=1 filter=167 channel=16
    32, 13, 12, 0, -8, -2, -69, -38, -48,
    -- layer=1 filter=167 channel=17
    33, 20, 19, 7, 12, 0, -8, -16, -29,
    -- layer=1 filter=167 channel=18
    40, 21, 9, 30, 26, 12, 23, 0, -1,
    -- layer=1 filter=167 channel=19
    9, 0, 33, 0, -5, -38, 41, 23, 14,
    -- layer=1 filter=167 channel=20
    12, 15, 16, 0, 19, 17, 5, 7, -1,
    -- layer=1 filter=167 channel=21
    -5, 6, -14, -17, 2, 5, -17, -4, 6,
    -- layer=1 filter=167 channel=22
    12, -3, 0, 4, 16, 24, -5, 3, -3,
    -- layer=1 filter=167 channel=23
    0, 0, -15, -26, -47, -33, -22, -49, -54,
    -- layer=1 filter=167 channel=24
    -9, -19, -3, -26, -21, -26, -16, -18, -24,
    -- layer=1 filter=167 channel=25
    5, -33, -4, -5, -19, -15, -43, -73, -63,
    -- layer=1 filter=167 channel=26
    32, 33, 20, 33, 21, -18, 0, -6, -48,
    -- layer=1 filter=167 channel=27
    22, 34, 36, 5, 18, 24, 1, 11, 0,
    -- layer=1 filter=167 channel=28
    -12, -39, -16, -12, -52, -7, -24, -64, -31,
    -- layer=1 filter=167 channel=29
    -11, 5, 8, -6, 2, -12, 6, -14, -23,
    -- layer=1 filter=167 channel=30
    27, 10, 3, 21, 38, 22, 50, 27, -1,
    -- layer=1 filter=167 channel=31
    -18, -23, -16, 10, 16, 9, -6, 7, 0,
    -- layer=1 filter=167 channel=32
    19, 1, -21, 30, 2, -44, 16, -2, -38,
    -- layer=1 filter=167 channel=33
    2, 15, -8, 0, 9, 14, 6, -14, -15,
    -- layer=1 filter=167 channel=34
    -15, -7, -8, -19, 7, 6, 13, 18, -5,
    -- layer=1 filter=167 channel=35
    -1, 1, -3, -3, -8, -2, -15, -1, -3,
    -- layer=1 filter=167 channel=36
    27, 7, 12, 2, -6, 1, -18, -1, -15,
    -- layer=1 filter=167 channel=37
    23, -4, 1, -8, -7, -13, -60, -11, -19,
    -- layer=1 filter=167 channel=38
    4, 1, 9, 9, 20, 29, 16, 13, 17,
    -- layer=1 filter=167 channel=39
    20, 3, 8, 0, -6, -17, -14, -4, 0,
    -- layer=1 filter=167 channel=40
    7, -9, -3, 19, 14, 32, 34, 14, 24,
    -- layer=1 filter=167 channel=41
    48, 29, -2, 39, -38, -56, 15, -24, -80,
    -- layer=1 filter=167 channel=42
    -21, -20, -11, -29, -17, -6, -21, -34, -23,
    -- layer=1 filter=167 channel=43
    27, -5, -12, -3, 2, -14, -75, -53, -37,
    -- layer=1 filter=167 channel=44
    21, 10, -6, 30, 6, -49, 1, -6, -47,
    -- layer=1 filter=167 channel=45
    -11, -1, -3, -16, -9, -6, -18, -2, -16,
    -- layer=1 filter=167 channel=46
    -31, -47, 0, -35, -29, -47, 9, 23, 38,
    -- layer=1 filter=167 channel=47
    -56, -25, -35, -17, -27, -45, 0, -12, -15,
    -- layer=1 filter=167 channel=48
    -9, 0, 1, -9, -8, 18, 9, 5, 11,
    -- layer=1 filter=167 channel=49
    -34, -25, -19, -1, 0, -15, 12, 1, -8,
    -- layer=1 filter=167 channel=50
    -3, 15, 17, 15, 10, 7, -8, -23, -32,
    -- layer=1 filter=167 channel=51
    -13, -29, -2, 5, -5, 27, 7, -4, 27,
    -- layer=1 filter=167 channel=52
    8, -3, -12, -16, -14, -3, 0, -12, 4,
    -- layer=1 filter=167 channel=53
    8, 9, 9, 2, 17, 0, 12, 14, -3,
    -- layer=1 filter=167 channel=54
    2, -25, -20, 11, -8, -8, -30, -59, -44,
    -- layer=1 filter=167 channel=55
    17, -4, 8, 0, -9, -9, -23, -15, -13,
    -- layer=1 filter=167 channel=56
    -4, 7, -1, 3, -6, 9, 6, 0, -7,
    -- layer=1 filter=167 channel=57
    -43, -72, -40, -20, -48, 9, 1, -14, -7,
    -- layer=1 filter=167 channel=58
    -38, -63, -43, -58, -101, -62, -3, -66, -69,
    -- layer=1 filter=167 channel=59
    -14, 5, -13, -9, -14, -7, -4, 0, -1,
    -- layer=1 filter=167 channel=60
    13, 1, -2, -2, 16, 3, 16, 3, 14,
    -- layer=1 filter=167 channel=61
    2, -4, 8, 12, -3, -3, 9, 7, 4,
    -- layer=1 filter=167 channel=62
    32, 7, 18, 8, 0, 12, -84, -34, -42,
    -- layer=1 filter=167 channel=63
    17, 10, 5, -3, -6, -1, -9, -7, -25,
    -- layer=1 filter=167 channel=64
    -7, 1, 1, -6, 10, -3, 0, 5, -2,
    -- layer=1 filter=167 channel=65
    1, -2, 13, -2, 5, 19, 0, -1, 14,
    -- layer=1 filter=167 channel=66
    15, 9, -3, 10, -1, -16, -8, -14, -18,
    -- layer=1 filter=167 channel=67
    -88, -75, -81, -29, -30, -38, -28, -11, -8,
    -- layer=1 filter=167 channel=68
    17, 2, -4, 38, -2, -38, -9, -13, -44,
    -- layer=1 filter=167 channel=69
    14, -15, -19, -24, -25, -39, -48, -15, -46,
    -- layer=1 filter=167 channel=70
    -36, -47, -57, 0, 6, -4, 0, 9, 13,
    -- layer=1 filter=167 channel=71
    0, -5, -17, -10, -5, 2, -19, -5, -1,
    -- layer=1 filter=167 channel=72
    -8, 1, 24, 5, 6, -1, 25, 12, 21,
    -- layer=1 filter=167 channel=73
    -2, 2, 2, -9, -1, 4, -12, -13, -3,
    -- layer=1 filter=167 channel=74
    29, 5, -24, 24, 15, -24, 16, -19, -10,
    -- layer=1 filter=167 channel=75
    -11, -27, -33, -36, -39, -3, -18, -28, -16,
    -- layer=1 filter=167 channel=76
    12, 10, -2, 13, 12, -9, 23, 1, -31,
    -- layer=1 filter=167 channel=77
    2, -4, 5, -6, -8, 8, -8, -4, -1,
    -- layer=1 filter=167 channel=78
    7, 0, -9, 1, -16, -19, -10, -9, -15,
    -- layer=1 filter=167 channel=79
    34, 9, 12, 10, -3, 8, -69, -22, -28,
    -- layer=1 filter=167 channel=80
    -3, -5, 1, 10, 8, 7, 7, 7, 0,
    -- layer=1 filter=167 channel=81
    -8, 9, 19, -22, -3, 0, -23, -20, -25,
    -- layer=1 filter=167 channel=82
    -16, 3, -3, 8, 16, 13, -8, 21, 14,
    -- layer=1 filter=167 channel=83
    13, -19, 14, -17, -27, -14, -11, -17, -22,
    -- layer=1 filter=167 channel=84
    52, 43, 32, 56, 54, 31, 47, 6, -21,
    -- layer=1 filter=167 channel=85
    0, -29, -19, -12, -42, -26, 20, -42, -39,
    -- layer=1 filter=167 channel=86
    14, 23, 10, 13, -13, -10, -25, -12, -23,
    -- layer=1 filter=167 channel=87
    -38, 8, 0, -24, 0, -55, 25, -3, 4,
    -- layer=1 filter=167 channel=88
    -24, -15, -28, -6, 0, -7, 0, -7, 2,
    -- layer=1 filter=167 channel=89
    2, 11, -4, 6, 12, 0, 6, 17, 8,
    -- layer=1 filter=167 channel=90
    8, -22, -8, 0, -38, -47, -8, -34, -70,
    -- layer=1 filter=167 channel=91
    7, -11, 9, 9, 22, 19, 26, 22, 22,
    -- layer=1 filter=167 channel=92
    6, -38, -7, -6, -66, -68, -1, -30, -75,
    -- layer=1 filter=167 channel=93
    8, -6, -1, -7, -3, 4, 1, -14, -1,
    -- layer=1 filter=167 channel=94
    13, 17, 10, 12, -8, 8, -15, -12, -21,
    -- layer=1 filter=167 channel=95
    35, 16, 9, 48, 27, 31, 38, 8, -6,
    -- layer=1 filter=167 channel=96
    8, 5, 6, -1, 1, 10, -1, 7, 0,
    -- layer=1 filter=167 channel=97
    22, 21, 12, 4, -2, 0, -11, -1, -8,
    -- layer=1 filter=167 channel=98
    23, -2, 5, 9, 20, 20, -51, -31, -17,
    -- layer=1 filter=167 channel=99
    -28, -70, -27, 0, -42, -46, 18, -31, -35,
    -- layer=1 filter=167 channel=100
    17, 17, 7, 17, 18, 14, -12, 5, -10,
    -- layer=1 filter=167 channel=101
    10, -1, 1, 20, 26, 27, 12, 26, 13,
    -- layer=1 filter=167 channel=102
    27, 20, 11, 29, 0, 17, 16, -4, 12,
    -- layer=1 filter=167 channel=103
    19, 5, 23, 12, 4, 13, -8, 0, 0,
    -- layer=1 filter=167 channel=104
    -7, 0, -5, 12, -7, -25, 31, -22, -17,
    -- layer=1 filter=167 channel=105
    22, 7, 14, 7, -9, -6, -15, -20, -22,
    -- layer=1 filter=167 channel=106
    -2, 1, -12, 18, 39, 12, 32, 30, 7,
    -- layer=1 filter=167 channel=107
    12, 8, -2, 4, 11, 6, 5, -4, -5,
    -- layer=1 filter=167 channel=108
    2, -14, -18, 11, -26, -69, -2, -25, -99,
    -- layer=1 filter=167 channel=109
    3, 5, -9, 0, 0, -4, -5, -4, -5,
    -- layer=1 filter=167 channel=110
    0, 10, -8, 9, -3, 5, -5, 0, -3,
    -- layer=1 filter=167 channel=111
    38, 28, 7, 27, 26, 36, 41, 26, -22,
    -- layer=1 filter=167 channel=112
    20, 6, -12, 43, 14, 5, 10, 3, -18,
    -- layer=1 filter=167 channel=113
    -40, -47, -21, -5, -22, 0, 13, -4, 2,
    -- layer=1 filter=167 channel=114
    5, 8, 4, 0, -10, -30, -34, -13, -25,
    -- layer=1 filter=167 channel=115
    7, -3, 0, 8, -8, 7, -21, -26, -10,
    -- layer=1 filter=167 channel=116
    6, 8, -3, 4, -2, 5, -11, 4, -7,
    -- layer=1 filter=167 channel=117
    24, -3, 2, 44, 32, 22, 14, -2, -21,
    -- layer=1 filter=167 channel=118
    26, 25, 10, 22, 44, 15, 47, 13, -1,
    -- layer=1 filter=167 channel=119
    11, -22, -6, 10, -11, -50, 2, -26, -76,
    -- layer=1 filter=167 channel=120
    -6, 0, 0, -9, 0, 20, -16, -5, 5,
    -- layer=1 filter=167 channel=121
    -23, -27, -20, -10, 0, 2, -4, 0, 8,
    -- layer=1 filter=167 channel=122
    9, -1, -7, -8, -4, 2, -7, 7, 0,
    -- layer=1 filter=167 channel=123
    11, -8, 4, 2, -7, 19, 12, -9, 8,
    -- layer=1 filter=167 channel=124
    -2, -3, -10, -15, -3, -9, -15, -5, -6,
    -- layer=1 filter=167 channel=125
    -33, -61, -50, -15, -12, -11, 3, 10, 24,
    -- layer=1 filter=167 channel=126
    -4, -22, -5, -4, 13, 25, -63, -17, -7,
    -- layer=1 filter=167 channel=127
    38, 32, 6, 46, 56, 30, 45, 16, 13,
    -- layer=1 filter=168 channel=0
    -21, -10, -12, 2, -8, -24, 2, 0, -3,
    -- layer=1 filter=168 channel=1
    -5, -14, -30, 0, -14, 7, 17, 0, 14,
    -- layer=1 filter=168 channel=2
    -29, -29, 13, -57, -7, -12, -2, 13, -6,
    -- layer=1 filter=168 channel=3
    1, -9, 0, -2, -20, -10, -9, -11, -7,
    -- layer=1 filter=168 channel=4
    -5, 8, 3, -5, 8, 8, -6, -4, -2,
    -- layer=1 filter=168 channel=5
    18, 11, -2, 17, 5, 22, 15, -4, 13,
    -- layer=1 filter=168 channel=6
    37, 54, 35, 33, 8, -13, 20, 9, -5,
    -- layer=1 filter=168 channel=7
    5, 20, 14, -6, -6, 75, -33, -32, 55,
    -- layer=1 filter=168 channel=8
    23, -10, 2, 9, 19, 23, 24, 8, 17,
    -- layer=1 filter=168 channel=9
    -4, 2, -19, -18, 43, -15, -2, 62, -34,
    -- layer=1 filter=168 channel=10
    -12, 7, 39, -9, -20, 62, -62, -55, 38,
    -- layer=1 filter=168 channel=11
    -20, 17, 11, 0, 17, -6, 6, 26, 5,
    -- layer=1 filter=168 channel=12
    -48, -70, -12, -59, -77, -53, 48, 18, 12,
    -- layer=1 filter=168 channel=13
    26, 22, 20, 12, 28, -35, 19, 2, -19,
    -- layer=1 filter=168 channel=14
    -18, -26, 13, -3, -6, 35, -19, -34, 57,
    -- layer=1 filter=168 channel=15
    1, 38, 14, 18, 48, 16, 15, 16, -10,
    -- layer=1 filter=168 channel=16
    31, 9, 0, 7, 4, 34, 30, 16, 14,
    -- layer=1 filter=168 channel=17
    -9, -27, -2, 0, 20, -5, 11, 19, 0,
    -- layer=1 filter=168 channel=18
    -25, 4, 21, -8, -2, -16, 0, -7, -3,
    -- layer=1 filter=168 channel=19
    22, -3, 31, 4, 8, 43, 12, 36, 6,
    -- layer=1 filter=168 channel=20
    13, 5, -4, 11, -11, -9, 22, 2, -20,
    -- layer=1 filter=168 channel=21
    9, -18, -37, -16, -41, -42, 7, -16, 6,
    -- layer=1 filter=168 channel=22
    23, 12, -12, 13, 9, -2, 26, 13, -2,
    -- layer=1 filter=168 channel=23
    9, 45, 28, 13, 29, 87, -27, 31, 50,
    -- layer=1 filter=168 channel=24
    -10, -30, -8, -22, -12, -28, -14, 5, -36,
    -- layer=1 filter=168 channel=25
    1, 2, 12, -4, 4, 68, -19, -35, 42,
    -- layer=1 filter=168 channel=26
    10, 25, 22, 0, 40, -12, 4, 37, -43,
    -- layer=1 filter=168 channel=27
    -15, -16, 23, -35, -12, -20, -4, -22, -21,
    -- layer=1 filter=168 channel=28
    -16, -7, 1, -24, -15, 41, -36, -49, 25,
    -- layer=1 filter=168 channel=29
    4, -2, 9, -4, -3, 11, 21, 13, 28,
    -- layer=1 filter=168 channel=30
    -37, -16, 16, -30, -31, -6, -42, -3, -46,
    -- layer=1 filter=168 channel=31
    -13, 23, 20, 7, 4, 0, 4, 16, -8,
    -- layer=1 filter=168 channel=32
    10, 24, 27, 6, 57, 6, -7, 24, -18,
    -- layer=1 filter=168 channel=33
    12, 15, -4, 0, -2, -5, 8, -8, -17,
    -- layer=1 filter=168 channel=34
    16, 43, 15, 20, 5, -10, 20, 19, -24,
    -- layer=1 filter=168 channel=35
    -1, 10, 16, 2, 8, 14, 15, 0, 4,
    -- layer=1 filter=168 channel=36
    -22, 6, -2, -6, 13, 0, -1, 0, 2,
    -- layer=1 filter=168 channel=37
    21, 16, 14, 0, 6, 16, 11, 4, 7,
    -- layer=1 filter=168 channel=38
    14, 2, 2, -6, -22, -38, 5, -18, -20,
    -- layer=1 filter=168 channel=39
    -17, -20, -4, 4, 8, 6, 14, 18, 1,
    -- layer=1 filter=168 channel=40
    2, 9, 26, -1, -3, -2, -3, -35, -17,
    -- layer=1 filter=168 channel=41
    -7, -20, 54, -34, 40, 9, -13, 75, 18,
    -- layer=1 filter=168 channel=42
    -33, -29, -24, -64, -42, -4, -24, -20, 13,
    -- layer=1 filter=168 channel=43
    0, -14, -18, 0, -25, 17, 17, 1, 29,
    -- layer=1 filter=168 channel=44
    2, 27, 15, -3, 57, -7, 9, -5, -33,
    -- layer=1 filter=168 channel=45
    20, -3, -19, 9, 4, -17, 14, -7, -8,
    -- layer=1 filter=168 channel=46
    15, -1, 16, 15, -12, 22, 29, 13, 2,
    -- layer=1 filter=168 channel=47
    14, 35, 68, 5, 40, 49, -28, 38, 12,
    -- layer=1 filter=168 channel=48
    -2, -35, -17, -5, -46, -36, -12, -35, -19,
    -- layer=1 filter=168 channel=49
    22, 15, 6, 2, 12, -12, 6, 30, -13,
    -- layer=1 filter=168 channel=50
    2, 4, -7, -7, -4, 0, 1, -13, -16,
    -- layer=1 filter=168 channel=51
    5, -17, 0, -10, -44, 13, -14, -58, 3,
    -- layer=1 filter=168 channel=52
    1, 17, -4, 10, 20, 0, 4, 23, 0,
    -- layer=1 filter=168 channel=53
    0, 28, -24, 0, -1, 9, -7, 13, 15,
    -- layer=1 filter=168 channel=54
    12, -12, 20, -12, 0, 53, -8, -29, 32,
    -- layer=1 filter=168 channel=55
    -13, 9, 32, 5, 25, 13, -13, 8, 0,
    -- layer=1 filter=168 channel=56
    5, 8, 10, 1, -3, 16, 9, 12, 13,
    -- layer=1 filter=168 channel=57
    -5, 0, 27, 0, -12, 61, -41, -53, 25,
    -- layer=1 filter=168 channel=58
    37, 51, 81, 8, 40, 112, -45, 24, 58,
    -- layer=1 filter=168 channel=59
    8, 12, 5, -2, 8, 8, 2, 14, -1,
    -- layer=1 filter=168 channel=60
    0, 1, 13, 23, 9, 14, 3, -3, 21,
    -- layer=1 filter=168 channel=61
    0, -3, -10, 12, -5, 1, 12, 5, -6,
    -- layer=1 filter=168 channel=62
    11, -11, -7, -6, -7, 38, 24, 10, 4,
    -- layer=1 filter=168 channel=63
    -2, 1, 0, -10, 8, -15, 7, 1, 5,
    -- layer=1 filter=168 channel=64
    13, 8, -13, -5, -6, -15, 14, 0, 0,
    -- layer=1 filter=168 channel=65
    -6, -30, -39, -25, -47, -33, -9, -33, -7,
    -- layer=1 filter=168 channel=66
    1, -4, -1, -3, -20, -11, -10, -13, 0,
    -- layer=1 filter=168 channel=67
    51, 55, 59, 28, -2, -28, 35, -9, -39,
    -- layer=1 filter=168 channel=68
    24, 36, -8, 26, 61, -19, 17, 14, -21,
    -- layer=1 filter=168 channel=69
    -11, 8, 10, -7, 6, -3, 11, 26, 0,
    -- layer=1 filter=168 channel=70
    33, 49, 27, 40, 21, 7, 40, 21, -16,
    -- layer=1 filter=168 channel=71
    -22, -41, -37, -29, -47, -5, -3, -36, 6,
    -- layer=1 filter=168 channel=72
    11, -1, 44, -13, -24, 26, 17, 37, -18,
    -- layer=1 filter=168 channel=73
    0, 4, 1, 12, 4, 13, -7, -6, 1,
    -- layer=1 filter=168 channel=74
    3, 33, -11, 4, 21, -14, 3, -6, 9,
    -- layer=1 filter=168 channel=75
    -39, -15, -21, -9, -17, -11, 18, -22, 4,
    -- layer=1 filter=168 channel=76
    -16, 2, -1, -10, -5, -46, -3, -20, -38,
    -- layer=1 filter=168 channel=77
    -2, -20, -43, -25, -46, -48, -10, -30, -22,
    -- layer=1 filter=168 channel=78
    -9, -7, 24, -7, 6, 29, -15, -9, 26,
    -- layer=1 filter=168 channel=79
    1, 4, -12, -7, -6, 27, 14, 11, 14,
    -- layer=1 filter=168 channel=80
    -2, -4, -1, 2, 5, 21, -1, 20, 11,
    -- layer=1 filter=168 channel=81
    -14, -38, -39, -4, -34, -17, -12, -13, -21,
    -- layer=1 filter=168 channel=82
    1, -25, -23, -23, -50, -53, -6, -33, -35,
    -- layer=1 filter=168 channel=83
    -1, -5, -12, 12, 16, -10, 17, 20, -7,
    -- layer=1 filter=168 channel=84
    3, 4, -6, -1, 17, -37, -10, 0, -34,
    -- layer=1 filter=168 channel=85
    51, 33, 68, -2, 26, 91, -45, 34, 50,
    -- layer=1 filter=168 channel=86
    -9, 6, 2, 6, 7, 9, -8, -6, 5,
    -- layer=1 filter=168 channel=87
    29, 0, 29, 18, 4, 51, 17, 59, -17,
    -- layer=1 filter=168 channel=88
    4, -13, -12, 5, -25, -27, 0, -14, -24,
    -- layer=1 filter=168 channel=89
    -5, -25, -33, -19, -45, -57, 5, -56, -40,
    -- layer=1 filter=168 channel=90
    14, 29, 24, 9, 72, 6, 21, 37, -12,
    -- layer=1 filter=168 channel=91
    18, 16, 1, 12, -14, -22, 4, -15, -29,
    -- layer=1 filter=168 channel=92
    -5, 37, 35, 7, 67, 2, 15, 16, -15,
    -- layer=1 filter=168 channel=93
    -14, -63, -54, -19, -51, -36, -8, -44, -16,
    -- layer=1 filter=168 channel=94
    -10, -7, -23, -2, -12, -13, -10, -6, -12,
    -- layer=1 filter=168 channel=95
    -12, 8, -13, -25, -4, -48, -19, -7, -19,
    -- layer=1 filter=168 channel=96
    13, 7, -1, 6, -5, -4, 12, -5, -5,
    -- layer=1 filter=168 channel=97
    -22, -42, -50, -19, -30, -22, -2, -21, -17,
    -- layer=1 filter=168 channel=98
    8, -19, -13, -16, -27, 20, 11, 12, 24,
    -- layer=1 filter=168 channel=99
    10, 37, 46, 1, 35, 29, -64, -35, 42,
    -- layer=1 filter=168 channel=100
    -14, 12, 16, -2, 10, -22, -2, 14, -6,
    -- layer=1 filter=168 channel=101
    -1, 4, -14, 1, -31, -49, 1, -26, -19,
    -- layer=1 filter=168 channel=102
    -21, -5, -20, -26, -25, -31, -6, -29, -29,
    -- layer=1 filter=168 channel=103
    -7, 4, 15, -8, -2, -9, -2, 20, -9,
    -- layer=1 filter=168 channel=104
    2, 24, 63, 1, 40, 56, -19, 36, 38,
    -- layer=1 filter=168 channel=105
    -36, -30, -31, -14, -41, -24, -4, -35, -9,
    -- layer=1 filter=168 channel=106
    23, 20, 5, 16, 22, -33, 15, -11, -35,
    -- layer=1 filter=168 channel=107
    0, -10, -3, -2, -8, -2, 0, 4, 16,
    -- layer=1 filter=168 channel=108
    14, 29, 30, -3, 44, -7, 13, 43, -18,
    -- layer=1 filter=168 channel=109
    4, -8, 0, -10, -5, 6, 4, 3, 3,
    -- layer=1 filter=168 channel=110
    -2, -9, -7, -2, -9, 2, -8, 2, 4,
    -- layer=1 filter=168 channel=111
    -41, -20, 1, -20, -5, -20, -40, -21, -40,
    -- layer=1 filter=168 channel=112
    -18, 8, -21, 23, 20, -22, -15, -24, -17,
    -- layer=1 filter=168 channel=113
    23, 24, 11, 12, 11, 26, 17, -3, 24,
    -- layer=1 filter=168 channel=114
    16, 21, 17, 19, 17, 10, 34, 21, 22,
    -- layer=1 filter=168 channel=115
    -23, -13, 1, -9, -26, 27, -33, -41, 22,
    -- layer=1 filter=168 channel=116
    3, -6, -1, -8, 0, 7, 9, -6, -6,
    -- layer=1 filter=168 channel=117
    -19, -14, 15, 40, 10, 31, -27, -48, -3,
    -- layer=1 filter=168 channel=118
    -18, 12, -1, -22, -13, -66, -8, -13, -26,
    -- layer=1 filter=168 channel=119
    14, 16, 37, 4, 65, -4, 13, 37, -25,
    -- layer=1 filter=168 channel=120
    7, -11, -21, -8, -26, 3, -6, -23, -4,
    -- layer=1 filter=168 channel=121
    -25, 10, 18, -23, 12, 2, -2, 16, 24,
    -- layer=1 filter=168 channel=122
    9, -5, -3, -1, -6, 1, -8, -4, 0,
    -- layer=1 filter=168 channel=123
    -37, 4, 41, -14, 3, 18, -8, -2, 17,
    -- layer=1 filter=168 channel=124
    3, -3, -2, 3, 0, 17, 2, 3, 16,
    -- layer=1 filter=168 channel=125
    23, 29, 31, 57, 20, 37, 32, 17, 9,
    -- layer=1 filter=168 channel=126
    -5, -20, -9, 11, 0, 15, 1, -6, 4,
    -- layer=1 filter=168 channel=127
    -11, 23, 4, -2, -8, -39, -9, -17, -9,
    -- layer=1 filter=169 channel=0
    1, 1, 1, 3, 1, 1, -10, 3, -4,
    -- layer=1 filter=169 channel=1
    7, 5, 1, 6, 6, 2, 6, -8, 4,
    -- layer=1 filter=169 channel=2
    0, 4, 0, -9, 0, -3, 0, -11, -11,
    -- layer=1 filter=169 channel=3
    -4, 2, -2, -3, 2, 0, 0, -7, -9,
    -- layer=1 filter=169 channel=4
    0, 2, 3, 5, 1, -11, 2, -6, 6,
    -- layer=1 filter=169 channel=5
    -4, 1, 5, -14, -4, 8, -4, 8, -6,
    -- layer=1 filter=169 channel=6
    -3, 1, -9, 2, -9, 0, -9, 6, 3,
    -- layer=1 filter=169 channel=7
    7, -14, 10, -13, 5, -9, 7, -11, -12,
    -- layer=1 filter=169 channel=8
    -4, -11, 0, -6, -9, 7, -1, -11, 0,
    -- layer=1 filter=169 channel=9
    -9, -8, 6, 8, 2, 1, 3, -9, -6,
    -- layer=1 filter=169 channel=10
    -8, 0, -9, -10, -8, -10, -12, 2, -1,
    -- layer=1 filter=169 channel=11
    8, -10, -10, 1, -2, -9, -1, 2, -8,
    -- layer=1 filter=169 channel=12
    -5, 1, 3, -6, -1, 2, -6, -2, -10,
    -- layer=1 filter=169 channel=13
    -2, -6, -4, -1, 5, -10, 5, -12, 7,
    -- layer=1 filter=169 channel=14
    -6, 2, 7, -6, 2, -3, 4, -6, -3,
    -- layer=1 filter=169 channel=15
    -11, -9, -5, 2, -8, -7, -1, 5, 2,
    -- layer=1 filter=169 channel=16
    -5, 2, 6, 1, -6, 1, -10, 0, 6,
    -- layer=1 filter=169 channel=17
    0, -1, 8, -11, 6, 1, -12, 6, -12,
    -- layer=1 filter=169 channel=18
    0, -5, -11, 8, 0, -1, 3, 5, -8,
    -- layer=1 filter=169 channel=19
    1, 5, 5, 5, 2, 5, -5, -5, 7,
    -- layer=1 filter=169 channel=20
    4, 1, -1, 1, 3, -9, -7, -3, -9,
    -- layer=1 filter=169 channel=21
    -4, -1, 7, 6, 1, -2, -3, 8, -6,
    -- layer=1 filter=169 channel=22
    -11, -9, 7, -2, -9, -9, 3, 5, 8,
    -- layer=1 filter=169 channel=23
    -1, -8, 0, -11, -10, -3, -1, -10, 7,
    -- layer=1 filter=169 channel=24
    6, -1, 7, -7, -2, 7, -7, -8, 5,
    -- layer=1 filter=169 channel=25
    8, 0, 1, -1, -1, -10, -11, -2, -12,
    -- layer=1 filter=169 channel=26
    -10, -12, 1, 4, -5, -3, 0, -1, -10,
    -- layer=1 filter=169 channel=27
    -1, 4, 4, 0, 6, -12, -14, 0, -9,
    -- layer=1 filter=169 channel=28
    6, 0, -11, 2, -2, -1, 5, -2, -1,
    -- layer=1 filter=169 channel=29
    -7, 1, -10, -11, 4, 6, 7, 0, 8,
    -- layer=1 filter=169 channel=30
    2, -9, -2, 2, -1, -3, -3, -8, -10,
    -- layer=1 filter=169 channel=31
    6, 5, -1, -12, -9, 3, -11, 2, 8,
    -- layer=1 filter=169 channel=32
    1, -6, -2, 0, -1, -11, -4, -4, -3,
    -- layer=1 filter=169 channel=33
    0, 0, -5, -5, -8, 6, 7, 11, -2,
    -- layer=1 filter=169 channel=34
    6, -1, 7, -2, -4, 4, 1, 8, 7,
    -- layer=1 filter=169 channel=35
    1, -8, -11, -6, 6, 6, 2, 2, 3,
    -- layer=1 filter=169 channel=36
    0, 4, 2, 8, -8, 9, -1, 7, 4,
    -- layer=1 filter=169 channel=37
    -3, -10, -5, 1, 3, 3, -3, -8, -2,
    -- layer=1 filter=169 channel=38
    -2, -7, 6, -12, -13, 7, 1, 6, -8,
    -- layer=1 filter=169 channel=39
    3, -8, -11, 6, 2, 0, -1, -2, 6,
    -- layer=1 filter=169 channel=40
    -11, 4, 1, -9, 1, 0, 3, -5, -3,
    -- layer=1 filter=169 channel=41
    7, 4, 1, -10, 7, 5, 7, 0, 8,
    -- layer=1 filter=169 channel=42
    -16, 4, 3, -2, 2, 0, -7, -9, 6,
    -- layer=1 filter=169 channel=43
    -5, -11, 0, -9, 0, 5, -2, -8, -9,
    -- layer=1 filter=169 channel=44
    7, 1, -10, -12, 2, -9, 1, 1, -11,
    -- layer=1 filter=169 channel=45
    4, -11, 5, 6, -8, -12, -2, 0, 2,
    -- layer=1 filter=169 channel=46
    -11, -8, -8, -6, -4, 0, -7, 0, 2,
    -- layer=1 filter=169 channel=47
    -7, -7, 2, 0, -1, 2, -6, -6, -10,
    -- layer=1 filter=169 channel=48
    -1, -9, -8, -8, -8, -10, -5, -4, 1,
    -- layer=1 filter=169 channel=49
    8, -7, -11, -3, 7, 3, 0, 3, -4,
    -- layer=1 filter=169 channel=50
    -7, -7, 0, -2, 3, 0, 4, 0, 3,
    -- layer=1 filter=169 channel=51
    0, 6, 4, -9, -9, 0, -5, -12, -4,
    -- layer=1 filter=169 channel=52
    0, -1, -11, -11, 3, 7, -7, -11, -1,
    -- layer=1 filter=169 channel=53
    -11, 3, 2, 8, -6, -3, 0, -2, -9,
    -- layer=1 filter=169 channel=54
    2, 5, -1, -11, -12, -11, -1, 2, 0,
    -- layer=1 filter=169 channel=55
    -13, 0, -15, 3, 3, 0, -4, -7, -7,
    -- layer=1 filter=169 channel=56
    6, -7, 5, -10, 3, -2, 6, 7, -10,
    -- layer=1 filter=169 channel=57
    6, 3, 6, -6, -4, 0, 1, 0, 5,
    -- layer=1 filter=169 channel=58
    -2, 1, -1, -1, 2, -5, -3, -12, 4,
    -- layer=1 filter=169 channel=59
    -6, 5, -4, -7, -4, -2, -7, -5, 6,
    -- layer=1 filter=169 channel=60
    -6, 2, 5, 1, -10, 0, -1, -2, 0,
    -- layer=1 filter=169 channel=61
    7, -6, 2, 6, -4, -11, 2, -4, 3,
    -- layer=1 filter=169 channel=62
    5, 6, 4, -14, 0, 4, 0, -4, -2,
    -- layer=1 filter=169 channel=63
    8, -10, 3, -7, 2, -2, 0, 2, -4,
    -- layer=1 filter=169 channel=64
    8, -11, -2, 4, 0, 8, -7, -7, -3,
    -- layer=1 filter=169 channel=65
    5, -8, -10, -6, 8, 1, 7, -11, -5,
    -- layer=1 filter=169 channel=66
    0, 7, 1, -7, -8, 4, -12, 4, 0,
    -- layer=1 filter=169 channel=67
    -1, 2, 4, -3, -6, -8, 9, 8, -8,
    -- layer=1 filter=169 channel=68
    -3, 3, -10, -6, -1, -1, -7, -4, -9,
    -- layer=1 filter=169 channel=69
    3, 0, -17, -3, -5, -1, -1, 7, -12,
    -- layer=1 filter=169 channel=70
    3, -9, 0, 3, -6, -5, -11, 3, 4,
    -- layer=1 filter=169 channel=71
    6, 4, -6, 0, -10, 1, 2, 6, 4,
    -- layer=1 filter=169 channel=72
    7, -6, 6, 2, -4, -8, -7, -1, 5,
    -- layer=1 filter=169 channel=73
    5, -3, 1, 0, -8, -1, -11, -5, -10,
    -- layer=1 filter=169 channel=74
    2, 0, 5, -8, -10, -2, 1, -11, 2,
    -- layer=1 filter=169 channel=75
    -5, -4, 1, -1, -1, -8, -3, -8, 0,
    -- layer=1 filter=169 channel=76
    -5, 5, -2, 2, 3, -5, -1, -5, -7,
    -- layer=1 filter=169 channel=77
    7, -2, 6, -8, -2, 2, -10, -5, -1,
    -- layer=1 filter=169 channel=78
    6, 3, 6, -4, -11, -11, -11, -11, 0,
    -- layer=1 filter=169 channel=79
    -3, 4, 1, -2, -6, -8, 1, -1, -13,
    -- layer=1 filter=169 channel=80
    -8, -9, 6, -1, 8, 1, -1, 9, -8,
    -- layer=1 filter=169 channel=81
    -8, -3, -9, -6, -7, 4, -9, -11, 5,
    -- layer=1 filter=169 channel=82
    -9, 1, 5, -9, -8, 5, -5, 2, 5,
    -- layer=1 filter=169 channel=83
    -7, -2, -12, -10, -2, 3, -1, -3, 4,
    -- layer=1 filter=169 channel=84
    0, -1, -12, -12, -3, -4, 5, -11, 2,
    -- layer=1 filter=169 channel=85
    -5, 3, -11, -12, -8, -6, -6, -4, -2,
    -- layer=1 filter=169 channel=86
    2, -8, 4, -8, 6, 0, -6, 0, 1,
    -- layer=1 filter=169 channel=87
    8, 8, 0, 8, 4, 3, 3, 5, 5,
    -- layer=1 filter=169 channel=88
    0, 5, 5, -4, 3, 4, -8, -5, -2,
    -- layer=1 filter=169 channel=89
    -10, 1, -3, -10, -9, 7, -4, 7, 8,
    -- layer=1 filter=169 channel=90
    -2, 4, 6, 6, 0, -2, -1, -7, 8,
    -- layer=1 filter=169 channel=91
    -11, -1, 6, -1, -5, 6, -3, 1, 3,
    -- layer=1 filter=169 channel=92
    -11, 0, -7, -8, 0, -11, -3, 0, -2,
    -- layer=1 filter=169 channel=93
    7, -4, -8, 6, -9, 0, -11, -2, -1,
    -- layer=1 filter=169 channel=94
    1, 3, 6, -9, 5, -6, 1, -9, -10,
    -- layer=1 filter=169 channel=95
    4, -13, 4, -3, 0, -10, -3, 4, 8,
    -- layer=1 filter=169 channel=96
    0, 7, -6, 7, -4, -11, 0, -3, -8,
    -- layer=1 filter=169 channel=97
    -3, -3, 3, -3, -4, -8, -10, 4, -9,
    -- layer=1 filter=169 channel=98
    -5, 0, -5, -4, -1, 0, -10, 5, -4,
    -- layer=1 filter=169 channel=99
    7, 3, 2, -7, -11, -7, -9, 3, 1,
    -- layer=1 filter=169 channel=100
    -11, -4, -5, -5, -6, -11, 1, 0, 4,
    -- layer=1 filter=169 channel=101
    -6, -12, -12, -2, -5, 6, 1, 3, -6,
    -- layer=1 filter=169 channel=102
    -10, -1, -8, 0, -4, -10, -2, -4, -10,
    -- layer=1 filter=169 channel=103
    2, -4, -10, -9, -5, -5, 0, -7, 5,
    -- layer=1 filter=169 channel=104
    5, -10, -12, 5, 9, 7, 8, 2, 5,
    -- layer=1 filter=169 channel=105
    -8, 7, -7, 2, 4, 0, -10, -10, -3,
    -- layer=1 filter=169 channel=106
    -3, -11, 7, -2, -2, 2, 0, -5, 3,
    -- layer=1 filter=169 channel=107
    -2, 2, 2, 6, -6, 0, -4, 3, 1,
    -- layer=1 filter=169 channel=108
    3, -15, -1, 0, 3, -5, -3, -6, -5,
    -- layer=1 filter=169 channel=109
    -8, -6, -1, 7, 3, 1, -4, -2, 8,
    -- layer=1 filter=169 channel=110
    0, -3, -3, -10, 8, 3, 1, 2, -12,
    -- layer=1 filter=169 channel=111
    -5, -12, -5, 1, 2, -7, 0, -7, 3,
    -- layer=1 filter=169 channel=112
    -8, -11, 5, 7, -11, -7, -7, -11, 8,
    -- layer=1 filter=169 channel=113
    -2, 6, 4, 4, 1, 5, -10, -1, -8,
    -- layer=1 filter=169 channel=114
    -1, -8, -4, -11, -2, -7, -8, -2, -3,
    -- layer=1 filter=169 channel=115
    8, -6, -1, -11, 1, 6, 1, 3, -6,
    -- layer=1 filter=169 channel=116
    -5, 3, 9, -7, 5, -1, 9, -3, 7,
    -- layer=1 filter=169 channel=117
    -9, -3, 4, 6, 6, 4, 4, -3, 3,
    -- layer=1 filter=169 channel=118
    3, -5, 0, -8, 4, -8, 2, -11, 2,
    -- layer=1 filter=169 channel=119
    0, 5, 5, 0, 5, 0, 2, 0, -1,
    -- layer=1 filter=169 channel=120
    -5, 7, -9, -11, -11, -12, -2, 6, -4,
    -- layer=1 filter=169 channel=121
    -18, 0, -9, -11, -4, -15, -13, -8, -3,
    -- layer=1 filter=169 channel=122
    7, 8, 1, -3, -10, 7, -10, -1, -4,
    -- layer=1 filter=169 channel=123
    -12, -11, 3, 3, 0, 7, 1, 0, -1,
    -- layer=1 filter=169 channel=124
    7, -11, 2, -7, 2, 0, -9, 0, 3,
    -- layer=1 filter=169 channel=125
    0, 0, -1, -11, -7, -9, 3, 0, -6,
    -- layer=1 filter=169 channel=126
    1, -3, 0, -1, -9, -10, 4, 6, 0,
    -- layer=1 filter=169 channel=127
    0, -8, 2, -9, -6, -6, 4, 3, -3,
    -- layer=1 filter=170 channel=0
    14, 17, 11, 12, 5, -3, -4, -12, -12,
    -- layer=1 filter=170 channel=1
    39, 1, -3, -34, -11, -2, 16, -1, 7,
    -- layer=1 filter=170 channel=2
    -13, -5, 16, 14, -10, -4, 39, 3, 15,
    -- layer=1 filter=170 channel=3
    -8, -13, 7, -1, -8, -5, -5, 0, 12,
    -- layer=1 filter=170 channel=4
    0, 4, -7, 0, 5, -1, 0, -2, 0,
    -- layer=1 filter=170 channel=5
    36, -9, -3, -33, -25, -20, 4, -17, 3,
    -- layer=1 filter=170 channel=6
    2, -6, 11, 6, 0, 3, 3, 10, 22,
    -- layer=1 filter=170 channel=7
    -21, 6, -11, -2, 19, -6, 29, -1, 8,
    -- layer=1 filter=170 channel=8
    24, -3, 2, -33, -19, -34, 4, -2, 10,
    -- layer=1 filter=170 channel=9
    4, 31, -8, 47, -3, 40, 0, 7, 0,
    -- layer=1 filter=170 channel=10
    -18, 8, -5, 5, 9, 8, 24, 5, 10,
    -- layer=1 filter=170 channel=11
    18, 15, 3, -3, 8, 5, -12, -20, -19,
    -- layer=1 filter=170 channel=12
    -1, 0, -17, -22, -35, -29, 3, 7, 41,
    -- layer=1 filter=170 channel=13
    -18, -11, -11, -1, 0, 11, -9, 0, -2,
    -- layer=1 filter=170 channel=14
    -31, -15, -11, -23, 23, -24, -3, -8, 3,
    -- layer=1 filter=170 channel=15
    0, 0, -8, -61, -32, -14, 8, 6, 8,
    -- layer=1 filter=170 channel=16
    17, -12, -19, -18, -20, -12, -4, 1, 1,
    -- layer=1 filter=170 channel=17
    12, 0, 22, -12, -18, -19, -17, -15, -10,
    -- layer=1 filter=170 channel=18
    3, -2, 4, 15, -1, 13, -15, -12, -12,
    -- layer=1 filter=170 channel=19
    38, 65, 0, 63, 28, 35, 34, 54, 9,
    -- layer=1 filter=170 channel=20
    1, -2, 11, -24, 0, -2, -4, -1, 9,
    -- layer=1 filter=170 channel=21
    -4, -19, -7, -28, 5, -2, 1, 0, 0,
    -- layer=1 filter=170 channel=22
    -6, 11, 15, -20, -5, -12, -14, 3, -13,
    -- layer=1 filter=170 channel=23
    -5, 37, -9, 4, -33, 1, 20, 0, 11,
    -- layer=1 filter=170 channel=24
    0, -3, -15, -3, -22, -14, -15, 6, -3,
    -- layer=1 filter=170 channel=25
    2, 2, 1, 0, 13, 15, 34, 14, 21,
    -- layer=1 filter=170 channel=26
    -12, 3, 0, 19, 0, 6, -8, -2, 2,
    -- layer=1 filter=170 channel=27
    57, 52, 39, 19, 2, 1, -27, -32, -21,
    -- layer=1 filter=170 channel=28
    -14, 19, 10, -13, 10, -2, 4, 8, 5,
    -- layer=1 filter=170 channel=29
    31, 0, 13, -11, -5, 5, -23, -16, -20,
    -- layer=1 filter=170 channel=30
    -1, 6, -14, 24, -2, 16, -3, 8, -14,
    -- layer=1 filter=170 channel=31
    -3, 3, 6, -6, -3, -10, -16, 0, 7,
    -- layer=1 filter=170 channel=32
    0, 8, -6, 30, -4, 21, 9, 18, 1,
    -- layer=1 filter=170 channel=33
    8, 19, 6, 10, 3, -1, -2, -18, 0,
    -- layer=1 filter=170 channel=34
    -11, 9, 13, 1, 10, -16, 15, 0, -14,
    -- layer=1 filter=170 channel=35
    -9, 2, 3, -4, -1, -11, -13, -8, 1,
    -- layer=1 filter=170 channel=36
    9, 20, 1, 4, 7, -5, -14, -26, -24,
    -- layer=1 filter=170 channel=37
    35, -11, -21, -19, -3, -13, 0, -12, 7,
    -- layer=1 filter=170 channel=38
    -21, -3, 1, -9, 1, 6, -2, 0, 5,
    -- layer=1 filter=170 channel=39
    23, 18, 6, 10, 7, -10, -22, -2, -10,
    -- layer=1 filter=170 channel=40
    -2, -5, 8, 7, 7, 0, -4, -5, -4,
    -- layer=1 filter=170 channel=41
    -13, 33, -35, 53, -9, 50, -14, 40, -7,
    -- layer=1 filter=170 channel=42
    -41, -24, -5, -7, -3, -9, 10, 9, 24,
    -- layer=1 filter=170 channel=43
    26, 19, 0, -28, -14, -7, 30, 7, 11,
    -- layer=1 filter=170 channel=44
    -10, 9, -1, 4, 4, 11, -3, 4, 17,
    -- layer=1 filter=170 channel=45
    -18, -9, -5, -23, -17, -3, -14, 0, -2,
    -- layer=1 filter=170 channel=46
    49, 42, 0, 3, -12, -18, 12, 19, 9,
    -- layer=1 filter=170 channel=47
    -30, 0, -14, 36, -7, 48, 14, 25, 26,
    -- layer=1 filter=170 channel=48
    -9, 2, 0, -1, -10, 3, -9, 3, -6,
    -- layer=1 filter=170 channel=49
    -7, 3, 0, 14, 1, 6, 6, 8, -4,
    -- layer=1 filter=170 channel=50
    4, 5, 14, 16, 7, 4, -6, 0, 0,
    -- layer=1 filter=170 channel=51
    -7, 1, -4, 0, 0, 12, 11, -7, 6,
    -- layer=1 filter=170 channel=52
    -5, 0, -8, 1, 3, -7, 12, 14, 9,
    -- layer=1 filter=170 channel=53
    -1, -14, 0, -18, 0, -10, -11, -1, 11,
    -- layer=1 filter=170 channel=54
    17, 0, -11, 11, 21, 8, 35, 25, 23,
    -- layer=1 filter=170 channel=55
    20, 20, 6, 19, 1, -17, -13, -6, 0,
    -- layer=1 filter=170 channel=56
    5, -8, -10, 7, -3, -1, -3, 10, 3,
    -- layer=1 filter=170 channel=57
    -9, 17, -2, -6, 7, 11, 9, 4, 9,
    -- layer=1 filter=170 channel=58
    0, 17, -1, 42, -10, 16, 26, 23, 24,
    -- layer=1 filter=170 channel=59
    -9, 8, 4, -6, 4, -9, -5, -4, 4,
    -- layer=1 filter=170 channel=60
    0, 5, 7, 22, 3, 11, 4, -3, 26,
    -- layer=1 filter=170 channel=61
    0, 1, 0, 6, 0, 0, -6, -4, -8,
    -- layer=1 filter=170 channel=62
    17, -4, -19, -24, -13, -31, 9, -5, 3,
    -- layer=1 filter=170 channel=63
    21, 15, -4, 14, 4, 0, -13, -25, -29,
    -- layer=1 filter=170 channel=64
    9, 4, 6, -12, 7, -11, -8, -9, 1,
    -- layer=1 filter=170 channel=65
    8, 12, 0, -2, 10, 10, 4, -7, -12,
    -- layer=1 filter=170 channel=66
    20, 9, 4, -2, -3, -6, -14, -20, -13,
    -- layer=1 filter=170 channel=67
    15, 12, 6, 12, 17, 9, 25, 28, 16,
    -- layer=1 filter=170 channel=68
    1, -5, -9, 16, 1, 29, -4, 10, 24,
    -- layer=1 filter=170 channel=69
    -3, -18, -20, -20, -26, -27, 1, 8, 13,
    -- layer=1 filter=170 channel=70
    16, 7, 0, 3, 1, 2, 21, 12, 8,
    -- layer=1 filter=170 channel=71
    20, 14, 5, -20, -13, -22, 0, -6, -1,
    -- layer=1 filter=170 channel=72
    11, 24, -16, 53, 5, 33, 9, 15, -13,
    -- layer=1 filter=170 channel=73
    0, 7, 7, 11, 6, -4, 1, -4, -12,
    -- layer=1 filter=170 channel=74
    9, -5, -3, 1, -16, 28, -23, 10, 30,
    -- layer=1 filter=170 channel=75
    -35, -28, -9, -29, -17, -18, -17, -30, 17,
    -- layer=1 filter=170 channel=76
    5, 6, -4, 19, -5, 16, -6, -21, -9,
    -- layer=1 filter=170 channel=77
    2, 5, 0, -21, 0, 1, -11, -8, 3,
    -- layer=1 filter=170 channel=78
    2, 7, 2, -5, 7, 1, -13, 4, 5,
    -- layer=1 filter=170 channel=79
    13, 0, -15, -3, -12, -30, 8, -8, 15,
    -- layer=1 filter=170 channel=80
    -3, 0, -4, 6, -6, -2, 2, 0, -3,
    -- layer=1 filter=170 channel=81
    10, 30, 12, -12, -28, -15, -23, -21, -25,
    -- layer=1 filter=170 channel=82
    1, -3, 6, -19, 1, -4, 1, -2, -7,
    -- layer=1 filter=170 channel=83
    15, -3, -7, -20, -19, -17, -10, -14, 11,
    -- layer=1 filter=170 channel=84
    31, 6, 26, 56, 27, 39, 4, 9, 28,
    -- layer=1 filter=170 channel=85
    -10, 36, -2, 19, -15, 5, 7, 14, 14,
    -- layer=1 filter=170 channel=86
    18, 10, 2, 1, -9, -14, -26, -28, -4,
    -- layer=1 filter=170 channel=87
    11, 43, -37, 66, -3, 13, 5, 47, 8,
    -- layer=1 filter=170 channel=88
    -9, 4, -6, 5, -6, 7, 9, 5, -13,
    -- layer=1 filter=170 channel=89
    -7, 8, 8, 8, 2, 4, 3, 3, 1,
    -- layer=1 filter=170 channel=90
    -16, -1, 0, 0, -13, 15, -16, 7, 9,
    -- layer=1 filter=170 channel=91
    -21, 3, 9, 2, -7, 14, 1, 3, 3,
    -- layer=1 filter=170 channel=92
    -33, 35, -4, 1, -6, 43, -27, 12, 38,
    -- layer=1 filter=170 channel=93
    -4, 4, -2, -12, 3, -5, -11, -7, -9,
    -- layer=1 filter=170 channel=94
    12, -1, 4, 3, 1, 6, -21, -14, -17,
    -- layer=1 filter=170 channel=95
    22, 10, 19, 36, 17, 33, 0, 14, 21,
    -- layer=1 filter=170 channel=96
    14, 5, 3, -9, 0, 3, 5, -8, 3,
    -- layer=1 filter=170 channel=97
    5, 3, 19, -1, 5, -19, -18, -15, -1,
    -- layer=1 filter=170 channel=98
    22, 12, 3, -19, -7, -13, 11, 13, 10,
    -- layer=1 filter=170 channel=99
    -8, -7, -11, -2, 20, 7, -21, 14, 0,
    -- layer=1 filter=170 channel=100
    24, 2, 2, 0, -2, -1, -16, -22, -9,
    -- layer=1 filter=170 channel=101
    -11, -11, 1, -1, -3, 0, -14, 9, 3,
    -- layer=1 filter=170 channel=102
    -8, 4, 13, 0, -8, 14, -22, -23, -22,
    -- layer=1 filter=170 channel=103
    30, 27, 16, 10, 7, 21, -10, -3, 2,
    -- layer=1 filter=170 channel=104
    -17, 15, -7, -3, -7, -6, 25, 20, 22,
    -- layer=1 filter=170 channel=105
    -2, 13, 16, -1, 0, -12, -19, -20, -21,
    -- layer=1 filter=170 channel=106
    -1, -7, 4, 11, 0, 7, -14, 0, 11,
    -- layer=1 filter=170 channel=107
    -15, -8, -11, -20, -21, -1, 2, -8, -11,
    -- layer=1 filter=170 channel=108
    -14, -10, -13, 12, -5, -9, 1, 25, -7,
    -- layer=1 filter=170 channel=109
    6, -10, -6, -4, -3, 0, -8, -2, 5,
    -- layer=1 filter=170 channel=110
    4, -2, -5, -4, -2, 1, -8, -3, -14,
    -- layer=1 filter=170 channel=111
    6, -3, 0, 39, -13, 17, 1, 0, 1,
    -- layer=1 filter=170 channel=112
    15, -6, 1, 8, 22, -8, 7, 6, 21,
    -- layer=1 filter=170 channel=113
    -6, 10, 1, -23, 16, 5, -1, -4, -5,
    -- layer=1 filter=170 channel=114
    18, -13, -11, -35, -38, -23, 0, -9, -21,
    -- layer=1 filter=170 channel=115
    9, 25, 6, -15, -6, -5, 0, -24, -2,
    -- layer=1 filter=170 channel=116
    -1, 1, -13, 3, -1, 7, 7, 5, 5,
    -- layer=1 filter=170 channel=117
    23, 0, 17, 50, 21, -2, 22, 15, 33,
    -- layer=1 filter=170 channel=118
    15, -1, 10, 21, 5, 19, -8, 1, 4,
    -- layer=1 filter=170 channel=119
    -2, 4, -3, 31, 5, 32, 6, 12, 2,
    -- layer=1 filter=170 channel=120
    -11, 3, -13, -8, -11, -1, -1, -6, 15,
    -- layer=1 filter=170 channel=121
    17, 0, -3, -25, -26, -20, -18, 1, -19,
    -- layer=1 filter=170 channel=122
    -1, 4, 8, 0, 1, 2, -2, 1, 0,
    -- layer=1 filter=170 channel=123
    10, 28, 0, -6, -4, -21, -10, -1, -5,
    -- layer=1 filter=170 channel=124
    -5, 6, -9, -11, -12, -4, 12, 7, -1,
    -- layer=1 filter=170 channel=125
    3, 0, -12, 2, 8, 5, -14, -2, -6,
    -- layer=1 filter=170 channel=126
    32, 10, -4, -20, -11, -19, 13, 28, 11,
    -- layer=1 filter=170 channel=127
    8, -6, -1, 24, 12, 23, 1, 16, 5,
    -- layer=1 filter=171 channel=0
    8, 0, 0, -6, 3, 5, 0, 2, -2,
    -- layer=1 filter=171 channel=1
    -6, -4, 8, 7, 7, -4, -10, -9, -9,
    -- layer=1 filter=171 channel=2
    -1, -10, 0, -10, 5, 2, -11, -10, 7,
    -- layer=1 filter=171 channel=3
    7, 4, 7, -4, -7, 3, -1, -2, -10,
    -- layer=1 filter=171 channel=4
    -6, -1, 5, 1, 6, -10, -4, -1, -9,
    -- layer=1 filter=171 channel=5
    -9, -9, 0, -4, -5, 2, 0, 3, -10,
    -- layer=1 filter=171 channel=6
    -6, -8, -10, -11, 0, -8, -9, 6, -2,
    -- layer=1 filter=171 channel=7
    -11, -7, -10, -1, 5, -9, -6, -3, -6,
    -- layer=1 filter=171 channel=8
    4, 0, -1, -9, 0, 0, -4, 0, -3,
    -- layer=1 filter=171 channel=9
    -9, -6, -11, 8, -11, 6, -1, 6, -12,
    -- layer=1 filter=171 channel=10
    4, -3, -9, -5, -6, -6, -13, 0, 6,
    -- layer=1 filter=171 channel=11
    0, 0, 8, -11, 5, -1, 5, 4, -11,
    -- layer=1 filter=171 channel=12
    -9, 2, 10, 0, 9, 8, -7, 2, 1,
    -- layer=1 filter=171 channel=13
    -3, -6, -4, 0, 6, -11, -2, 5, 10,
    -- layer=1 filter=171 channel=14
    -4, 8, 4, 0, 3, -1, 1, 5, -6,
    -- layer=1 filter=171 channel=15
    -2, 2, 4, -2, -4, -9, 1, -11, -3,
    -- layer=1 filter=171 channel=16
    -10, 5, 1, 0, -2, -5, 2, -8, -1,
    -- layer=1 filter=171 channel=17
    3, 4, -2, 0, 4, -11, 8, 2, 5,
    -- layer=1 filter=171 channel=18
    0, -4, -10, 0, 8, 2, 3, 0, -11,
    -- layer=1 filter=171 channel=19
    -1, -7, 5, 4, -2, 4, -1, -2, 0,
    -- layer=1 filter=171 channel=20
    -5, -5, -3, 2, -11, -9, 8, -12, -1,
    -- layer=1 filter=171 channel=21
    3, 5, 4, -3, -7, 0, -3, -4, 0,
    -- layer=1 filter=171 channel=22
    -3, -9, -1, 3, -10, 4, 0, -2, -9,
    -- layer=1 filter=171 channel=23
    -6, 5, 0, 6, 4, 3, 0, -7, -4,
    -- layer=1 filter=171 channel=24
    5, -2, -12, 5, -10, -3, -10, -2, -5,
    -- layer=1 filter=171 channel=25
    -5, -2, 11, -8, -10, -5, 9, 6, -10,
    -- layer=1 filter=171 channel=26
    -1, -5, 1, 7, 0, -5, -1, 7, 0,
    -- layer=1 filter=171 channel=27
    1, -3, 2, 2, -2, 4, -6, -3, -2,
    -- layer=1 filter=171 channel=28
    5, 1, 7, 0, -1, 4, -2, 3, -8,
    -- layer=1 filter=171 channel=29
    6, -8, 1, 2, 2, 2, -3, -12, -3,
    -- layer=1 filter=171 channel=30
    -10, -3, 0, -10, 1, -5, 5, 7, 3,
    -- layer=1 filter=171 channel=31
    4, -7, 6, -9, 2, 3, -3, 1, -2,
    -- layer=1 filter=171 channel=32
    2, 1, -1, 0, 3, -9, -8, -6, 5,
    -- layer=1 filter=171 channel=33
    10, -6, 6, 8, 5, -5, 8, 6, 7,
    -- layer=1 filter=171 channel=34
    -11, 7, -6, -2, -10, -3, 1, 4, 2,
    -- layer=1 filter=171 channel=35
    -7, -5, -10, 4, 0, -9, 8, -10, 5,
    -- layer=1 filter=171 channel=36
    7, 4, -2, -10, -2, 3, 3, -10, -2,
    -- layer=1 filter=171 channel=37
    -5, -11, 7, -1, 4, 6, 3, -13, -1,
    -- layer=1 filter=171 channel=38
    1, -5, 10, 8, -6, 10, 2, -5, 4,
    -- layer=1 filter=171 channel=39
    -1, 3, -8, 3, -1, -11, -11, -5, -10,
    -- layer=1 filter=171 channel=40
    -6, -8, -6, -8, 5, 8, -3, -5, -1,
    -- layer=1 filter=171 channel=41
    0, 5, 7, -2, -8, 0, 4, -9, 1,
    -- layer=1 filter=171 channel=42
    -5, 4, 4, -5, 0, -5, 1, -6, -3,
    -- layer=1 filter=171 channel=43
    8, 0, 1, 0, -8, 4, 3, 4, -4,
    -- layer=1 filter=171 channel=44
    -11, -1, -1, 1, 0, 3, -9, 0, 2,
    -- layer=1 filter=171 channel=45
    0, -6, 3, -5, 1, -10, -1, -5, -3,
    -- layer=1 filter=171 channel=46
    5, -6, 5, -6, -4, 8, 6, 6, 4,
    -- layer=1 filter=171 channel=47
    -12, 0, -7, -5, 0, -1, -8, 4, -10,
    -- layer=1 filter=171 channel=48
    8, 3, -7, 4, -11, 3, -5, -5, -8,
    -- layer=1 filter=171 channel=49
    8, -6, 9, -3, 0, 3, -8, 0, 8,
    -- layer=1 filter=171 channel=50
    2, 5, 2, -3, 1, -4, -10, -5, -9,
    -- layer=1 filter=171 channel=51
    8, -8, -9, -4, -7, -11, 0, 5, -6,
    -- layer=1 filter=171 channel=52
    0, 6, 9, -2, -9, -6, 0, -1, 10,
    -- layer=1 filter=171 channel=53
    -4, 7, -2, 3, 1, -3, -1, -2, -3,
    -- layer=1 filter=171 channel=54
    6, 4, 0, -6, 1, 0, -13, -13, -3,
    -- layer=1 filter=171 channel=55
    2, 6, 1, 0, -1, 6, 3, -2, -3,
    -- layer=1 filter=171 channel=56
    8, 1, 2, 1, 2, -4, -10, 2, 2,
    -- layer=1 filter=171 channel=57
    2, 2, -6, 5, -2, 3, -9, -14, 1,
    -- layer=1 filter=171 channel=58
    2, 0, 5, -2, 5, 5, 2, -5, -10,
    -- layer=1 filter=171 channel=59
    -2, 0, -4, -9, 8, 0, -7, 0, -8,
    -- layer=1 filter=171 channel=60
    -8, -2, -4, 1, 5, 8, -7, 8, -8,
    -- layer=1 filter=171 channel=61
    8, -3, -7, -3, 6, -2, -8, -9, 4,
    -- layer=1 filter=171 channel=62
    -1, 5, -7, 6, -2, 0, -12, 2, 9,
    -- layer=1 filter=171 channel=63
    -4, 4, 0, -8, -4, -4, -6, 1, -11,
    -- layer=1 filter=171 channel=64
    -1, 0, -5, -3, 0, -5, -6, -7, 5,
    -- layer=1 filter=171 channel=65
    -2, -10, -2, -10, 0, 0, -4, 0, 5,
    -- layer=1 filter=171 channel=66
    1, -10, 8, 5, 4, -7, 4, -3, -6,
    -- layer=1 filter=171 channel=67
    4, 10, 0, 6, 0, -9, 3, -10, 6,
    -- layer=1 filter=171 channel=68
    -8, -4, 0, -11, 8, 7, 5, -10, 4,
    -- layer=1 filter=171 channel=69
    3, 9, 7, 7, -4, 1, 2, -11, -10,
    -- layer=1 filter=171 channel=70
    7, 11, 3, -7, -1, 2, 7, 5, 3,
    -- layer=1 filter=171 channel=71
    6, 10, -1, -4, 5, 6, -7, -7, 6,
    -- layer=1 filter=171 channel=72
    -11, 7, -10, -7, -5, -5, 7, 8, -6,
    -- layer=1 filter=171 channel=73
    -5, -9, 8, -12, 8, -10, -1, 6, 6,
    -- layer=1 filter=171 channel=74
    3, 2, 6, 6, 5, -3, -11, -6, 5,
    -- layer=1 filter=171 channel=75
    -7, 0, 1, 2, 0, 9, 5, 1, -11,
    -- layer=1 filter=171 channel=76
    1, -10, 2, -5, 6, 5, 0, -3, -5,
    -- layer=1 filter=171 channel=77
    -10, 7, -6, 0, -3, 5, -3, -3, -9,
    -- layer=1 filter=171 channel=78
    7, 5, 0, 7, -11, -6, 7, 4, 2,
    -- layer=1 filter=171 channel=79
    7, -6, -8, -10, 1, 3, -6, 5, 4,
    -- layer=1 filter=171 channel=80
    -5, -3, -4, -2, -3, 6, 8, 8, -9,
    -- layer=1 filter=171 channel=81
    -4, -3, 1, -6, -8, -4, -1, -8, -12,
    -- layer=1 filter=171 channel=82
    -4, -4, 0, -6, 6, -1, 0, 1, 3,
    -- layer=1 filter=171 channel=83
    -5, -8, -3, -12, 0, 1, -4, -6, 2,
    -- layer=1 filter=171 channel=84
    -4, -3, -5, -9, -4, 7, -9, -2, 3,
    -- layer=1 filter=171 channel=85
    2, 7, -7, 5, 2, 1, -3, -3, 4,
    -- layer=1 filter=171 channel=86
    5, 0, -1, -1, 1, -7, 1, -3, -11,
    -- layer=1 filter=171 channel=87
    -8, -4, 0, -11, -11, 8, -2, -9, -9,
    -- layer=1 filter=171 channel=88
    6, -4, -1, 0, -3, -10, -6, 4, 2,
    -- layer=1 filter=171 channel=89
    2, 7, -12, -6, 0, -1, -4, 5, 6,
    -- layer=1 filter=171 channel=90
    6, -8, 5, -2, -9, -11, 7, -7, -12,
    -- layer=1 filter=171 channel=91
    8, -4, -5, 2, -6, -7, -11, -5, -7,
    -- layer=1 filter=171 channel=92
    5, 1, 0, -6, -10, 5, -12, -4, 0,
    -- layer=1 filter=171 channel=93
    -2, 2, 1, -8, -1, -4, -7, -2, -11,
    -- layer=1 filter=171 channel=94
    -1, 2, -10, 6, -1, -3, 4, 2, 7,
    -- layer=1 filter=171 channel=95
    -4, 5, 6, -5, -5, 2, -4, -9, -2,
    -- layer=1 filter=171 channel=96
    -6, -6, -5, -10, 3, -10, 3, -7, -7,
    -- layer=1 filter=171 channel=97
    -5, -8, -7, -8, -7, 0, -11, -1, -8,
    -- layer=1 filter=171 channel=98
    -6, 9, -8, 7, 0, -8, -11, -5, -3,
    -- layer=1 filter=171 channel=99
    7, -5, 3, -3, -6, 0, 3, -2, -10,
    -- layer=1 filter=171 channel=100
    -4, 1, -11, -2, -11, -8, -6, 8, 1,
    -- layer=1 filter=171 channel=101
    -8, 3, -1, 5, -12, -4, -5, 0, 9,
    -- layer=1 filter=171 channel=102
    -12, -9, -1, 6, -3, -9, -2, 1, -2,
    -- layer=1 filter=171 channel=103
    8, -4, 6, -5, -6, -10, -6, 0, 7,
    -- layer=1 filter=171 channel=104
    -10, -6, 5, -7, 4, 3, 7, 7, 3,
    -- layer=1 filter=171 channel=105
    -4, -9, 1, -5, -5, -3, -3, -9, 0,
    -- layer=1 filter=171 channel=106
    -2, -8, -4, -7, 0, 5, -7, -3, -6,
    -- layer=1 filter=171 channel=107
    4, -11, 9, -6, -6, 4, -4, -3, -10,
    -- layer=1 filter=171 channel=108
    -8, 2, -4, -10, 0, -8, 9, -5, -5,
    -- layer=1 filter=171 channel=109
    -3, -9, -4, -3, 4, 7, 0, -8, 6,
    -- layer=1 filter=171 channel=110
    2, -4, 5, 5, -2, -6, -12, -7, -4,
    -- layer=1 filter=171 channel=111
    -5, -2, -1, 1, 6, -10, -7, 4, 6,
    -- layer=1 filter=171 channel=112
    -7, -9, 3, 5, 3, 2, -5, -8, -8,
    -- layer=1 filter=171 channel=113
    1, 8, -6, -9, -8, -2, -4, 4, -2,
    -- layer=1 filter=171 channel=114
    -4, -9, 6, -7, 0, -13, -8, -4, 1,
    -- layer=1 filter=171 channel=115
    -11, -7, -1, 2, 0, -10, 0, -8, 0,
    -- layer=1 filter=171 channel=116
    8, 4, 0, -8, -6, 6, 0, 9, 0,
    -- layer=1 filter=171 channel=117
    0, 7, 7, -1, -11, 8, -2, -10, 6,
    -- layer=1 filter=171 channel=118
    -1, 7, -7, -3, -2, 2, -6, 7, -5,
    -- layer=1 filter=171 channel=119
    4, -8, -12, -2, -7, -2, -5, -5, -10,
    -- layer=1 filter=171 channel=120
    -3, 8, 1, -10, -6, 6, 0, 6, 4,
    -- layer=1 filter=171 channel=121
    6, 4, -5, -8, -9, 4, -2, 2, -5,
    -- layer=1 filter=171 channel=122
    6, 5, -10, 0, 3, 9, -5, 0, 0,
    -- layer=1 filter=171 channel=123
    6, -12, 4, 3, 8, -8, -1, 4, 8,
    -- layer=1 filter=171 channel=124
    4, 8, -9, -5, 6, 2, -3, -6, -8,
    -- layer=1 filter=171 channel=125
    -8, 0, -3, -6, 5, -4, -8, 9, 3,
    -- layer=1 filter=171 channel=126
    0, 1, 3, 2, -8, -3, 1, 6, -4,
    -- layer=1 filter=171 channel=127
    -8, 4, 7, -2, 4, -10, 2, -3, -2,
    -- layer=1 filter=172 channel=0
    14, 7, 8, 12, 2, 4, -6, 7, 7,
    -- layer=1 filter=172 channel=1
    -18, -11, -5, 21, 23, -5, 9, 12, 13,
    -- layer=1 filter=172 channel=2
    -29, -46, -56, -54, -59, -67, 47, 66, 59,
    -- layer=1 filter=172 channel=3
    -14, 6, 9, 2, 7, 4, 7, -5, 3,
    -- layer=1 filter=172 channel=4
    1, 3, -8, -2, 3, 2, -8, -11, -1,
    -- layer=1 filter=172 channel=5
    2, 0, 13, -6, -6, -29, 4, 18, 6,
    -- layer=1 filter=172 channel=6
    -95, -77, -93, -6, 2, -1, 46, 30, 46,
    -- layer=1 filter=172 channel=7
    -15, -14, -33, -53, -96, -103, -43, -107, -43,
    -- layer=1 filter=172 channel=8
    14, 27, 18, 41, 24, 0, 0, 29, 22,
    -- layer=1 filter=172 channel=9
    18, 0, 1, 35, -18, -3, 15, -19, -30,
    -- layer=1 filter=172 channel=10
    -20, -48, -46, -81, -118, -91, -30, -91, -45,
    -- layer=1 filter=172 channel=11
    21, 20, 6, -3, 0, 0, -33, -13, 0,
    -- layer=1 filter=172 channel=12
    7, -30, 27, -7, -2, 8, 10, 29, 78,
    -- layer=1 filter=172 channel=13
    -28, -39, -25, 25, 10, 7, 42, 33, 33,
    -- layer=1 filter=172 channel=14
    -1, 0, 18, -26, -65, -78, -13, -28, -20,
    -- layer=1 filter=172 channel=15
    -6, -39, -45, -4, -2, -9, -10, -26, -4,
    -- layer=1 filter=172 channel=16
    32, 27, 28, 34, 26, 21, 21, 18, 16,
    -- layer=1 filter=172 channel=17
    8, 4, 0, 17, 11, -2, 10, 25, 15,
    -- layer=1 filter=172 channel=18
    16, -2, 11, 24, -20, -23, -23, -35, -6,
    -- layer=1 filter=172 channel=19
    45, 41, 18, 12, 12, 9, -2, -47, -44,
    -- layer=1 filter=172 channel=20
    -21, -29, -26, 24, 23, -2, 52, 44, 33,
    -- layer=1 filter=172 channel=21
    -24, -19, -38, 18, 5, -7, 28, 28, 14,
    -- layer=1 filter=172 channel=22
    -42, -26, -24, 32, 14, 2, 40, 32, 32,
    -- layer=1 filter=172 channel=23
    -19, 27, -26, -49, -36, -59, -74, -79, -47,
    -- layer=1 filter=172 channel=24
    16, -12, 2, -3, -17, 4, -25, -3, -7,
    -- layer=1 filter=172 channel=25
    -8, 5, -16, -7, -53, -43, -2, -46, -29,
    -- layer=1 filter=172 channel=26
    29, 22, 0, 10, 13, 6, 4, -3, 7,
    -- layer=1 filter=172 channel=27
    0, 13, 18, -39, -6, 3, -30, -18, -3,
    -- layer=1 filter=172 channel=28
    19, -27, -22, 14, -39, -43, -2, -38, -18,
    -- layer=1 filter=172 channel=29
    -15, 5, 5, -16, -12, -9, -47, -25, -25,
    -- layer=1 filter=172 channel=30
    59, 25, 5, -4, -23, -47, -9, -18, -12,
    -- layer=1 filter=172 channel=31
    -15, -37, -33, -12, -33, -27, 34, 41, 34,
    -- layer=1 filter=172 channel=32
    16, -7, -14, -34, -39, -63, -49, -34, -29,
    -- layer=1 filter=172 channel=33
    -15, 6, -4, -4, -7, -8, 0, -6, -14,
    -- layer=1 filter=172 channel=34
    -42, -20, -26, -8, 0, 28, 17, 1, -8,
    -- layer=1 filter=172 channel=35
    -4, 7, -3, -3, 0, 2, 7, 6, 1,
    -- layer=1 filter=172 channel=36
    38, 23, 33, 11, 1, 4, -13, -5, -9,
    -- layer=1 filter=172 channel=37
    9, 6, 3, -5, -9, -11, 0, 6, 4,
    -- layer=1 filter=172 channel=38
    -26, -27, -38, 1, 3, -7, 34, 41, 37,
    -- layer=1 filter=172 channel=39
    9, 16, 17, 21, 22, 8, -1, 10, 4,
    -- layer=1 filter=172 channel=40
    -45, -70, -42, 27, 0, 3, 30, 37, 42,
    -- layer=1 filter=172 channel=41
    68, 14, 9, 4, -53, -59, -67, -77, -33,
    -- layer=1 filter=172 channel=42
    -13, -35, -39, -47, -31, -72, 61, 81, 45,
    -- layer=1 filter=172 channel=43
    -2, 9, 4, 43, 14, 0, 13, 26, 10,
    -- layer=1 filter=172 channel=44
    23, -6, -12, -14, -7, -42, -47, -5, -10,
    -- layer=1 filter=172 channel=45
    -15, -33, -12, 7, -2, -5, 22, 32, 28,
    -- layer=1 filter=172 channel=46
    25, 29, 16, -8, 9, 7, 49, 14, 19,
    -- layer=1 filter=172 channel=47
    -35, -24, -29, -59, -56, -75, -31, -17, -21,
    -- layer=1 filter=172 channel=48
    -20, -10, -22, 7, 7, 2, 34, 18, 14,
    -- layer=1 filter=172 channel=49
    -40, -38, -42, -4, -7, -15, 50, 24, 37,
    -- layer=1 filter=172 channel=50
    -14, -9, 5, 8, 9, 10, 11, -9, 11,
    -- layer=1 filter=172 channel=51
    -40, -30, -33, -6, -15, -13, 16, 14, 9,
    -- layer=1 filter=172 channel=52
    -14, -2, 1, -1, -8, 7, 3, 9, 0,
    -- layer=1 filter=172 channel=53
    18, 2, 1, 6, 0, 9, 8, 9, 23,
    -- layer=1 filter=172 channel=54
    0, -8, -9, -36, -49, -22, -5, -57, -33,
    -- layer=1 filter=172 channel=55
    12, 17, 17, -14, 8, -1, -47, -25, -20,
    -- layer=1 filter=172 channel=56
    6, 6, -8, 4, -8, 1, 0, 4, 6,
    -- layer=1 filter=172 channel=57
    -52, -62, -73, -36, -71, -31, 0, -18, 16,
    -- layer=1 filter=172 channel=58
    -49, -43, -65, -129, -132, -144, -53, -127, -69,
    -- layer=1 filter=172 channel=59
    -15, -4, -8, -8, 8, -1, -6, 6, -3,
    -- layer=1 filter=172 channel=60
    12, -9, -4, 11, 5, 0, 4, 7, 0,
    -- layer=1 filter=172 channel=61
    0, -2, -8, 15, 3, -1, 7, 7, 3,
    -- layer=1 filter=172 channel=62
    6, 17, 7, 40, 19, 22, 2, 28, 31,
    -- layer=1 filter=172 channel=63
    16, 17, 20, -11, 0, 6, -26, -21, -9,
    -- layer=1 filter=172 channel=64
    -18, -16, -22, 11, -9, -12, 18, 17, 17,
    -- layer=1 filter=172 channel=65
    -11, -8, -26, 5, 5, 4, 26, 19, 18,
    -- layer=1 filter=172 channel=66
    11, 9, 16, -9, 1, 13, -12, -9, -6,
    -- layer=1 filter=172 channel=67
    -113, -92, -82, -62, -44, -40, 64, 48, 11,
    -- layer=1 filter=172 channel=68
    27, -13, 9, -34, -52, -51, -55, -37, -12,
    -- layer=1 filter=172 channel=69
    18, 13, 0, 3, 23, -2, -3, 15, 18,
    -- layer=1 filter=172 channel=70
    -64, -55, -67, -48, -53, -31, 86, 70, 72,
    -- layer=1 filter=172 channel=71
    -13, -6, -7, -7, -7, -19, -21, -10, -12,
    -- layer=1 filter=172 channel=72
    31, -12, -7, 15, -7, -44, -9, -51, -17,
    -- layer=1 filter=172 channel=73
    4, -13, -9, 2, 4, -4, -12, -3, 4,
    -- layer=1 filter=172 channel=74
    14, -10, 12, -3, -30, -30, -3, -33, -13,
    -- layer=1 filter=172 channel=75
    4, -3, -11, -13, -51, -59, -24, -20, 27,
    -- layer=1 filter=172 channel=76
    38, 20, 5, 4, -12, -6, -22, -13, -17,
    -- layer=1 filter=172 channel=77
    -25, -25, -30, 9, -7, -2, 8, 13, 4,
    -- layer=1 filter=172 channel=78
    6, 2, 5, 1, -11, -24, 14, -13, -14,
    -- layer=1 filter=172 channel=79
    23, 22, 10, 30, 26, 15, 18, 31, 30,
    -- layer=1 filter=172 channel=80
    -8, 4, 9, 5, 0, -9, -2, -8, -6,
    -- layer=1 filter=172 channel=81
    3, -2, -18, 10, 0, 13, -1, 3, 1,
    -- layer=1 filter=172 channel=82
    -29, -19, -28, 5, 4, -15, 26, 34, 29,
    -- layer=1 filter=172 channel=83
    3, -17, 0, 16, 3, -9, 12, 17, 18,
    -- layer=1 filter=172 channel=84
    30, 22, 28, 34, 8, -7, -22, -29, -1,
    -- layer=1 filter=172 channel=85
    -10, 2, -48, -41, -59, -61, -37, -63, -42,
    -- layer=1 filter=172 channel=86
    9, 18, 16, -15, -6, 3, -6, -3, -6,
    -- layer=1 filter=172 channel=87
    26, 3, -14, 12, 2, -16, 49, -3, -20,
    -- layer=1 filter=172 channel=88
    -15, -15, -2, 8, 1, 2, 33, 19, 30,
    -- layer=1 filter=172 channel=89
    -17, -12, -13, 17, -5, -3, 20, 37, 20,
    -- layer=1 filter=172 channel=90
    26, -17, -3, -3, -24, -36, -37, -23, -5,
    -- layer=1 filter=172 channel=91
    -22, -32, -41, 8, 5, 9, 37, 39, 34,
    -- layer=1 filter=172 channel=92
    28, -17, -6, -32, -56, -11, -4, -32, -58,
    -- layer=1 filter=172 channel=93
    -4, -3, -17, 16, 3, -4, 12, 0, 14,
    -- layer=1 filter=172 channel=94
    29, 5, 22, 9, 8, 18, -3, 7, -5,
    -- layer=1 filter=172 channel=95
    41, 26, 34, 2, -12, -7, -30, -22, -9,
    -- layer=1 filter=172 channel=96
    3, -4, -9, 4, 12, 0, 0, 8, -4,
    -- layer=1 filter=172 channel=97
    15, 12, 16, 14, 4, 9, -4, 13, 3,
    -- layer=1 filter=172 channel=98
    3, 0, 5, 42, 24, 16, 16, 21, 31,
    -- layer=1 filter=172 channel=99
    -12, -94, -5, -34, -111, -92, -5, -53, -73,
    -- layer=1 filter=172 channel=100
    25, 22, 30, -19, 4, 3, -19, -12, 3,
    -- layer=1 filter=172 channel=101
    -37, -30, -21, 11, 12, -10, 37, 47, 29,
    -- layer=1 filter=172 channel=102
    19, -4, 7, -5, 7, -5, 28, 12, 7,
    -- layer=1 filter=172 channel=103
    3, 15, 17, 1, 11, 18, -10, -8, 13,
    -- layer=1 filter=172 channel=104
    -4, 3, -30, -26, -1, -64, -39, -19, -17,
    -- layer=1 filter=172 channel=105
    16, 8, 12, 12, -8, 8, 2, -4, -4,
    -- layer=1 filter=172 channel=106
    -37, -28, -31, -5, 10, -12, 50, 36, 42,
    -- layer=1 filter=172 channel=107
    11, -6, 5, 0, -2, -1, 3, 11, 0,
    -- layer=1 filter=172 channel=108
    21, -3, -39, -11, -23, -40, -56, -31, -25,
    -- layer=1 filter=172 channel=109
    -4, 5, -3, -5, -8, 4, 0, -1, 3,
    -- layer=1 filter=172 channel=110
    -5, 3, 1, -7, -2, -8, -7, -2, 3,
    -- layer=1 filter=172 channel=111
    64, 26, 18, 8, -8, -8, -5, -12, -3,
    -- layer=1 filter=172 channel=112
    18, 25, 44, 41, 21, 33, -26, -15, -5,
    -- layer=1 filter=172 channel=113
    -60, -74, -71, -6, -41, -34, 18, 35, 4,
    -- layer=1 filter=172 channel=114
    19, 30, 22, 18, 17, 16, -12, 7, 11,
    -- layer=1 filter=172 channel=115
    10, -9, 5, 4, -5, -9, -7, -27, -16,
    -- layer=1 filter=172 channel=116
    2, -10, -8, -7, -3, 0, -2, -9, -3,
    -- layer=1 filter=172 channel=117
    40, 16, 53, 53, 31, 43, -11, -3, 4,
    -- layer=1 filter=172 channel=118
    32, 27, 31, 8, -25, -30, -8, -13, 2,
    -- layer=1 filter=172 channel=119
    15, -8, -18, -32, -37, -76, -68, -39, -33,
    -- layer=1 filter=172 channel=120
    -29, -9, -36, 0, -7, -12, 26, 7, 25,
    -- layer=1 filter=172 channel=121
    24, 25, 8, -8, -10, -14, 7, -24, 5,
    -- layer=1 filter=172 channel=122
    -7, -2, 5, 10, -7, -5, -3, -2, -7,
    -- layer=1 filter=172 channel=123
    7, 9, 14, -29, -4, 0, -21, -29, -13,
    -- layer=1 filter=172 channel=124
    6, -2, 4, 2, 11, 2, 0, -8, -2,
    -- layer=1 filter=172 channel=125
    -99, -83, -98, -48, -28, -22, 78, 74, 56,
    -- layer=1 filter=172 channel=126
    -13, -8, 0, 47, 34, 15, 24, 39, 34,
    -- layer=1 filter=172 channel=127
    44, 24, 33, 27, -24, -30, -10, -12, 12,
    -- layer=1 filter=173 channel=0
    9, -3, 10, 14, 4, -2, 9, 2, 9,
    -- layer=1 filter=173 channel=1
    -28, -51, -38, -13, -33, -20, -27, -5, -21,
    -- layer=1 filter=173 channel=2
    -11, -8, 4, -16, -4, 0, 0, 0, -9,
    -- layer=1 filter=173 channel=3
    0, -10, 10, -2, -9, -10, -3, 7, 4,
    -- layer=1 filter=173 channel=4
    8, 11, -7, 8, 0, -4, -6, 10, 3,
    -- layer=1 filter=173 channel=5
    -47, -65, -57, -54, -41, -31, -60, -26, -50,
    -- layer=1 filter=173 channel=6
    32, 24, 20, 11, 14, 11, 35, -4, -20,
    -- layer=1 filter=173 channel=7
    -84, -123, -82, -23, -157, -122, 25, -33, -71,
    -- layer=1 filter=173 channel=8
    -65, -99, -47, -91, -99, -75, -80, -85, -68,
    -- layer=1 filter=173 channel=9
    -4, -21, -8, -26, -14, -9, -14, -4, 13,
    -- layer=1 filter=173 channel=10
    -56, -95, -73, -9, -117, -75, 54, -20, -56,
    -- layer=1 filter=173 channel=11
    8, 19, 1, 13, 18, 5, 26, 18, 18,
    -- layer=1 filter=173 channel=12
    -14, -32, 0, -30, -25, -32, 48, 39, 17,
    -- layer=1 filter=173 channel=13
    13, -1, -6, 21, 7, -12, 9, 4, -16,
    -- layer=1 filter=173 channel=14
    -49, -49, 0, -15, -93, -42, 31, -5, -79,
    -- layer=1 filter=173 channel=15
    17, -17, -13, 11, -53, -21, 18, -68, -30,
    -- layer=1 filter=173 channel=16
    -83, -74, -60, -92, -111, -90, -79, -90, -89,
    -- layer=1 filter=173 channel=17
    18, 13, 1, 24, 17, 20, 1, 20, 9,
    -- layer=1 filter=173 channel=18
    -23, -24, -23, 1, -27, -20, 42, 29, 0,
    -- layer=1 filter=173 channel=19
    7, -27, -7, -42, -126, -89, -59, -91, -100,
    -- layer=1 filter=173 channel=20
    27, 19, 16, 9, 12, 5, 7, 0, 15,
    -- layer=1 filter=173 channel=21
    -23, -12, -22, -16, -12, -1, -2, -21, -15,
    -- layer=1 filter=173 channel=22
    9, 0, 0, 1, 8, 2, 3, -1, 0,
    -- layer=1 filter=173 channel=23
    11, -31, -1, -5, -23, -21, -4, -4, -26,
    -- layer=1 filter=173 channel=24
    -13, -22, -15, 5, -17, -15, 0, -12, -20,
    -- layer=1 filter=173 channel=25
    -80, -70, -57, -51, -122, -84, -6, -58, -108,
    -- layer=1 filter=173 channel=26
    12, -27, -8, 6, -22, -40, 14, -20, -29,
    -- layer=1 filter=173 channel=27
    16, 21, -4, 20, 29, 16, 29, 44, 26,
    -- layer=1 filter=173 channel=28
    -32, -30, -20, 2, -68, -25, 25, -17, -44,
    -- layer=1 filter=173 channel=29
    -1, 6, 1, 2, 6, 1, -13, -3, 10,
    -- layer=1 filter=173 channel=30
    -28, -77, -54, -30, -104, -71, -3, -30, -66,
    -- layer=1 filter=173 channel=31
    -25, -50, -54, -35, -27, -52, 25, 6, -36,
    -- layer=1 filter=173 channel=32
    20, -79, -49, 23, -65, -64, 30, -43, -26,
    -- layer=1 filter=173 channel=33
    4, -5, -11, -8, 8, 0, 9, 2, 8,
    -- layer=1 filter=173 channel=34
    12, 4, 10, 2, -2, 2, 13, 6, -7,
    -- layer=1 filter=173 channel=35
    -4, -8, -15, -10, -4, -8, -10, -16, -4,
    -- layer=1 filter=173 channel=36
    32, 33, 13, 18, 34, 32, 25, 31, 34,
    -- layer=1 filter=173 channel=37
    -73, -53, -68, -85, -46, -52, -55, -74, -74,
    -- layer=1 filter=173 channel=38
    23, 8, 17, 8, 6, 9, 18, 9, -12,
    -- layer=1 filter=173 channel=39
    -1, 2, -3, -7, -9, -4, 2, 15, -3,
    -- layer=1 filter=173 channel=40
    -64, -52, -31, -16, -44, -29, 48, 10, -39,
    -- layer=1 filter=173 channel=41
    23, -9, -8, 10, -9, -31, 1, -45, -15,
    -- layer=1 filter=173 channel=42
    -22, -19, 4, -9, -3, 5, 33, -9, -36,
    -- layer=1 filter=173 channel=43
    -53, -64, -55, -97, -107, -64, -78, -90, -72,
    -- layer=1 filter=173 channel=44
    4, -94, -53, -3, -87, -72, 26, -46, -26,
    -- layer=1 filter=173 channel=45
    20, -2, 4, 8, 4, -4, 23, 8, -15,
    -- layer=1 filter=173 channel=46
    -12, -7, 30, -86, -98, -78, -64, -90, -101,
    -- layer=1 filter=173 channel=47
    9, -22, -25, 28, -20, -19, 12, -11, -55,
    -- layer=1 filter=173 channel=48
    8, -8, 0, 14, 3, 4, 10, -6, -7,
    -- layer=1 filter=173 channel=49
    -6, -2, 1, -22, -5, -9, -9, -19, -30,
    -- layer=1 filter=173 channel=50
    1, -2, 4, 2, 2, 0, -4, 3, 4,
    -- layer=1 filter=173 channel=51
    -5, 8, 17, 2, -19, -2, 35, -4, -24,
    -- layer=1 filter=173 channel=52
    0, 6, 6, -2, 0, -2, 7, -11, -4,
    -- layer=1 filter=173 channel=53
    -19, -8, -14, -12, -1, -14, -15, -4, -8,
    -- layer=1 filter=173 channel=54
    -50, -34, -24, -42, -67, -54, -8, -41, -72,
    -- layer=1 filter=173 channel=55
    23, 27, 16, 28, 26, 33, 23, 43, 24,
    -- layer=1 filter=173 channel=56
    -6, -1, -1, 8, -3, -2, 7, 3, -4,
    -- layer=1 filter=173 channel=57
    -76, -77, -64, -20, -104, -59, 63, 6, -52,
    -- layer=1 filter=173 channel=58
    -41, -92, -49, -24, -90, -73, 17, 4, -80,
    -- layer=1 filter=173 channel=59
    2, -6, -15, -14, -7, 4, -5, -13, 5,
    -- layer=1 filter=173 channel=60
    -7, -18, -6, -2, -3, -6, -12, -8, -14,
    -- layer=1 filter=173 channel=61
    -9, 0, -9, 3, 2, 7, 0, 7, -7,
    -- layer=1 filter=173 channel=62
    -110, -110, -73, -147, -137, -111, -104, -114, -105,
    -- layer=1 filter=173 channel=63
    7, 11, 5, 11, 27, 6, 27, 27, 16,
    -- layer=1 filter=173 channel=64
    6, 7, -5, -9, -10, -6, -9, 1, 12,
    -- layer=1 filter=173 channel=65
    -10, 9, 0, 2, -15, -7, 1, -6, -3,
    -- layer=1 filter=173 channel=66
    8, 19, 7, 8, 12, 12, 0, 19, 6,
    -- layer=1 filter=173 channel=67
    6, -21, -29, -22, -18, -17, -14, -52, -30,
    -- layer=1 filter=173 channel=68
    -14, -108, -76, -11, -103, -91, 16, -58, -36,
    -- layer=1 filter=173 channel=69
    -5, -32, -29, -6, -39, -42, -12, -23, -63,
    -- layer=1 filter=173 channel=70
    20, 1, -11, -15, -13, -39, 28, -16, -34,
    -- layer=1 filter=173 channel=71
    -12, -12, 0, -24, -11, -5, -20, -12, -6,
    -- layer=1 filter=173 channel=72
    34, 7, 37, -22, -68, -37, 0, -20, -17,
    -- layer=1 filter=173 channel=73
    6, 3, 10, 13, 11, 2, 4, -2, 9,
    -- layer=1 filter=173 channel=74
    8, -43, -26, -10, -53, -51, 9, -2, 3,
    -- layer=1 filter=173 channel=75
    -23, -49, -11, -56, -100, -59, 43, 7, 7,
    -- layer=1 filter=173 channel=76
    3, 7, -12, 0, 8, -11, 0, 3, -9,
    -- layer=1 filter=173 channel=77
    -15, -29, -10, -12, -20, -12, -2, -13, -20,
    -- layer=1 filter=173 channel=78
    -2, -3, 12, 21, 6, 6, 8, 14, 0,
    -- layer=1 filter=173 channel=79
    -43, -64, -57, -86, -87, -91, -60, -58, -66,
    -- layer=1 filter=173 channel=80
    7, 2, -4, -8, -5, -3, -7, -2, 0,
    -- layer=1 filter=173 channel=81
    -12, -16, -22, -6, -12, -13, 2, -8, 6,
    -- layer=1 filter=173 channel=82
    -19, -12, -6, -20, -24, -8, -11, -23, -23,
    -- layer=1 filter=173 channel=83
    2, -18, -22, 8, -13, -20, 0, -20, -33,
    -- layer=1 filter=173 channel=84
    -74, -87, -68, -37, -58, -62, 23, -18, -4,
    -- layer=1 filter=173 channel=85
    -2, -48, -5, -1, -19, -8, 13, 14, -33,
    -- layer=1 filter=173 channel=86
    10, 19, 25, 8, 27, 14, 12, 20, 13,
    -- layer=1 filter=173 channel=87
    27, -23, -6, -39, -38, -72, -6, -75, -49,
    -- layer=1 filter=173 channel=88
    -31, -25, -27, -30, -21, -23, -10, -19, -33,
    -- layer=1 filter=173 channel=89
    -12, -28, -17, -20, -12, -26, -8, -33, -25,
    -- layer=1 filter=173 channel=90
    -6, -105, -54, 0, -94, -86, 35, -76, -51,
    -- layer=1 filter=173 channel=91
    24, 19, 21, 23, 14, 8, 26, 3, 2,
    -- layer=1 filter=173 channel=92
    50, -27, 16, 46, -35, -34, 65, -49, -4,
    -- layer=1 filter=173 channel=93
    -3, 14, 6, -2, -2, 19, 7, 2, 11,
    -- layer=1 filter=173 channel=94
    11, 2, 12, 25, 14, 7, 17, 7, 18,
    -- layer=1 filter=173 channel=95
    -91, -76, -71, -52, -67, -67, -3, -32, -38,
    -- layer=1 filter=173 channel=96
    -4, 14, 7, 12, 16, 13, 1, 25, 13,
    -- layer=1 filter=173 channel=97
    22, 19, 18, 15, 5, 7, 1, 5, 19,
    -- layer=1 filter=173 channel=98
    -25, -44, -42, -51, -64, -45, -58, -41, -43,
    -- layer=1 filter=173 channel=99
    -44, -56, -65, -1, -57, -46, 49, -2, -49,
    -- layer=1 filter=173 channel=100
    20, 9, 0, 8, 8, 8, 10, 17, 3,
    -- layer=1 filter=173 channel=101
    7, 17, 7, 17, 18, 13, 6, 19, 16,
    -- layer=1 filter=173 channel=102
    15, 20, 14, 24, 5, 21, 19, 5, 20,
    -- layer=1 filter=173 channel=103
    0, 19, 12, -7, 10, 7, 17, 18, 6,
    -- layer=1 filter=173 channel=104
    -3, -18, 13, -16, 4, -3, -15, 18, -5,
    -- layer=1 filter=173 channel=105
    16, 19, 14, 21, 15, 21, 11, 23, 19,
    -- layer=1 filter=173 channel=106
    18, 8, 7, 35, 15, -6, 13, -9, 2,
    -- layer=1 filter=173 channel=107
    2, -4, 1, 2, 13, 7, -1, -9, -3,
    -- layer=1 filter=173 channel=108
    -27, -128, -63, -20, -124, -98, -1, -91, -53,
    -- layer=1 filter=173 channel=109
    7, 2, -5, -7, 0, -3, -5, 0, -5,
    -- layer=1 filter=173 channel=110
    4, 1, 3, -8, -5, 6, 2, 5, -1,
    -- layer=1 filter=173 channel=111
    -74, -63, -32, -8, -39, -36, 53, 23, -13,
    -- layer=1 filter=173 channel=112
    -31, -4, 0, -2, -27, -11, 59, 29, 22,
    -- layer=1 filter=173 channel=113
    -13, -34, -31, -25, -43, -39, -2, -52, -38,
    -- layer=1 filter=173 channel=114
    -28, -15, -37, 4, 9, 0, -15, 10, -16,
    -- layer=1 filter=173 channel=115
    8, 22, 17, 18, 10, 29, 16, 23, 25,
    -- layer=1 filter=173 channel=116
    -2, 1, 9, 4, 9, -9, -5, -1, 1,
    -- layer=1 filter=173 channel=117
    -119, -91, -59, -38, -78, -53, 63, 55, -10,
    -- layer=1 filter=173 channel=118
    -46, -57, -47, -10, -62, -49, 22, -15, -12,
    -- layer=1 filter=173 channel=119
    -25, -102, -61, -5, -96, -100, 7, -78, -56,
    -- layer=1 filter=173 channel=120
    -16, 1, 0, -9, -10, -3, 23, 1, -6,
    -- layer=1 filter=173 channel=121
    23, 14, 31, 10, 8, 13, 6, -10, -13,
    -- layer=1 filter=173 channel=122
    -3, 0, 1, 7, 7, 9, -5, -5, 6,
    -- layer=1 filter=173 channel=123
    7, 23, 23, 17, 20, 25, 33, 35, 9,
    -- layer=1 filter=173 channel=124
    -9, -3, -5, -17, -8, -8, -1, -12, -15,
    -- layer=1 filter=173 channel=125
    21, -11, -25, 7, -21, -27, 34, -32, -42,
    -- layer=1 filter=173 channel=126
    -50, -91, -74, -65, -95, -58, -64, -63, -54,
    -- layer=1 filter=173 channel=127
    -56, -81, -44, -27, -40, -60, 31, -14, -14,
    -- layer=1 filter=174 channel=0
    -7, -10, -1, -6, -7, -9, -1, -7, -10,
    -- layer=1 filter=174 channel=1
    -3, -10, 4, 4, 5, -1, 8, -9, 6,
    -- layer=1 filter=174 channel=2
    -4, -5, -1, -10, -10, 6, 8, -6, 3,
    -- layer=1 filter=174 channel=3
    8, 1, -6, -6, -3, -2, 9, -6, -2,
    -- layer=1 filter=174 channel=4
    -5, -9, -9, -3, 0, -5, -5, -5, 0,
    -- layer=1 filter=174 channel=5
    -6, -3, -6, -9, 7, -2, -2, 3, -1,
    -- layer=1 filter=174 channel=6
    0, -3, 8, -10, -5, 4, 5, 3, 1,
    -- layer=1 filter=174 channel=7
    -2, -1, -1, 0, -1, 6, 0, -7, -9,
    -- layer=1 filter=174 channel=8
    2, 3, -3, -9, -1, -10, -12, -11, 6,
    -- layer=1 filter=174 channel=9
    -2, 0, 0, 0, 3, 6, -7, 5, -1,
    -- layer=1 filter=174 channel=10
    -6, 4, 7, 2, -3, -3, 5, -8, -3,
    -- layer=1 filter=174 channel=11
    2, -2, -2, -7, 3, -1, -7, 1, -1,
    -- layer=1 filter=174 channel=12
    3, -2, 4, -5, 2, 2, 8, -8, 7,
    -- layer=1 filter=174 channel=13
    -6, -12, 2, -9, 3, -11, 8, -12, 1,
    -- layer=1 filter=174 channel=14
    9, -4, 1, -4, -3, 3, -9, 7, 8,
    -- layer=1 filter=174 channel=15
    -2, -2, -9, -1, -6, 0, -7, 8, 0,
    -- layer=1 filter=174 channel=16
    5, -2, -10, -9, 2, 1, -7, -10, 4,
    -- layer=1 filter=174 channel=17
    -11, 6, -1, 3, 5, 5, -3, 8, -1,
    -- layer=1 filter=174 channel=18
    -5, 8, -8, 5, -4, -7, 6, -5, 8,
    -- layer=1 filter=174 channel=19
    -2, 3, -10, -3, -6, 0, -2, 0, -8,
    -- layer=1 filter=174 channel=20
    -2, -4, -3, 4, 1, -1, -8, -12, 0,
    -- layer=1 filter=174 channel=21
    5, -3, 4, 2, -5, 0, -6, 2, 1,
    -- layer=1 filter=174 channel=22
    7, -10, 2, 7, -6, 4, 8, -10, 0,
    -- layer=1 filter=174 channel=23
    -10, 0, 4, 0, -5, -7, -8, -10, 5,
    -- layer=1 filter=174 channel=24
    -1, 5, -4, -8, -11, 6, 0, -11, 0,
    -- layer=1 filter=174 channel=25
    -3, -7, -7, 2, 8, 4, -3, 1, 1,
    -- layer=1 filter=174 channel=26
    4, -8, 6, -1, -11, -6, -2, 0, -8,
    -- layer=1 filter=174 channel=27
    -4, -6, 9, 3, -3, -6, 4, -1, 8,
    -- layer=1 filter=174 channel=28
    3, -10, -2, -8, -9, 1, 6, -3, 7,
    -- layer=1 filter=174 channel=29
    9, -8, 9, -3, 7, 8, 2, 8, -8,
    -- layer=1 filter=174 channel=30
    6, -3, 2, -1, 6, 10, 5, 2, 1,
    -- layer=1 filter=174 channel=31
    -7, 5, -1, -4, 7, 1, 7, -3, -3,
    -- layer=1 filter=174 channel=32
    -11, 5, -5, 5, -6, -1, 6, -6, -6,
    -- layer=1 filter=174 channel=33
    10, -2, -3, 1, 1, -6, -5, -7, -8,
    -- layer=1 filter=174 channel=34
    0, 3, 2, -4, -7, 1, -1, 0, 8,
    -- layer=1 filter=174 channel=35
    -3, 7, 5, -7, 7, 4, 4, 2, 9,
    -- layer=1 filter=174 channel=36
    5, -3, -9, -4, 0, -7, 7, -2, 0,
    -- layer=1 filter=174 channel=37
    -3, 6, -9, 4, -8, -4, -1, -10, 6,
    -- layer=1 filter=174 channel=38
    -6, 7, 8, -2, -4, 8, -12, 8, 0,
    -- layer=1 filter=174 channel=39
    0, 8, 8, -7, -8, -5, 2, -2, -7,
    -- layer=1 filter=174 channel=40
    0, 10, -7, -6, -12, 2, -1, -7, 1,
    -- layer=1 filter=174 channel=41
    -9, -7, 5, 0, -11, 4, 3, 6, -9,
    -- layer=1 filter=174 channel=42
    7, 6, 8, -4, -1, -2, -6, 8, 9,
    -- layer=1 filter=174 channel=43
    -5, 2, -9, -2, -7, 8, -4, 0, -2,
    -- layer=1 filter=174 channel=44
    -8, -3, -8, -3, 7, 4, -5, -1, 0,
    -- layer=1 filter=174 channel=45
    -14, -9, -2, -4, 5, 0, -11, 8, 0,
    -- layer=1 filter=174 channel=46
    4, 6, -1, 6, -8, 7, 10, -3, -6,
    -- layer=1 filter=174 channel=47
    -8, -6, -8, -2, 5, 9, 5, 2, 6,
    -- layer=1 filter=174 channel=48
    3, 3, -4, -8, 2, 6, -6, -2, 6,
    -- layer=1 filter=174 channel=49
    -4, -11, 0, -10, 6, -8, 2, 8, -10,
    -- layer=1 filter=174 channel=50
    0, 0, -2, 4, -5, -9, -10, -12, -4,
    -- layer=1 filter=174 channel=51
    1, -8, -9, -10, -7, 5, 8, 1, 4,
    -- layer=1 filter=174 channel=52
    -7, -6, -7, -6, 3, -1, 8, 1, 5,
    -- layer=1 filter=174 channel=53
    7, -3, -11, -10, 6, -5, 8, 7, 2,
    -- layer=1 filter=174 channel=54
    8, -1, 1, -8, -7, -8, 0, -1, -3,
    -- layer=1 filter=174 channel=55
    7, 2, -2, 2, 0, 3, 5, -5, 6,
    -- layer=1 filter=174 channel=56
    8, 0, 4, 6, -4, 2, -9, -1, -11,
    -- layer=1 filter=174 channel=57
    5, -9, 0, -5, -10, 1, -10, -6, 0,
    -- layer=1 filter=174 channel=58
    -10, -1, -10, -2, -11, 4, -1, 2, 3,
    -- layer=1 filter=174 channel=59
    -10, -3, -9, 7, -7, 0, 0, -8, 7,
    -- layer=1 filter=174 channel=60
    8, -10, -5, 7, -1, -2, -1, 0, 3,
    -- layer=1 filter=174 channel=61
    5, 0, 0, -9, -4, 0, 4, 6, 2,
    -- layer=1 filter=174 channel=62
    -10, -12, -3, -4, 8, -8, 0, -10, 4,
    -- layer=1 filter=174 channel=63
    -7, -8, 2, -7, 4, -2, -10, -5, 0,
    -- layer=1 filter=174 channel=64
    2, -5, 4, -2, -9, 0, 0, 1, -3,
    -- layer=1 filter=174 channel=65
    -10, 1, -1, -1, 8, -11, 0, -9, 1,
    -- layer=1 filter=174 channel=66
    -9, -11, -10, 4, 4, -8, 7, -8, -6,
    -- layer=1 filter=174 channel=67
    -11, -9, 8, 9, 9, -1, 9, -1, 1,
    -- layer=1 filter=174 channel=68
    -5, -9, -11, -2, 2, 3, -2, -9, -1,
    -- layer=1 filter=174 channel=69
    -3, -9, 10, 4, 5, 6, -9, 3, -8,
    -- layer=1 filter=174 channel=70
    2, -9, 2, 1, 0, -7, 0, 0, -2,
    -- layer=1 filter=174 channel=71
    -8, 3, -9, -2, 5, 3, 3, 2, -1,
    -- layer=1 filter=174 channel=72
    -2, 4, -11, 1, -9, 5, -3, -11, 5,
    -- layer=1 filter=174 channel=73
    5, -11, -3, -10, 2, -2, -7, 7, -1,
    -- layer=1 filter=174 channel=74
    2, -6, -2, 0, 6, 0, -7, 1, 0,
    -- layer=1 filter=174 channel=75
    3, -5, 8, -1, -7, 6, 8, 7, 5,
    -- layer=1 filter=174 channel=76
    6, 1, -2, 3, 1, 1, -7, -8, 0,
    -- layer=1 filter=174 channel=77
    6, -10, 7, 8, -11, 7, 2, 8, -11,
    -- layer=1 filter=174 channel=78
    -3, 4, -9, -9, -10, -12, 0, 0, -8,
    -- layer=1 filter=174 channel=79
    0, -8, 10, 1, 7, 9, 0, 4, 1,
    -- layer=1 filter=174 channel=80
    8, 3, 9, -8, -3, -10, 1, -10, -9,
    -- layer=1 filter=174 channel=81
    3, -1, -9, -3, 8, -10, 7, -7, 1,
    -- layer=1 filter=174 channel=82
    2, 6, 7, -4, -8, -4, 7, 6, -4,
    -- layer=1 filter=174 channel=83
    7, 0, -7, 4, -1, -3, -2, -4, 5,
    -- layer=1 filter=174 channel=84
    -9, -10, 2, -1, -1, 1, 5, -1, 2,
    -- layer=1 filter=174 channel=85
    -10, 9, -9, 7, -10, -10, -9, 0, -4,
    -- layer=1 filter=174 channel=86
    3, -5, -11, 3, -6, 5, 1, 0, -5,
    -- layer=1 filter=174 channel=87
    -4, 0, -11, 7, 6, -11, -3, 8, -7,
    -- layer=1 filter=174 channel=88
    0, -7, -6, -8, -1, 5, 5, -2, -7,
    -- layer=1 filter=174 channel=89
    -1, -11, -9, -7, 3, 0, 6, -2, -11,
    -- layer=1 filter=174 channel=90
    0, -6, -4, -5, 4, 7, -3, -8, 0,
    -- layer=1 filter=174 channel=91
    -7, 6, -1, -1, 3, -7, -8, -1, -1,
    -- layer=1 filter=174 channel=92
    8, -5, 2, -6, -7, -4, -7, -9, 3,
    -- layer=1 filter=174 channel=93
    2, -1, -8, 8, 8, -9, -10, -6, 1,
    -- layer=1 filter=174 channel=94
    -10, -3, -3, 5, 0, 6, 8, 1, -9,
    -- layer=1 filter=174 channel=95
    -7, 2, -3, -7, -11, -1, 0, 0, -5,
    -- layer=1 filter=174 channel=96
    -7, -2, 0, -7, -7, 7, 4, -1, -8,
    -- layer=1 filter=174 channel=97
    1, 6, 8, 5, 0, -5, -3, -2, 6,
    -- layer=1 filter=174 channel=98
    -4, 0, 10, -8, -10, -9, 3, -9, -2,
    -- layer=1 filter=174 channel=99
    0, 2, 0, 4, -7, 4, -8, 5, -2,
    -- layer=1 filter=174 channel=100
    0, 8, -5, 0, 4, 2, -7, 8, 1,
    -- layer=1 filter=174 channel=101
    -3, -1, -7, 4, -6, 1, 2, -10, -11,
    -- layer=1 filter=174 channel=102
    5, -5, 0, -7, -7, -2, 2, 2, -10,
    -- layer=1 filter=174 channel=103
    5, 3, 2, 7, 1, 4, -2, 7, -5,
    -- layer=1 filter=174 channel=104
    7, 1, 7, 1, 7, -11, -1, 2, -5,
    -- layer=1 filter=174 channel=105
    -10, -4, -1, -6, -7, 1, -7, -2, -10,
    -- layer=1 filter=174 channel=106
    4, -7, 0, 7, 3, -8, 0, 4, -8,
    -- layer=1 filter=174 channel=107
    -9, 7, -9, -10, -10, 4, -4, -8, 7,
    -- layer=1 filter=174 channel=108
    5, -6, -2, -4, -10, 2, 6, 5, 9,
    -- layer=1 filter=174 channel=109
    -5, 2, 9, 0, 1, 2, -7, -8, -10,
    -- layer=1 filter=174 channel=110
    8, 5, -8, 6, -2, -3, 2, 4, 9,
    -- layer=1 filter=174 channel=111
    -9, 8, -5, 6, 10, 7, 0, 4, -8,
    -- layer=1 filter=174 channel=112
    0, 0, 6, -5, -4, -2, 1, 3, 8,
    -- layer=1 filter=174 channel=113
    1, 8, -10, 8, 6, -7, 6, 0, -9,
    -- layer=1 filter=174 channel=114
    -1, 5, 1, 6, 8, -6, 7, -5, -2,
    -- layer=1 filter=174 channel=115
    0, 4, 0, -11, -10, -7, -12, -2, -9,
    -- layer=1 filter=174 channel=116
    -7, -4, 2, -9, -5, -1, 3, -5, -5,
    -- layer=1 filter=174 channel=117
    -2, -5, -7, -8, -6, -9, 5, -5, 1,
    -- layer=1 filter=174 channel=118
    6, -7, 8, 3, 1, -10, -7, 2, -9,
    -- layer=1 filter=174 channel=119
    5, 6, 8, -10, -2, -5, 0, 2, 0,
    -- layer=1 filter=174 channel=120
    1, -2, -6, 0, 0, -5, 6, -4, 7,
    -- layer=1 filter=174 channel=121
    2, -1, -9, -8, -13, 0, 3, 8, 7,
    -- layer=1 filter=174 channel=122
    -1, 3, -8, -8, -8, 5, -8, 2, 2,
    -- layer=1 filter=174 channel=123
    -9, -7, 8, -9, 5, -12, -5, -3, 7,
    -- layer=1 filter=174 channel=124
    4, 9, 4, 4, 6, 1, -10, -11, 4,
    -- layer=1 filter=174 channel=125
    1, 1, 9, -9, -4, 6, 3, 7, 4,
    -- layer=1 filter=174 channel=126
    0, -7, -3, -10, 7, -3, -2, -7, -8,
    -- layer=1 filter=174 channel=127
    -6, 3, 0, 7, -7, -2, 0, -6, -4,
    -- layer=1 filter=175 channel=0
    -4, 1, -7, -10, 0, -6, -5, 4, -9,
    -- layer=1 filter=175 channel=1
    -1, -5, 2, 0, -6, 5, 0, 4, 5,
    -- layer=1 filter=175 channel=2
    2, -1, -7, -4, 3, 2, 6, -6, 2,
    -- layer=1 filter=175 channel=3
    0, -10, -2, 6, 4, -5, -7, 9, -4,
    -- layer=1 filter=175 channel=4
    3, -12, 7, 7, -4, -3, 2, -1, -3,
    -- layer=1 filter=175 channel=5
    3, 0, -7, -2, -7, 4, -5, 2, -5,
    -- layer=1 filter=175 channel=6
    4, -1, 8, -9, -4, -9, -9, 7, -7,
    -- layer=1 filter=175 channel=7
    0, -3, -2, -2, 1, -10, -4, 0, -3,
    -- layer=1 filter=175 channel=8
    0, 0, -6, -10, -6, 2, 3, -9, 5,
    -- layer=1 filter=175 channel=9
    0, 4, -6, -10, -2, 6, 4, 2, -2,
    -- layer=1 filter=175 channel=10
    -5, -7, 8, -2, 7, -5, -3, -10, -3,
    -- layer=1 filter=175 channel=11
    -6, 0, -12, 6, -10, -5, -11, -7, -1,
    -- layer=1 filter=175 channel=12
    2, -4, -8, -3, -5, 2, -2, 2, -6,
    -- layer=1 filter=175 channel=13
    -8, -9, 0, -6, -12, -10, 1, -3, 4,
    -- layer=1 filter=175 channel=14
    4, -5, 4, 0, 0, 1, 6, 0, 0,
    -- layer=1 filter=175 channel=15
    6, -6, 0, 4, 1, -3, 5, -3, -2,
    -- layer=1 filter=175 channel=16
    -1, -10, 1, -3, 5, -3, 1, 7, 5,
    -- layer=1 filter=175 channel=17
    7, 5, -3, -11, 9, 6, -5, 7, 8,
    -- layer=1 filter=175 channel=18
    -2, -9, -11, -7, 7, 0, -9, -10, 6,
    -- layer=1 filter=175 channel=19
    7, -11, 4, -10, 1, 4, -6, -7, -9,
    -- layer=1 filter=175 channel=20
    5, -9, -8, 0, 2, 6, -13, -3, 2,
    -- layer=1 filter=175 channel=21
    6, 3, 6, -4, 8, -9, -4, -8, -1,
    -- layer=1 filter=175 channel=22
    -4, 5, 8, 7, -3, 8, -7, 3, -1,
    -- layer=1 filter=175 channel=23
    -1, 3, -2, 7, 9, 10, -9, 10, -9,
    -- layer=1 filter=175 channel=24
    1, 6, -6, -3, -6, -3, 8, -3, 3,
    -- layer=1 filter=175 channel=25
    2, 0, 3, 5, -10, -5, 0, -5, -3,
    -- layer=1 filter=175 channel=26
    -13, 0, 7, -12, 4, -1, -10, 2, 4,
    -- layer=1 filter=175 channel=27
    -5, -8, -1, -6, 6, -8, 4, 5, -2,
    -- layer=1 filter=175 channel=28
    -3, -5, -5, -9, -3, -6, -7, 1, 5,
    -- layer=1 filter=175 channel=29
    -4, -9, 7, 5, -11, -4, 4, -1, -9,
    -- layer=1 filter=175 channel=30
    -9, -9, 4, -12, 0, 8, 4, 2, -12,
    -- layer=1 filter=175 channel=31
    9, 2, 0, -8, 0, -9, 3, 7, -10,
    -- layer=1 filter=175 channel=32
    -12, 5, -5, -14, 1, 0, -7, -8, -12,
    -- layer=1 filter=175 channel=33
    0, 2, 5, 1, -8, 5, 9, 5, 2,
    -- layer=1 filter=175 channel=34
    8, 1, -3, 6, 1, 3, 0, -6, 6,
    -- layer=1 filter=175 channel=35
    -2, -5, -7, 2, -9, -9, -9, 4, -5,
    -- layer=1 filter=175 channel=36
    -9, -2, -10, 6, -11, 8, 3, 0, -7,
    -- layer=1 filter=175 channel=37
    -4, -12, -1, 5, 0, 0, 2, 3, -6,
    -- layer=1 filter=175 channel=38
    4, -6, 8, -1, -8, 0, -10, -4, 0,
    -- layer=1 filter=175 channel=39
    0, -7, 1, -8, -3, -6, 6, -2, -9,
    -- layer=1 filter=175 channel=40
    -7, -1, 10, -6, -10, -6, 0, -11, 5,
    -- layer=1 filter=175 channel=41
    6, -6, 1, -3, 6, 0, -4, -8, -10,
    -- layer=1 filter=175 channel=42
    5, 0, -1, 1, 4, 2, -5, -2, 2,
    -- layer=1 filter=175 channel=43
    4, -7, -11, -6, 3, -1, 3, 10, -3,
    -- layer=1 filter=175 channel=44
    3, -12, 3, 7, 4, -7, -2, -4, 0,
    -- layer=1 filter=175 channel=45
    5, -11, -12, -5, 6, -8, -1, 0, -6,
    -- layer=1 filter=175 channel=46
    -2, -7, 2, -10, -7, 3, 5, 7, -8,
    -- layer=1 filter=175 channel=47
    0, 2, -11, -2, -7, 7, 3, -12, -5,
    -- layer=1 filter=175 channel=48
    -8, 2, -6, -1, 4, -1, 6, -5, 3,
    -- layer=1 filter=175 channel=49
    7, -5, -11, -11, -3, 7, 1, 3, 4,
    -- layer=1 filter=175 channel=50
    -6, -12, -5, 1, -4, -3, -4, -3, -4,
    -- layer=1 filter=175 channel=51
    5, 5, 8, -7, -4, -4, 3, 6, 4,
    -- layer=1 filter=175 channel=52
    8, 6, 0, 5, -8, 1, 2, -8, 3,
    -- layer=1 filter=175 channel=53
    5, 4, -11, -8, -2, -10, -3, 4, 5,
    -- layer=1 filter=175 channel=54
    -11, 8, 4, -11, 4, 6, -10, 0, 0,
    -- layer=1 filter=175 channel=55
    -3, -7, -7, 2, 5, -9, 0, -14, 0,
    -- layer=1 filter=175 channel=56
    4, 2, -6, 3, -6, 6, -4, 2, 0,
    -- layer=1 filter=175 channel=57
    0, 0, -5, -4, 3, -4, -9, -4, -6,
    -- layer=1 filter=175 channel=58
    3, 6, 0, 1, 1, 7, -12, -10, -3,
    -- layer=1 filter=175 channel=59
    -10, 0, 6, -3, -10, -4, 7, 3, 8,
    -- layer=1 filter=175 channel=60
    -6, -2, -7, 3, -10, 4, 0, 5, 7,
    -- layer=1 filter=175 channel=61
    -5, -9, 0, 0, -5, 0, 1, 8, -6,
    -- layer=1 filter=175 channel=62
    -10, 2, 1, 7, -11, -8, -9, -11, 3,
    -- layer=1 filter=175 channel=63
    -6, 0, -11, -11, 2, -1, 3, -6, 2,
    -- layer=1 filter=175 channel=64
    6, 2, -2, 0, 8, 0, 5, 6, -11,
    -- layer=1 filter=175 channel=65
    -7, 4, 3, -7, 3, 2, 4, 3, 0,
    -- layer=1 filter=175 channel=66
    -11, 8, -12, -6, -3, -1, -4, -8, 5,
    -- layer=1 filter=175 channel=67
    -1, 8, 6, 0, 2, 7, -1, -9, -2,
    -- layer=1 filter=175 channel=68
    -7, 3, 0, -4, 7, 1, -3, -5, 5,
    -- layer=1 filter=175 channel=69
    -5, 1, 7, -7, -1, 6, -6, -6, 3,
    -- layer=1 filter=175 channel=70
    2, 1, 0, -2, 4, 6, 1, -8, 5,
    -- layer=1 filter=175 channel=71
    -12, -7, 0, 1, 4, -1, -7, 0, 6,
    -- layer=1 filter=175 channel=72
    -1, -8, 6, -6, -7, -5, 7, 3, -6,
    -- layer=1 filter=175 channel=73
    1, -1, 2, -6, -1, -1, 1, 0, -3,
    -- layer=1 filter=175 channel=74
    -8, 6, -5, 5, 0, -10, 0, 2, -1,
    -- layer=1 filter=175 channel=75
    6, -8, -4, -1, 11, -5, 4, -1, 3,
    -- layer=1 filter=175 channel=76
    0, 0, -9, -1, 4, -7, 3, -2, 3,
    -- layer=1 filter=175 channel=77
    -8, -10, -1, 5, -1, 7, 7, 5, -8,
    -- layer=1 filter=175 channel=78
    -12, -5, -9, -8, -4, 0, 0, 6, -9,
    -- layer=1 filter=175 channel=79
    2, -8, -11, 7, 2, 4, -3, -7, -9,
    -- layer=1 filter=175 channel=80
    -5, 4, 2, 0, -2, -3, 2, 0, -7,
    -- layer=1 filter=175 channel=81
    3, -11, -8, -5, -3, 0, 0, 8, 1,
    -- layer=1 filter=175 channel=82
    0, -8, 8, 0, 8, 5, -2, -2, 0,
    -- layer=1 filter=175 channel=83
    4, -5, 0, 6, 3, -7, 7, -5, -9,
    -- layer=1 filter=175 channel=84
    -2, -7, 2, 0, -4, -1, 4, -3, -11,
    -- layer=1 filter=175 channel=85
    -12, -10, -4, 0, -4, -1, -7, -1, 5,
    -- layer=1 filter=175 channel=86
    4, -9, -8, -3, 6, 7, 1, -5, -9,
    -- layer=1 filter=175 channel=87
    6, 2, 1, -11, -3, 5, -10, -7, -4,
    -- layer=1 filter=175 channel=88
    8, -7, 5, 0, 2, -7, -8, -2, -7,
    -- layer=1 filter=175 channel=89
    1, 6, -5, -2, -5, -11, -1, 0, 9,
    -- layer=1 filter=175 channel=90
    -9, -8, -1, -10, 5, 3, 9, -3, 2,
    -- layer=1 filter=175 channel=91
    -3, -10, -9, 6, -8, 0, 7, -11, -4,
    -- layer=1 filter=175 channel=92
    -10, 4, 1, 1, -3, 3, 6, 0, -5,
    -- layer=1 filter=175 channel=93
    0, -7, 6, -1, -8, 5, -1, -6, -5,
    -- layer=1 filter=175 channel=94
    4, -9, 2, -11, -6, -12, 6, 5, 7,
    -- layer=1 filter=175 channel=95
    -9, -4, -5, 7, 2, -7, 4, 7, 5,
    -- layer=1 filter=175 channel=96
    1, 5, -2, 3, -9, -4, 7, 0, -3,
    -- layer=1 filter=175 channel=97
    -9, -7, 7, 3, -6, 0, 1, -5, -7,
    -- layer=1 filter=175 channel=98
    0, 0, 0, -11, -2, -3, -7, 2, 0,
    -- layer=1 filter=175 channel=99
    -5, 3, -8, 0, 1, -8, -6, -3, 8,
    -- layer=1 filter=175 channel=100
    8, 2, -10, 6, 1, 5, 6, 1, 1,
    -- layer=1 filter=175 channel=101
    -4, 5, -7, -1, -12, 6, -7, 4, -3,
    -- layer=1 filter=175 channel=102
    -12, 2, 3, -3, 7, 1, -12, -10, -2,
    -- layer=1 filter=175 channel=103
    -6, -10, 2, 8, 8, -11, 2, 7, 2,
    -- layer=1 filter=175 channel=104
    1, -8, 4, 3, -4, 3, 0, -4, -7,
    -- layer=1 filter=175 channel=105
    -10, -7, 5, -10, 9, -10, 1, 8, 2,
    -- layer=1 filter=175 channel=106
    5, -11, -12, 0, -3, -12, -12, 1, -1,
    -- layer=1 filter=175 channel=107
    -2, -3, -6, 5, -4, 0, -6, -8, 4,
    -- layer=1 filter=175 channel=108
    -4, 0, 0, 0, -3, 9, 1, -3, -1,
    -- layer=1 filter=175 channel=109
    -10, 6, 3, -5, -7, 0, -7, 6, 6,
    -- layer=1 filter=175 channel=110
    2, -6, -12, 3, 2, -10, 2, -2, -11,
    -- layer=1 filter=175 channel=111
    -7, 3, 0, -6, -4, 7, 3, 0, 0,
    -- layer=1 filter=175 channel=112
    5, -3, -10, -7, 0, -8, -5, -5, -5,
    -- layer=1 filter=175 channel=113
    7, 1, 7, -2, -2, -6, -7, -6, -7,
    -- layer=1 filter=175 channel=114
    -7, 0, -7, 5, -9, 4, 5, -2, 2,
    -- layer=1 filter=175 channel=115
    5, -4, -1, 3, -4, -12, -8, 2, 6,
    -- layer=1 filter=175 channel=116
    3, -7, 0, 0, -3, -1, -5, 9, 2,
    -- layer=1 filter=175 channel=117
    3, -5, -7, -4, 5, 5, 1, 1, -2,
    -- layer=1 filter=175 channel=118
    1, -9, 1, 0, -8, -5, 0, 7, -4,
    -- layer=1 filter=175 channel=119
    2, -4, -7, -6, 7, -4, 5, 7, 1,
    -- layer=1 filter=175 channel=120
    6, -11, -6, -4, -5, -5, -7, 0, -3,
    -- layer=1 filter=175 channel=121
    0, -3, -9, 5, 1, 2, -7, 2, 0,
    -- layer=1 filter=175 channel=122
    0, -4, 7, -7, -4, 5, -8, -3, -3,
    -- layer=1 filter=175 channel=123
    -4, -6, 3, 6, 4, 4, 4, -7, 3,
    -- layer=1 filter=175 channel=124
    2, -11, -9, -9, -9, 1, 5, -2, -11,
    -- layer=1 filter=175 channel=125
    -5, -4, 0, -7, -5, 8, -10, 4, -6,
    -- layer=1 filter=175 channel=126
    -3, -3, -4, -2, 0, -2, -7, 2, 5,
    -- layer=1 filter=175 channel=127
    -13, -7, -4, -2, -4, 5, 7, 2, -2,
    -- layer=1 filter=176 channel=0
    -14, -11, -8, -31, -16, -14, -11, -31, 1,
    -- layer=1 filter=176 channel=1
    0, 3, -26, -10, 0, -14, 5, 7, -3,
    -- layer=1 filter=176 channel=2
    -20, -22, 9, -23, 0, -20, 15, -2, -6,
    -- layer=1 filter=176 channel=3
    -7, -8, -9, 2, 3, -5, -8, -12, -1,
    -- layer=1 filter=176 channel=4
    -7, 1, 6, -2, -11, 0, 2, -11, -9,
    -- layer=1 filter=176 channel=5
    18, -3, 3, 3, -4, -23, 0, -9, -4,
    -- layer=1 filter=176 channel=6
    3, 17, 13, 7, 14, 9, 1, 20, -8,
    -- layer=1 filter=176 channel=7
    37, 36, 8, 40, 69, 26, 25, 37, 35,
    -- layer=1 filter=176 channel=8
    26, -4, -5, 1, -4, -8, 7, -3, 5,
    -- layer=1 filter=176 channel=9
    -4, -22, -13, 24, 8, -1, -25, 8, -2,
    -- layer=1 filter=176 channel=10
    30, 23, 0, 24, 55, 1, 17, 30, 24,
    -- layer=1 filter=176 channel=11
    -6, -7, -22, 6, 2, -2, 6, -8, 1,
    -- layer=1 filter=176 channel=12
    -40, -56, -19, -46, -37, -16, 16, -5, 8,
    -- layer=1 filter=176 channel=13
    1, 13, 10, 2, 16, 5, -8, 9, 0,
    -- layer=1 filter=176 channel=14
    -7, -24, -2, 11, 24, 10, 32, 4, 12,
    -- layer=1 filter=176 channel=15
    8, 18, 6, 20, 7, 18, 41, 36, -5,
    -- layer=1 filter=176 channel=16
    15, -26, -9, 15, 5, -5, 17, -14, 1,
    -- layer=1 filter=176 channel=17
    7, -10, 14, -16, -2, -2, -10, 0, -15,
    -- layer=1 filter=176 channel=18
    -1, 9, -4, -6, -5, -24, -18, -5, 7,
    -- layer=1 filter=176 channel=19
    3, -13, -13, 28, 1, 7, -1, 18, 7,
    -- layer=1 filter=176 channel=20
    3, 14, 9, 7, 15, -3, 0, 15, 1,
    -- layer=1 filter=176 channel=21
    -12, -15, -13, -3, -2, 7, -3, -6, -1,
    -- layer=1 filter=176 channel=22
    18, 28, -1, 10, 18, 21, 4, 8, 3,
    -- layer=1 filter=176 channel=23
    -6, 37, -31, 32, 18, 10, 23, 35, -1,
    -- layer=1 filter=176 channel=24
    -22, -48, -2, -16, -19, -5, 7, -9, -14,
    -- layer=1 filter=176 channel=25
    12, 5, -20, 15, 46, 11, 22, 0, 24,
    -- layer=1 filter=176 channel=26
    -11, 14, 23, 15, 22, 12, 17, 27, -16,
    -- layer=1 filter=176 channel=27
    0, -23, -25, -34, -48, -42, -38, -68, -53,
    -- layer=1 filter=176 channel=28
    -7, -3, -14, -12, 5, -5, -16, -12, 10,
    -- layer=1 filter=176 channel=29
    -1, 4, 8, 8, -27, -17, 10, -5, 1,
    -- layer=1 filter=176 channel=30
    -9, -10, 19, 8, 4, -10, -22, -1, -3,
    -- layer=1 filter=176 channel=31
    6, 19, 22, 16, 7, -8, 11, 22, 2,
    -- layer=1 filter=176 channel=32
    6, 21, 14, 22, 41, 20, 25, 37, 1,
    -- layer=1 filter=176 channel=33
    7, 20, 6, 6, 12, -6, 12, 12, -13,
    -- layer=1 filter=176 channel=34
    -11, -6, -1, -19, 6, -22, 13, 17, 2,
    -- layer=1 filter=176 channel=35
    7, 5, 8, -1, 18, 18, -4, -6, 11,
    -- layer=1 filter=176 channel=36
    -7, -39, -31, -10, -23, -14, -5, -36, -29,
    -- layer=1 filter=176 channel=37
    5, -14, -15, 5, -10, 0, -4, 5, -7,
    -- layer=1 filter=176 channel=38
    -3, 18, 18, -11, 20, 13, -8, 12, 1,
    -- layer=1 filter=176 channel=39
    -25, -7, -5, 0, -20, -20, -3, -9, -6,
    -- layer=1 filter=176 channel=40
    25, 32, 21, 6, 21, 1, 10, 24, 22,
    -- layer=1 filter=176 channel=41
    14, -7, -19, 21, 52, -28, 14, 29, -14,
    -- layer=1 filter=176 channel=42
    -20, -2, -17, -24, -22, -8, 20, -3, 7,
    -- layer=1 filter=176 channel=43
    5, -7, -19, -2, -2, -8, 17, 14, 3,
    -- layer=1 filter=176 channel=44
    -2, 20, 16, 7, 28, -4, 8, 8, -11,
    -- layer=1 filter=176 channel=45
    3, -14, 6, 16, 6, -1, 19, 3, 1,
    -- layer=1 filter=176 channel=46
    -29, -28, -20, 15, -3, -2, -3, 4, 13,
    -- layer=1 filter=176 channel=47
    0, 26, -11, 3, 19, -5, 0, 22, 5,
    -- layer=1 filter=176 channel=48
    -18, -7, 0, -16, 0, -4, -9, -16, 5,
    -- layer=1 filter=176 channel=49
    3, 0, -8, -2, 14, 2, -3, -4, -2,
    -- layer=1 filter=176 channel=50
    -14, -1, -10, -12, -15, -15, -6, -7, -29,
    -- layer=1 filter=176 channel=51
    11, -7, 0, -7, 18, 4, -11, -5, 16,
    -- layer=1 filter=176 channel=52
    5, -4, -3, -7, 17, 0, 15, 19, -3,
    -- layer=1 filter=176 channel=53
    8, -8, 0, 5, 7, -5, 6, 3, 5,
    -- layer=1 filter=176 channel=54
    9, 2, -10, 18, 24, 3, 16, 12, 34,
    -- layer=1 filter=176 channel=55
    0, 0, -12, 8, 4, -4, 16, -2, -14,
    -- layer=1 filter=176 channel=56
    0, -5, 7, 3, -1, 10, 8, 8, 13,
    -- layer=1 filter=176 channel=57
    31, 25, 21, 20, 44, 16, 8, 20, 18,
    -- layer=1 filter=176 channel=58
    30, 66, -5, 55, 82, 26, 39, 71, 41,
    -- layer=1 filter=176 channel=59
    7, 4, -4, -5, 5, -8, 0, 3, 6,
    -- layer=1 filter=176 channel=60
    15, 7, 17, 0, 18, 5, 10, 16, 10,
    -- layer=1 filter=176 channel=61
    8, -11, -7, 2, -18, -15, -8, 1, -14,
    -- layer=1 filter=176 channel=62
    11, -5, -9, 3, -3, 8, 13, 9, 6,
    -- layer=1 filter=176 channel=63
    -26, -25, -40, -16, -25, -40, -5, -38, -14,
    -- layer=1 filter=176 channel=64
    -6, 2, 4, 0, -9, 0, -10, -4, 2,
    -- layer=1 filter=176 channel=65
    -6, -13, 10, -7, 0, 9, -3, 2, 3,
    -- layer=1 filter=176 channel=66
    -16, -10, -16, -16, -19, -15, -16, -35, -22,
    -- layer=1 filter=176 channel=67
    -34, -41, -25, -38, -48, -45, -35, -41, -9,
    -- layer=1 filter=176 channel=68
    11, 19, 28, 25, 39, 15, 21, 21, 19,
    -- layer=1 filter=176 channel=69
    5, -4, 23, 4, -3, 21, 14, 25, 6,
    -- layer=1 filter=176 channel=70
    -27, -13, -3, -23, -1, -23, -21, -7, -21,
    -- layer=1 filter=176 channel=71
    -33, -39, -19, -31, -30, -28, -12, -12, 1,
    -- layer=1 filter=176 channel=72
    13, -12, 2, 24, 24, 17, -23, 8, -1,
    -- layer=1 filter=176 channel=73
    11, 4, 7, 8, 2, 13, 7, -6, 6,
    -- layer=1 filter=176 channel=74
    -4, -10, -17, 1, -6, 10, -16, -1, 14,
    -- layer=1 filter=176 channel=75
    -43, -13, -18, -10, 6, 1, -1, 1, -12,
    -- layer=1 filter=176 channel=76
    -26, -22, -23, -16, 0, -40, -14, -27, -15,
    -- layer=1 filter=176 channel=77
    -30, -36, -3, -28, -37, -8, -14, -15, 13,
    -- layer=1 filter=176 channel=78
    -5, -17, 5, -9, 7, -3, 0, -9, 13,
    -- layer=1 filter=176 channel=79
    13, 5, -12, 3, -8, 5, -1, 11, 8,
    -- layer=1 filter=176 channel=80
    -1, 5, 9, -1, -6, 16, -1, 9, 15,
    -- layer=1 filter=176 channel=81
    -29, -54, -37, -30, -58, -28, -18, -26, -8,
    -- layer=1 filter=176 channel=82
    -23, -13, -9, -23, -8, -11, -1, 2, -6,
    -- layer=1 filter=176 channel=83
    -10, 4, 0, -10, -11, -19, 12, 10, -22,
    -- layer=1 filter=176 channel=84
    6, 0, -10, 14, 15, -34, 13, 4, -12,
    -- layer=1 filter=176 channel=85
    3, 20, -11, 23, 21, -6, -2, 44, 8,
    -- layer=1 filter=176 channel=86
    15, 7, -8, 5, -3, 0, 10, 0, -3,
    -- layer=1 filter=176 channel=87
    24, -11, 2, 21, 25, 31, -2, 35, 17,
    -- layer=1 filter=176 channel=88
    15, -13, 6, -4, 0, -5, -4, 0, 6,
    -- layer=1 filter=176 channel=89
    -19, -18, -9, -21, -20, -4, -15, -4, 4,
    -- layer=1 filter=176 channel=90
    7, 15, 29, 0, 26, 14, 7, 19, 0,
    -- layer=1 filter=176 channel=91
    12, 23, 21, 6, 17, 17, 6, 10, 14,
    -- layer=1 filter=176 channel=92
    -23, 14, 11, -20, 25, -11, 15, -13, 5,
    -- layer=1 filter=176 channel=93
    -23, -30, -20, -23, -18, -18, -9, -5, -4,
    -- layer=1 filter=176 channel=94
    -4, 1, -13, -26, -21, -10, -18, -29, 0,
    -- layer=1 filter=176 channel=95
    -6, -13, -12, 2, -10, -27, 1, -17, -14,
    -- layer=1 filter=176 channel=96
    -5, -5, -12, 7, -9, 2, 0, 0, -16,
    -- layer=1 filter=176 channel=97
    -15, -22, -14, -17, -21, -9, -13, -16, -14,
    -- layer=1 filter=176 channel=98
    1, 4, 4, -6, 5, 0, 8, -5, 6,
    -- layer=1 filter=176 channel=99
    3, -10, 24, 16, -13, 8, 14, -2, 33,
    -- layer=1 filter=176 channel=100
    -3, -24, -27, -1, 5, -20, 12, -31, -32,
    -- layer=1 filter=176 channel=101
    -5, 4, 6, 0, 16, 8, -2, 9, 2,
    -- layer=1 filter=176 channel=102
    -6, -5, 0, -39, -13, -8, -28, -27, -14,
    -- layer=1 filter=176 channel=103
    -9, -27, -4, -3, -14, -15, 3, -4, -7,
    -- layer=1 filter=176 channel=104
    0, 21, -23, 24, 8, 0, 3, 25, -13,
    -- layer=1 filter=176 channel=105
    -1, -4, -5, -24, -27, -23, -13, -31, 2,
    -- layer=1 filter=176 channel=106
    1, 20, 15, -7, 22, 7, 1, 1, -10,
    -- layer=1 filter=176 channel=107
    -17, 2, -5, -14, -8, -23, -17, 5, -2,
    -- layer=1 filter=176 channel=108
    -10, -4, 5, 17, 26, -5, 22, 33, -13,
    -- layer=1 filter=176 channel=109
    -3, 5, 0, -9, -6, 1, 2, -5, 9,
    -- layer=1 filter=176 channel=110
    4, 11, 0, -7, 0, -11, -6, -3, -9,
    -- layer=1 filter=176 channel=111
    -15, 4, -3, -10, 5, -30, -18, -18, -1,
    -- layer=1 filter=176 channel=112
    0, -14, -33, -19, 2, -60, 14, -12, 4,
    -- layer=1 filter=176 channel=113
    -9, 15, -15, -23, 0, -15, 0, 15, -18,
    -- layer=1 filter=176 channel=114
    22, -16, 8, 16, -12, -10, 10, 3, -3,
    -- layer=1 filter=176 channel=115
    12, 27, 3, 24, 24, -8, 11, 0, 8,
    -- layer=1 filter=176 channel=116
    3, 9, 1, -4, 0, 7, -8, 9, -1,
    -- layer=1 filter=176 channel=117
    -20, -11, -21, 1, -20, -26, 0, -2, 16,
    -- layer=1 filter=176 channel=118
    -3, 1, 0, 5, -3, -9, -11, 12, 12,
    -- layer=1 filter=176 channel=119
    9, 4, 23, 19, 35, 7, 23, 33, -1,
    -- layer=1 filter=176 channel=120
    -2, -9, -22, -3, 7, 10, 1, -7, 8,
    -- layer=1 filter=176 channel=121
    -20, -11, 7, 5, 8, 2, -11, -12, -2,
    -- layer=1 filter=176 channel=122
    8, 3, -4, 8, 0, 2, -6, -2, 7,
    -- layer=1 filter=176 channel=123
    -23, -22, -11, -10, 0, -27, -7, 3, -16,
    -- layer=1 filter=176 channel=124
    16, 20, 12, 20, 11, 12, 7, 9, 4,
    -- layer=1 filter=176 channel=125
    -18, -23, 1, -2, 11, 3, -24, 8, 2,
    -- layer=1 filter=176 channel=126
    0, -10, -1, -29, -30, -5, -1, -13, -23,
    -- layer=1 filter=176 channel=127
    -1, 14, 14, 15, 6, -2, -1, 2, 12,
    -- layer=1 filter=177 channel=0
    5, -1, -3, 5, 0, -4, 6, 0, -2,
    -- layer=1 filter=177 channel=1
    -2, -6, -10, 6, -4, -11, -8, -12, 7,
    -- layer=1 filter=177 channel=2
    -1, 3, 10, 1, -2, -7, 2, -3, -8,
    -- layer=1 filter=177 channel=3
    1, 5, 5, 3, 0, 3, 0, 5, -9,
    -- layer=1 filter=177 channel=4
    -7, -5, 8, -9, -5, -8, -2, -5, -3,
    -- layer=1 filter=177 channel=5
    2, -8, -10, -6, 0, -2, -3, -6, -2,
    -- layer=1 filter=177 channel=6
    6, -9, 5, -10, -10, 0, -3, 7, 4,
    -- layer=1 filter=177 channel=7
    -8, -6, 0, 1, 0, 9, -11, -7, 0,
    -- layer=1 filter=177 channel=8
    -11, -6, -9, -3, -2, -6, -6, 0, -7,
    -- layer=1 filter=177 channel=9
    9, -5, 0, 4, -5, 7, -1, 1, -5,
    -- layer=1 filter=177 channel=10
    -6, 1, -3, -7, -1, 8, -8, 3, -6,
    -- layer=1 filter=177 channel=11
    0, -12, 4, 2, 5, 6, -5, -2, 7,
    -- layer=1 filter=177 channel=12
    -10, 5, -2, 6, -4, 0, -5, 6, 8,
    -- layer=1 filter=177 channel=13
    -4, -12, -3, -5, 2, -10, 0, -2, -9,
    -- layer=1 filter=177 channel=14
    3, -4, -1, 0, -9, -7, 8, 0, -7,
    -- layer=1 filter=177 channel=15
    8, -4, -5, -1, -7, -10, -5, -5, -2,
    -- layer=1 filter=177 channel=16
    0, -10, -7, -4, -4, 4, 6, 0, -12,
    -- layer=1 filter=177 channel=17
    -11, -3, -9, 0, -1, -11, 6, -6, -11,
    -- layer=1 filter=177 channel=18
    -2, 7, -3, -9, 0, -3, 1, 3, -12,
    -- layer=1 filter=177 channel=19
    -5, 2, 1, -5, 2, -3, 0, -3, -4,
    -- layer=1 filter=177 channel=20
    -3, 6, 4, -2, 7, -3, -2, -8, -3,
    -- layer=1 filter=177 channel=21
    -6, -3, -9, 0, 1, 0, 7, 0, 3,
    -- layer=1 filter=177 channel=22
    0, 6, -12, -12, -14, 0, -9, -5, -4,
    -- layer=1 filter=177 channel=23
    -2, -6, -3, -4, -5, -4, -1, -4, 6,
    -- layer=1 filter=177 channel=24
    -6, 0, 3, -1, 5, 6, -1, -8, 0,
    -- layer=1 filter=177 channel=25
    4, 3, 6, -2, -10, 0, -7, -7, 0,
    -- layer=1 filter=177 channel=26
    -6, -2, 6, -3, -8, -10, 3, 4, 8,
    -- layer=1 filter=177 channel=27
    6, 0, -4, -9, -8, 6, -5, 0, -8,
    -- layer=1 filter=177 channel=28
    0, 8, 1, 0, -6, -10, 9, 7, 3,
    -- layer=1 filter=177 channel=29
    0, 0, 9, 0, -5, -4, -3, -6, -4,
    -- layer=1 filter=177 channel=30
    -2, 4, 5, 5, 6, -6, 8, 1, -9,
    -- layer=1 filter=177 channel=31
    0, -9, 4, -7, -8, 7, -2, 0, -7,
    -- layer=1 filter=177 channel=32
    8, -2, -2, 2, -2, 4, -4, 2, 0,
    -- layer=1 filter=177 channel=33
    3, 7, 6, 0, 8, -7, -10, 3, -4,
    -- layer=1 filter=177 channel=34
    -2, -5, -9, -10, -10, 7, 7, -7, 1,
    -- layer=1 filter=177 channel=35
    -1, 0, -4, 8, -4, -12, -7, -4, -10,
    -- layer=1 filter=177 channel=36
    -8, -12, -13, -2, 5, -12, 4, -1, -1,
    -- layer=1 filter=177 channel=37
    2, -8, -6, -6, 4, 3, 1, -1, -2,
    -- layer=1 filter=177 channel=38
    6, -6, 0, 3, -2, 7, -9, 0, -9,
    -- layer=1 filter=177 channel=39
    2, -4, 0, -5, 4, 2, 5, -6, -11,
    -- layer=1 filter=177 channel=40
    4, 5, -6, -10, -6, 2, 0, 7, 3,
    -- layer=1 filter=177 channel=41
    -5, 9, 1, 2, 1, 5, 3, -3, 7,
    -- layer=1 filter=177 channel=42
    5, -8, -5, 2, -1, 0, -7, -1, 5,
    -- layer=1 filter=177 channel=43
    -3, -2, -3, 8, 6, -6, -10, -1, -2,
    -- layer=1 filter=177 channel=44
    -6, -7, 4, -1, -1, -4, -1, -5, 0,
    -- layer=1 filter=177 channel=45
    2, 0, 2, -3, 0, 5, 4, -6, 4,
    -- layer=1 filter=177 channel=46
    2, -2, -6, -7, -10, -9, -9, 10, -2,
    -- layer=1 filter=177 channel=47
    -5, 0, 8, 2, -6, -4, -5, -10, -2,
    -- layer=1 filter=177 channel=48
    -8, 8, -1, 6, -2, -5, 1, -12, 5,
    -- layer=1 filter=177 channel=49
    -3, -10, 5, 8, -10, 0, 2, 0, -6,
    -- layer=1 filter=177 channel=50
    -3, 1, -4, 3, -8, -9, 6, -9, 2,
    -- layer=1 filter=177 channel=51
    2, -7, 8, -6, -2, 0, 1, 9, -6,
    -- layer=1 filter=177 channel=52
    1, 5, 10, -13, 1, -2, -1, 8, -7,
    -- layer=1 filter=177 channel=53
    5, 1, -5, -10, 9, -4, -6, 6, 0,
    -- layer=1 filter=177 channel=54
    -7, 7, -10, 1, 0, 5, -3, -9, -2,
    -- layer=1 filter=177 channel=55
    -11, -11, -4, -9, -11, -12, -6, -6, -11,
    -- layer=1 filter=177 channel=56
    9, 4, -5, 3, 8, -5, -8, -8, 4,
    -- layer=1 filter=177 channel=57
    5, -1, 6, -11, -5, -4, 5, 0, 5,
    -- layer=1 filter=177 channel=58
    -6, 2, -7, 1, 3, -12, 8, 2, -6,
    -- layer=1 filter=177 channel=59
    6, -11, -4, -10, 5, 8, 2, 4, -9,
    -- layer=1 filter=177 channel=60
    -6, -5, 1, -6, -3, 1, -10, 4, -5,
    -- layer=1 filter=177 channel=61
    6, -9, 3, 8, 0, 4, 9, -1, 0,
    -- layer=1 filter=177 channel=62
    3, -5, 8, -7, 6, 7, 2, -13, -12,
    -- layer=1 filter=177 channel=63
    -7, 2, -4, 1, -5, -5, -1, -12, -10,
    -- layer=1 filter=177 channel=64
    8, 1, -5, 2, 2, -8, 4, -1, 2,
    -- layer=1 filter=177 channel=65
    6, 1, -4, -10, -3, -6, 8, 5, 4,
    -- layer=1 filter=177 channel=66
    5, -10, 4, -11, -2, -2, 1, 1, -6,
    -- layer=1 filter=177 channel=67
    7, 5, 7, 7, 12, 5, 4, -1, 7,
    -- layer=1 filter=177 channel=68
    2, 2, -9, 3, -10, -3, -1, -12, 0,
    -- layer=1 filter=177 channel=69
    4, -9, -3, -4, -7, 0, -3, 0, 5,
    -- layer=1 filter=177 channel=70
    5, 6, 3, -1, -4, 11, 3, 8, -5,
    -- layer=1 filter=177 channel=71
    -4, 2, -6, 0, 12, 5, 12, -6, -5,
    -- layer=1 filter=177 channel=72
    7, -11, -4, 1, 6, 3, -3, -2, -3,
    -- layer=1 filter=177 channel=73
    6, -11, 1, -6, 7, -8, -7, 4, -7,
    -- layer=1 filter=177 channel=74
    8, 6, 0, 6, 4, 3, 4, 8, -8,
    -- layer=1 filter=177 channel=75
    -6, 3, 5, -9, 7, -6, 9, 0, 5,
    -- layer=1 filter=177 channel=76
    1, 1, -7, -2, -1, 7, 3, -10, -7,
    -- layer=1 filter=177 channel=77
    0, 9, -1, -2, 4, -10, -7, -2, -9,
    -- layer=1 filter=177 channel=78
    -9, -10, 3, 0, -2, -7, -3, -1, 5,
    -- layer=1 filter=177 channel=79
    1, -6, -1, 4, 6, -12, 0, -1, 5,
    -- layer=1 filter=177 channel=80
    -6, -5, -4, -3, -3, 4, -8, -2, 8,
    -- layer=1 filter=177 channel=81
    -8, 8, 1, 1, -9, -1, 0, -7, -12,
    -- layer=1 filter=177 channel=82
    -1, -7, 5, 5, 7, 9, 10, -2, 1,
    -- layer=1 filter=177 channel=83
    3, 1, -8, -12, 5, 5, 3, 5, 4,
    -- layer=1 filter=177 channel=84
    -5, -1, -7, 4, -3, 7, -4, 7, -10,
    -- layer=1 filter=177 channel=85
    -9, -9, -10, -2, 0, -7, 0, -12, -1,
    -- layer=1 filter=177 channel=86
    5, 1, -13, 2, -13, 7, -5, -7, 0,
    -- layer=1 filter=177 channel=87
    0, -9, -6, -8, 4, -5, 5, 0, 3,
    -- layer=1 filter=177 channel=88
    3, -7, 6, 0, 4, -1, -7, 2, -9,
    -- layer=1 filter=177 channel=89
    -9, -3, -6, 0, -8, -5, 1, -1, 6,
    -- layer=1 filter=177 channel=90
    -10, -5, 8, 8, -7, 2, -4, -3, -3,
    -- layer=1 filter=177 channel=91
    3, -1, -11, -7, -10, -1, 7, 4, -4,
    -- layer=1 filter=177 channel=92
    -2, 2, 4, -4, -7, -6, 7, -2, -2,
    -- layer=1 filter=177 channel=93
    7, 2, 0, -6, 0, 0, -12, -4, 5,
    -- layer=1 filter=177 channel=94
    1, 7, 0, -10, -12, -7, 4, 1, 2,
    -- layer=1 filter=177 channel=95
    -4, 2, 0, -2, 8, -4, -10, 5, 2,
    -- layer=1 filter=177 channel=96
    4, 2, -9, 1, 3, 3, 0, 6, 0,
    -- layer=1 filter=177 channel=97
    -1, 0, -4, 8, 2, -2, 4, -3, -5,
    -- layer=1 filter=177 channel=98
    1, -10, -7, -3, -7, 7, 0, -1, -5,
    -- layer=1 filter=177 channel=99
    -1, -1, -9, 0, 7, 3, 1, 0, -3,
    -- layer=1 filter=177 channel=100
    5, 8, -5, -4, -1, -5, -12, 7, 7,
    -- layer=1 filter=177 channel=101
    8, 0, -7, 4, -7, 2, 5, -6, -2,
    -- layer=1 filter=177 channel=102
    -8, -6, 6, 3, -5, 0, -12, -9, 4,
    -- layer=1 filter=177 channel=103
    3, 1, -8, -13, 4, 2, -10, -2, 0,
    -- layer=1 filter=177 channel=104
    -11, 8, 0, -1, 0, -2, 1, 4, -9,
    -- layer=1 filter=177 channel=105
    -4, -4, -6, 8, 0, -2, -8, -11, -4,
    -- layer=1 filter=177 channel=106
    -1, -9, 6, 1, 1, -9, 0, -11, -5,
    -- layer=1 filter=177 channel=107
    3, 3, -8, -11, 6, 7, 0, 7, -7,
    -- layer=1 filter=177 channel=108
    7, 2, -5, -7, 8, 0, 8, 0, -8,
    -- layer=1 filter=177 channel=109
    -6, 2, -9, 3, 5, 6, -10, -6, -3,
    -- layer=1 filter=177 channel=110
    3, -11, -10, -4, 1, -8, -5, 8, 5,
    -- layer=1 filter=177 channel=111
    8, 8, -5, 6, 4, -10, 6, -1, 2,
    -- layer=1 filter=177 channel=112
    -11, 0, 3, 0, -4, -3, 0, 2, 0,
    -- layer=1 filter=177 channel=113
    -3, 0, 8, 1, -10, -2, 5, 9, 8,
    -- layer=1 filter=177 channel=114
    -3, 0, -4, 1, -2, 6, 5, 3, -7,
    -- layer=1 filter=177 channel=115
    -1, -8, 1, 5, -2, 2, -2, 4, -10,
    -- layer=1 filter=177 channel=116
    10, -4, -1, 8, -2, -1, 5, 1, 5,
    -- layer=1 filter=177 channel=117
    5, 8, -1, 6, 0, 0, 0, 0, 3,
    -- layer=1 filter=177 channel=118
    1, -3, -5, 6, 4, -3, -12, 3, -12,
    -- layer=1 filter=177 channel=119
    -4, -1, -8, -9, 5, 3, -4, 2, 0,
    -- layer=1 filter=177 channel=120
    -5, 2, 6, 0, 4, -11, -1, 6, 7,
    -- layer=1 filter=177 channel=121
    5, -3, -8, 1, 6, -7, -4, -4, -10,
    -- layer=1 filter=177 channel=122
    7, -7, 0, 4, 9, 2, -2, -2, -5,
    -- layer=1 filter=177 channel=123
    4, -2, -6, -7, -11, -5, -12, 3, -11,
    -- layer=1 filter=177 channel=124
    -4, -8, 4, 0, 3, -3, 7, 0, 3,
    -- layer=1 filter=177 channel=125
    -11, -13, -9, -2, 4, 4, 0, -11, -11,
    -- layer=1 filter=177 channel=126
    9, 0, -1, -5, -4, 2, -10, -1, 0,
    -- layer=1 filter=177 channel=127
    4, 0, -8, -3, 1, 6, -5, -14, -5,
    -- layer=1 filter=178 channel=0
    13, -20, -48, 14, -14, -46, 39, 1, -21,
    -- layer=1 filter=178 channel=1
    2, 6, -8, -10, 18, 10, -7, 36, 11,
    -- layer=1 filter=178 channel=2
    -19, 21, 61, -26, 0, 55, -29, -22, 30,
    -- layer=1 filter=178 channel=3
    8, 1, 18, 12, -1, -7, 8, -3, 10,
    -- layer=1 filter=178 channel=4
    9, 8, 15, 0, -3, 3, -13, -9, -9,
    -- layer=1 filter=178 channel=5
    4, 46, 7, 11, 11, 28, 13, 26, 8,
    -- layer=1 filter=178 channel=6
    19, 18, 4, -1, 16, 24, 12, 8, 29,
    -- layer=1 filter=178 channel=7
    -130, -126, -51, -87, -133, -70, -15, -108, -82,
    -- layer=1 filter=178 channel=8
    5, 27, -4, 18, 39, 31, 32, 53, 2,
    -- layer=1 filter=178 channel=9
    15, 26, 43, -56, 18, 30, -35, 7, -2,
    -- layer=1 filter=178 channel=10
    -104, -131, -37, -64, -127, -75, -6, -92, -108,
    -- layer=1 filter=178 channel=11
    13, 1, 15, -3, -10, -37, -3, -26, -50,
    -- layer=1 filter=178 channel=12
    63, 66, 73, -35, -49, 6, -6, 2, -41,
    -- layer=1 filter=178 channel=13
    9, 2, -6, 8, 24, 18, -1, 8, -4,
    -- layer=1 filter=178 channel=14
    -45, -30, 2, 5, -61, -10, -15, -82, -41,
    -- layer=1 filter=178 channel=15
    50, 56, 40, 38, 64, 74, 32, 71, 59,
    -- layer=1 filter=178 channel=16
    -7, 31, 1, 3, 14, 30, 1, 11, 2,
    -- layer=1 filter=178 channel=17
    29, -27, -75, 46, 17, -15, 51, 20, -24,
    -- layer=1 filter=178 channel=18
    18, 40, 9, 10, 10, 4, 7, 18, -17,
    -- layer=1 filter=178 channel=19
    -13, 12, -22, -44, -57, -2, -59, -53, -75,
    -- layer=1 filter=178 channel=20
    22, 8, -25, 15, 22, 3, 12, 16, 4,
    -- layer=1 filter=178 channel=21
    -15, 2, 22, -27, -11, 12, -26, -39, 12,
    -- layer=1 filter=178 channel=22
    16, 2, 1, 16, 16, 16, 26, 32, 14,
    -- layer=1 filter=178 channel=23
    -59, -7, -75, -58, -15, -31, -42, -26, -44,
    -- layer=1 filter=178 channel=24
    16, -4, 23, 6, -5, 13, -33, 14, 1,
    -- layer=1 filter=178 channel=25
    -118, -82, -40, -86, -36, -20, -36, -78, -71,
    -- layer=1 filter=178 channel=26
    42, 15, 17, 43, 42, 13, 10, 39, 9,
    -- layer=1 filter=178 channel=27
    32, 56, 33, 9, 32, 6, -20, -12, -8,
    -- layer=1 filter=178 channel=28
    -90, -140, -44, -80, -104, -51, 1, -88, -95,
    -- layer=1 filter=178 channel=29
    15, 15, 10, 14, 10, -9, 1, -22, -23,
    -- layer=1 filter=178 channel=30
    6, 6, 0, -15, -27, -2, 8, 6, -34,
    -- layer=1 filter=178 channel=31
    38, 20, 26, 7, -1, -5, 17, -6, 22,
    -- layer=1 filter=178 channel=32
    59, 21, 13, 14, 39, -5, 12, 41, 6,
    -- layer=1 filter=178 channel=33
    29, 6, 39, 23, 29, 5, 10, 5, -3,
    -- layer=1 filter=178 channel=34
    24, 30, 31, 43, 25, 38, 13, 7, 14,
    -- layer=1 filter=178 channel=35
    -7, 18, -39, 10, -20, 9, 12, 2, 16,
    -- layer=1 filter=178 channel=36
    12, -8, -10, 3, -27, -54, 14, -32, -55,
    -- layer=1 filter=178 channel=37
    -1, 29, 3, -18, 8, 22, 2, 3, -23,
    -- layer=1 filter=178 channel=38
    2, -6, -4, 6, -5, 6, 4, 9, -10,
    -- layer=1 filter=178 channel=39
    9, 18, 14, 21, -2, -7, 9, -8, -25,
    -- layer=1 filter=178 channel=40
    15, -6, -11, 4, -17, -6, 29, -9, 1,
    -- layer=1 filter=178 channel=41
    7, 11, 23, -23, 0, -21, -15, 2, -57,
    -- layer=1 filter=178 channel=42
    -30, 10, 50, -19, 5, 53, -32, -18, 29,
    -- layer=1 filter=178 channel=43
    -32, 0, -16, -28, -6, 9, -17, -11, -9,
    -- layer=1 filter=178 channel=44
    38, 11, 14, 37, 41, -4, 8, 36, 25,
    -- layer=1 filter=178 channel=45
    44, 18, 20, 17, 13, 18, -12, 16, 6,
    -- layer=1 filter=178 channel=46
    0, 50, 47, -17, 13, 49, 5, -10, -4,
    -- layer=1 filter=178 channel=47
    0, 35, 20, -41, 13, 4, -24, 3, 23,
    -- layer=1 filter=178 channel=48
    -10, -7, -4, 0, -3, 6, -12, -9, -13,
    -- layer=1 filter=178 channel=49
    -15, 25, 6, -16, -4, 14, -24, -10, 11,
    -- layer=1 filter=178 channel=50
    4, 16, 47, -26, -12, 2, 1, 5, 12,
    -- layer=1 filter=178 channel=51
    -24, -35, -13, -28, -50, -5, -8, -33, -45,
    -- layer=1 filter=178 channel=52
    -5, -4, -26, 29, 29, 18, 19, -10, -24,
    -- layer=1 filter=178 channel=53
    -12, 6, 2, -15, -11, 4, 5, -10, -6,
    -- layer=1 filter=178 channel=54
    -110, -39, -22, -79, -60, -26, -72, -82, -94,
    -- layer=1 filter=178 channel=55
    0, -8, 3, -17, -16, -1, 3, -8, 5,
    -- layer=1 filter=178 channel=56
    -2, 7, -4, 6, 3, 3, 1, 3, 0,
    -- layer=1 filter=178 channel=57
    -68, -96, -43, -31, -85, -47, 1, -51, -79,
    -- layer=1 filter=178 channel=58
    -189, -88, -66, -137, -119, -74, -63, -142, -95,
    -- layer=1 filter=178 channel=59
    0, -5, 6, -4, -3, 21, -8, 17, 3,
    -- layer=1 filter=178 channel=60
    35, 25, 18, -6, 3, 33, 2, 15, 35,
    -- layer=1 filter=178 channel=61
    0, -1, 2, 5, 8, 3, 10, 9, 12,
    -- layer=1 filter=178 channel=62
    11, 43, -7, 18, 15, 30, -4, 34, -18,
    -- layer=1 filter=178 channel=63
    12, 0, 0, -4, -34, -36, 7, -24, -37,
    -- layer=1 filter=178 channel=64
    2, 7, -4, 0, 20, 22, 15, 2, 4,
    -- layer=1 filter=178 channel=65
    -6, 4, 11, 0, 8, 0, 7, -5, -5,
    -- layer=1 filter=178 channel=66
    -2, -33, -48, 6, -46, -49, 14, -11, -28,
    -- layer=1 filter=178 channel=67
    19, 14, 24, -20, 0, 35, -9, 14, 45,
    -- layer=1 filter=178 channel=68
    59, 9, 23, 35, 23, -13, 16, 30, 12,
    -- layer=1 filter=178 channel=69
    33, 45, 29, 40, 45, 47, 2, 54, 9,
    -- layer=1 filter=178 channel=70
    23, 26, 9, 28, 5, 25, 11, 42, 39,
    -- layer=1 filter=178 channel=71
    -46, -11, -23, -59, -28, -18, -30, -12, -30,
    -- layer=1 filter=178 channel=72
    19, 23, 12, -22, -10, -10, -24, -2, -12,
    -- layer=1 filter=178 channel=73
    -12, 13, -16, -10, 7, 0, -2, 18, 1,
    -- layer=1 filter=178 channel=74
    19, 6, 11, -10, -8, -12, 6, -55, -20,
    -- layer=1 filter=178 channel=75
    39, 43, 9, -7, 7, 30, 37, -8, 19,
    -- layer=1 filter=178 channel=76
    20, -3, 15, 3, 9, -31, 24, 4, -41,
    -- layer=1 filter=178 channel=77
    0, -17, 13, 9, -1, 12, -10, -4, 5,
    -- layer=1 filter=178 channel=78
    -26, -22, -24, -22, -19, -26, 12, -13, -35,
    -- layer=1 filter=178 channel=79
    4, 48, 15, 10, 27, 30, 16, 44, 2,
    -- layer=1 filter=178 channel=80
    0, -1, -34, 36, 7, 19, -36, -11, 23,
    -- layer=1 filter=178 channel=81
    -11, -10, 11, -12, -14, 5, -20, -13, -6,
    -- layer=1 filter=178 channel=82
    -4, 8, 2, -18, -2, 16, -41, -13, 13,
    -- layer=1 filter=178 channel=83
    30, 4, -25, 60, 41, 21, 9, 52, 17,
    -- layer=1 filter=178 channel=84
    14, 8, 15, -35, -14, -25, 13, -22, -29,
    -- layer=1 filter=178 channel=85
    -63, -49, -39, -69, -58, -25, -49, -70, -27,
    -- layer=1 filter=178 channel=86
    -5, -30, -52, 11, -31, -56, 22, -9, -31,
    -- layer=1 filter=178 channel=87
    31, 60, 3, -40, -36, -38, -45, -41, 6,
    -- layer=1 filter=178 channel=88
    -18, 7, 21, -22, -6, 12, -22, -19, -3,
    -- layer=1 filter=178 channel=89
    -8, -6, 17, -10, 0, 11, -15, 0, 20,
    -- layer=1 filter=178 channel=90
    58, 24, 18, 59, 35, 33, 18, 59, 25,
    -- layer=1 filter=178 channel=91
    -8, 6, -15, 3, -1, -8, 2, 0, -8,
    -- layer=1 filter=178 channel=92
    25, 0, 55, 3, 26, 31, -32, 27, 34,
    -- layer=1 filter=178 channel=93
    -5, -11, -6, 3, -3, -15, -6, -8, -21,
    -- layer=1 filter=178 channel=94
    -15, -33, -46, 13, -32, -76, 27, -3, -29,
    -- layer=1 filter=178 channel=95
    7, 7, 15, -33, 9, 0, 23, -12, -23,
    -- layer=1 filter=178 channel=96
    -7, -9, 11, -4, -3, 1, -6, -3, 4,
    -- layer=1 filter=178 channel=97
    1, -31, -36, 12, -15, -25, 10, 9, -4,
    -- layer=1 filter=178 channel=98
    2, 7, -11, 9, 22, 41, 3, 28, -2,
    -- layer=1 filter=178 channel=99
    -39, -156, -64, -51, -154, -134, 19, -40, -144,
    -- layer=1 filter=178 channel=100
    28, 17, 16, 11, 7, 2, -1, -21, -28,
    -- layer=1 filter=178 channel=101
    1, -14, -19, 7, 5, -10, 8, -2, 1,
    -- layer=1 filter=178 channel=102
    -3, -43, -53, 31, 12, -19, 33, 24, -1,
    -- layer=1 filter=178 channel=103
    51, 38, 45, 13, 38, 25, 8, 0, -13,
    -- layer=1 filter=178 channel=104
    0, 33, 32, -29, 7, 0, 17, -6, -13,
    -- layer=1 filter=178 channel=105
    -4, -40, -61, 12, -45, -46, 24, 4, -43,
    -- layer=1 filter=178 channel=106
    14, 9, 7, 6, 34, 2, 4, 22, 9,
    -- layer=1 filter=178 channel=107
    5, 20, 5, 8, 23, 0, 7, 16, 15,
    -- layer=1 filter=178 channel=108
    44, 28, 36, 29, 44, 30, -5, 49, 40,
    -- layer=1 filter=178 channel=109
    -3, 7, -6, -9, -3, -7, 0, -1, 8,
    -- layer=1 filter=178 channel=110
    4, 22, 1, 7, -5, 0, 19, 7, -14,
    -- layer=1 filter=178 channel=111
    -5, 9, 12, -44, 4, -24, 11, -7, -46,
    -- layer=1 filter=178 channel=112
    38, 35, 27, 1, 9, -24, 9, -2, -22,
    -- layer=1 filter=178 channel=113
    24, 32, 54, 6, 10, 49, 8, 8, 12,
    -- layer=1 filter=178 channel=114
    8, 44, 22, 13, 27, 24, 38, 20, 10,
    -- layer=1 filter=178 channel=115
    -57, -85, -91, -34, -72, -58, 3, -39, -65,
    -- layer=1 filter=178 channel=116
    3, -4, 8, 0, -6, 2, 2, -6, 0,
    -- layer=1 filter=178 channel=117
    22, 28, 43, -16, 0, -43, -10, -25, -26,
    -- layer=1 filter=178 channel=118
    13, 5, -6, -28, -4, -24, 14, -14, -37,
    -- layer=1 filter=178 channel=119
    55, 13, 14, 29, 25, 14, 15, 51, 13,
    -- layer=1 filter=178 channel=120
    -21, 1, 23, -27, -7, 16, -31, -29, -4,
    -- layer=1 filter=178 channel=121
    23, 33, 17, -15, 13, 31, -12, -12, 6,
    -- layer=1 filter=178 channel=122
    3, -1, 0, -2, 0, 1, 3, 6, 8,
    -- layer=1 filter=178 channel=123
    -3, -7, 0, -23, 12, 14, -27, -32, -26,
    -- layer=1 filter=178 channel=124
    -4, 0, -2, 21, 18, 13, -3, 23, 8,
    -- layer=1 filter=178 channel=125
    24, 5, 23, -1, 0, 30, 14, 13, 30,
    -- layer=1 filter=178 channel=126
    4, -19, -25, 35, 48, 52, 16, 52, 27,
    -- layer=1 filter=178 channel=127
    26, 19, 11, -26, -25, -12, 4, 9, -26,
    -- layer=1 filter=179 channel=0
    -5, 4, -15, 5, 1, -2, -4, -6, 3,
    -- layer=1 filter=179 channel=1
    -5, -2, -4, -2, -9, 4, -8, -2, -7,
    -- layer=1 filter=179 channel=2
    1, -12, -13, 0, -18, 1, -8, 0, -13,
    -- layer=1 filter=179 channel=3
    3, 4, 3, 0, -9, 4, -8, -4, 4,
    -- layer=1 filter=179 channel=4
    4, 0, -4, 8, 0, 6, 6, -9, -6,
    -- layer=1 filter=179 channel=5
    -2, -9, 6, -2, 2, 12, 1, -8, 0,
    -- layer=1 filter=179 channel=6
    9, -11, -10, 10, 3, -11, -3, -5, -1,
    -- layer=1 filter=179 channel=7
    -18, -19, -7, -8, -5, -4, 1, -15, -8,
    -- layer=1 filter=179 channel=8
    -15, -10, -10, -6, -8, 6, -6, -9, -9,
    -- layer=1 filter=179 channel=9
    -3, 10, 3, 2, -4, -18, 0, 0, 1,
    -- layer=1 filter=179 channel=10
    -12, 0, 3, -12, -11, -3, 2, -1, -12,
    -- layer=1 filter=179 channel=11
    0, 5, 2, 6, 2, 5, 2, 0, 4,
    -- layer=1 filter=179 channel=12
    4, 3, -4, -8, -3, 0, 4, 10, 0,
    -- layer=1 filter=179 channel=13
    -6, -9, -14, 2, -9, -6, -3, -15, -1,
    -- layer=1 filter=179 channel=14
    5, -9, 3, -10, 2, -1, -7, -4, -9,
    -- layer=1 filter=179 channel=15
    0, 14, 0, 3, 8, -4, -11, 1, 4,
    -- layer=1 filter=179 channel=16
    1, -7, 7, -1, -2, -3, -12, -18, -12,
    -- layer=1 filter=179 channel=17
    5, 8, 0, -7, -5, -3, -12, -1, -3,
    -- layer=1 filter=179 channel=18
    2, -4, -5, -8, 0, -3, -11, -13, 1,
    -- layer=1 filter=179 channel=19
    -5, -1, 0, 0, -13, -3, 1, 4, 0,
    -- layer=1 filter=179 channel=20
    -6, 1, -8, 5, -4, -14, -3, -15, -6,
    -- layer=1 filter=179 channel=21
    -4, -7, -11, -17, -9, -1, -7, -1, -3,
    -- layer=1 filter=179 channel=22
    -9, -8, 4, -6, 0, -2, 0, -3, -15,
    -- layer=1 filter=179 channel=23
    -3, 10, -3, 8, -3, -6, 1, -2, -3,
    -- layer=1 filter=179 channel=24
    -4, -12, -18, -2, -8, -5, 0, -4, -10,
    -- layer=1 filter=179 channel=25
    -19, -6, 9, -11, -5, -3, 2, -19, -11,
    -- layer=1 filter=179 channel=26
    0, 0, 0, 2, 6, -11, 3, -2, 2,
    -- layer=1 filter=179 channel=27
    -1, 1, 13, 10, 4, -7, -9, -9, 0,
    -- layer=1 filter=179 channel=28
    -13, 1, -7, -1, 10, -12, -17, -11, -16,
    -- layer=1 filter=179 channel=29
    2, 1, 0, 0, -4, 3, 0, 8, -6,
    -- layer=1 filter=179 channel=30
    -2, -8, -1, 0, -5, -16, -4, -8, -12,
    -- layer=1 filter=179 channel=31
    -9, -7, 3, -5, -2, 6, -4, -8, 7,
    -- layer=1 filter=179 channel=32
    2, 13, -15, -1, 7, 3, 3, 9, -5,
    -- layer=1 filter=179 channel=33
    -7, 8, -5, -8, -12, 6, 7, 4, 7,
    -- layer=1 filter=179 channel=34
    -5, 0, 7, 5, -5, -9, 0, 0, 7,
    -- layer=1 filter=179 channel=35
    -10, 1, 1, -7, -12, -4, 0, 3, -4,
    -- layer=1 filter=179 channel=36
    14, 1, 0, -8, -4, -13, 5, -9, 9,
    -- layer=1 filter=179 channel=37
    -18, 0, -3, -8, 0, 12, -14, -11, -4,
    -- layer=1 filter=179 channel=38
    2, -9, -14, 10, -9, -16, 5, -9, -12,
    -- layer=1 filter=179 channel=39
    -8, -11, -1, -3, 8, -7, -4, 3, 6,
    -- layer=1 filter=179 channel=40
    10, -7, -13, -1, 0, 6, 7, -4, -2,
    -- layer=1 filter=179 channel=41
    4, 9, -12, 5, 2, -9, -2, 5, 2,
    -- layer=1 filter=179 channel=42
    4, -16, 5, -3, 0, -8, -2, -11, 1,
    -- layer=1 filter=179 channel=43
    -19, 0, 7, -8, 0, -4, 0, 0, -5,
    -- layer=1 filter=179 channel=44
    -2, 5, 3, -11, -1, 5, 5, 7, 3,
    -- layer=1 filter=179 channel=45
    -6, -10, -9, -13, -2, -15, -12, -6, -6,
    -- layer=1 filter=179 channel=46
    -15, 4, -4, 0, -5, 6, 1, -12, 9,
    -- layer=1 filter=179 channel=47
    -10, -1, 0, -10, -5, 3, -1, 10, -1,
    -- layer=1 filter=179 channel=48
    -10, -12, -8, -4, 1, -16, -8, 3, 0,
    -- layer=1 filter=179 channel=49
    3, -2, -9, -11, -6, -22, 8, 7, 0,
    -- layer=1 filter=179 channel=50
    -8, -6, -8, 8, -7, 6, 2, -5, -11,
    -- layer=1 filter=179 channel=51
    -20, -22, -10, -16, -10, -3, -13, 2, -16,
    -- layer=1 filter=179 channel=52
    7, -3, -9, -3, 6, 6, -4, -1, -2,
    -- layer=1 filter=179 channel=53
    -5, 4, -11, 6, -4, -6, -2, -6, -8,
    -- layer=1 filter=179 channel=54
    2, 0, -2, -9, 3, 12, 3, 3, -5,
    -- layer=1 filter=179 channel=55
    -17, 10, -4, -11, -1, -11, 1, 1, -15,
    -- layer=1 filter=179 channel=56
    8, 0, 0, 3, -7, 0, 2, 0, -4,
    -- layer=1 filter=179 channel=57
    -8, -16, 0, 3, -5, -1, 7, -14, -4,
    -- layer=1 filter=179 channel=58
    -13, -14, -1, -6, 2, -5, 2, -4, -2,
    -- layer=1 filter=179 channel=59
    -4, 3, -8, 1, 7, 8, 7, -4, -2,
    -- layer=1 filter=179 channel=60
    1, -5, -10, 2, -6, 0, 8, 8, -5,
    -- layer=1 filter=179 channel=61
    1, -6, -5, -4, 3, -3, 3, -2, 5,
    -- layer=1 filter=179 channel=62
    -9, -1, 10, -10, 0, 9, 2, -16, -4,
    -- layer=1 filter=179 channel=63
    3, 5, 1, 6, -2, -5, 5, -9, 8,
    -- layer=1 filter=179 channel=64
    -14, -1, -5, -13, 1, -10, -1, -9, -15,
    -- layer=1 filter=179 channel=65
    -11, -3, -9, 5, -10, -9, -13, -11, 2,
    -- layer=1 filter=179 channel=66
    -1, 0, -2, -7, 1, 4, -15, -5, 1,
    -- layer=1 filter=179 channel=67
    -1, 1, -1, -11, 1, 9, -11, 4, 7,
    -- layer=1 filter=179 channel=68
    12, -7, -11, 7, 2, 0, -13, -11, -9,
    -- layer=1 filter=179 channel=69
    -14, -3, 4, -16, -2, 13, -4, -17, -4,
    -- layer=1 filter=179 channel=70
    5, 7, 5, 6, 1, -4, 2, 1, -8,
    -- layer=1 filter=179 channel=71
    -20, -19, -5, -6, 1, 0, -9, 2, -5,
    -- layer=1 filter=179 channel=72
    -13, -10, 0, 0, -4, -4, -11, -9, 9,
    -- layer=1 filter=179 channel=73
    -6, 9, 0, -2, -4, 3, 8, -9, 7,
    -- layer=1 filter=179 channel=74
    -4, -7, -6, -8, -3, 5, -9, -19, 5,
    -- layer=1 filter=179 channel=75
    -3, -12, -7, -8, -13, 9, 4, -13, 1,
    -- layer=1 filter=179 channel=76
    8, 3, -3, 6, -2, 9, -4, 4, -3,
    -- layer=1 filter=179 channel=77
    -8, 1, -15, -8, 6, -2, -14, -7, -7,
    -- layer=1 filter=179 channel=78
    2, 8, 3, -14, -8, 1, -10, 1, -2,
    -- layer=1 filter=179 channel=79
    -1, 0, -10, -11, -13, -5, -11, -4, -13,
    -- layer=1 filter=179 channel=80
    -4, -6, 3, -3, -7, 1, 6, -1, 0,
    -- layer=1 filter=179 channel=81
    -17, -6, -2, -2, 5, 0, -9, -11, -5,
    -- layer=1 filter=179 channel=82
    -8, -4, -15, -15, -14, -16, -7, -7, -3,
    -- layer=1 filter=179 channel=83
    -10, 5, 9, -11, -2, -10, 2, -8, -3,
    -- layer=1 filter=179 channel=84
    -2, 4, -10, 0, 0, 3, -17, -9, 10,
    -- layer=1 filter=179 channel=85
    -2, 1, 12, -5, 6, 4, 2, -9, -12,
    -- layer=1 filter=179 channel=86
    0, -1, -4, -9, -9, -6, -9, -4, 3,
    -- layer=1 filter=179 channel=87
    -8, -7, -3, 7, 3, 4, -6, -1, 0,
    -- layer=1 filter=179 channel=88
    -14, -15, -6, -9, -15, -14, -8, -17, -7,
    -- layer=1 filter=179 channel=89
    0, 1, -7, -15, 1, -9, 0, -7, -10,
    -- layer=1 filter=179 channel=90
    1, -9, -7, -8, -4, 5, 0, -11, 1,
    -- layer=1 filter=179 channel=91
    6, -11, -1, 9, -3, -21, 0, -2, -19,
    -- layer=1 filter=179 channel=92
    -14, 2, -6, -13, 2, -8, -11, -9, -9,
    -- layer=1 filter=179 channel=93
    -17, -2, -13, -1, -18, -11, -13, -1, -18,
    -- layer=1 filter=179 channel=94
    -4, 0, -13, -15, -9, -2, -1, -5, -9,
    -- layer=1 filter=179 channel=95
    -9, 4, 0, -4, -11, -3, -11, -12, 5,
    -- layer=1 filter=179 channel=96
    -6, 5, 1, -2, -4, 4, -6, -9, 0,
    -- layer=1 filter=179 channel=97
    -7, -9, -6, -15, -3, -14, -3, 1, 5,
    -- layer=1 filter=179 channel=98
    -9, -5, 4, -5, 7, 0, 1, -12, -5,
    -- layer=1 filter=179 channel=99
    -12, -5, -6, -4, 7, 2, 2, 3, -12,
    -- layer=1 filter=179 channel=100
    10, -5, 0, 2, -15, -2, 0, -15, 0,
    -- layer=1 filter=179 channel=101
    -11, -12, -25, -3, -17, -14, -5, -15, -14,
    -- layer=1 filter=179 channel=102
    1, -6, -11, -3, -11, -9, -5, 0, -11,
    -- layer=1 filter=179 channel=103
    6, -4, -11, -1, 1, 5, -3, -7, 5,
    -- layer=1 filter=179 channel=104
    -9, 7, -5, -12, 7, -8, -2, -8, -13,
    -- layer=1 filter=179 channel=105
    -14, -10, -6, -15, -11, -11, -17, 8, -8,
    -- layer=1 filter=179 channel=106
    0, -5, -14, 10, 0, -2, 2, 6, -19,
    -- layer=1 filter=179 channel=107
    -7, -8, -4, 5, -7, 0, 6, -6, 8,
    -- layer=1 filter=179 channel=108
    0, 6, 7, -3, -1, 4, -3, 0, -18,
    -- layer=1 filter=179 channel=109
    3, -4, 0, -6, -10, -4, 2, -5, -9,
    -- layer=1 filter=179 channel=110
    -7, -11, -6, -2, 0, 0, -9, -1, 0,
    -- layer=1 filter=179 channel=111
    -3, 6, -7, 4, 9, 3, -15, -17, 0,
    -- layer=1 filter=179 channel=112
    -8, 2, 1, 0, -3, -4, -19, -1, 3,
    -- layer=1 filter=179 channel=113
    -11, 7, 3, 10, 5, 1, 7, -14, -6,
    -- layer=1 filter=179 channel=114
    -7, -7, 16, -11, 4, 4, -14, -10, -10,
    -- layer=1 filter=179 channel=115
    -3, -8, -5, -14, 4, 4, 3, 6, -14,
    -- layer=1 filter=179 channel=116
    0, 8, 5, 3, 9, -3, -9, -1, 0,
    -- layer=1 filter=179 channel=117
    -8, -4, -7, 2, 8, 11, -3, 10, -11,
    -- layer=1 filter=179 channel=118
    -5, -10, -5, -6, 3, 4, -4, 0, -7,
    -- layer=1 filter=179 channel=119
    2, 3, -4, -3, 1, -15, -3, 7, -10,
    -- layer=1 filter=179 channel=120
    -17, -20, 3, -12, -9, -18, -13, -2, -16,
    -- layer=1 filter=179 channel=121
    -15, -17, -13, 0, -13, -19, 4, -12, -11,
    -- layer=1 filter=179 channel=122
    0, 0, -1, 9, 8, 3, -1, 10, 3,
    -- layer=1 filter=179 channel=123
    -11, 0, 4, -7, 0, -16, -10, 3, -11,
    -- layer=1 filter=179 channel=124
    -2, -7, 0, -7, -9, 4, -7, -3, -1,
    -- layer=1 filter=179 channel=125
    3, 4, 0, 6, 8, 5, 3, -9, 0,
    -- layer=1 filter=179 channel=126
    -8, -6, 5, -11, -8, 0, -18, -16, 7,
    -- layer=1 filter=179 channel=127
    -8, -5, -6, 0, -2, 4, -11, -7, 3,
    -- layer=1 filter=180 channel=0
    8, -4, 5, -2, 4, -8, 1, -7, -5,
    -- layer=1 filter=180 channel=1
    1, 2, -3, 3, 4, 7, -8, 7, 7,
    -- layer=1 filter=180 channel=2
    -10, 2, -5, -3, 8, 1, -3, -6, -9,
    -- layer=1 filter=180 channel=3
    6, 8, -10, 1, 6, 0, 0, 0, 7,
    -- layer=1 filter=180 channel=4
    2, -8, 0, -4, -1, 5, 2, 7, 4,
    -- layer=1 filter=180 channel=5
    -15, 4, 0, -11, -14, -8, -4, 3, -8,
    -- layer=1 filter=180 channel=6
    3, -9, 5, 4, 4, 0, 3, -9, 8,
    -- layer=1 filter=180 channel=7
    -4, -7, 2, -2, 2, -6, -8, -11, -9,
    -- layer=1 filter=180 channel=8
    9, -5, 0, 5, -5, -5, 8, 2, 1,
    -- layer=1 filter=180 channel=9
    7, 5, 5, -5, 2, -6, 7, 3, 0,
    -- layer=1 filter=180 channel=10
    -10, 0, -2, 2, 5, -11, -4, -3, -1,
    -- layer=1 filter=180 channel=11
    -10, 0, 7, 6, -3, 5, -10, 6, -5,
    -- layer=1 filter=180 channel=12
    7, 2, -2, -6, -5, -3, -6, 2, -7,
    -- layer=1 filter=180 channel=13
    6, -3, 6, 7, -1, -9, 1, 0, -6,
    -- layer=1 filter=180 channel=14
    9, 0, 0, -6, -3, 9, -4, -1, 0,
    -- layer=1 filter=180 channel=15
    -7, 8, 9, -7, -2, -3, 8, 9, 9,
    -- layer=1 filter=180 channel=16
    -14, 4, -9, -3, -1, -1, -4, -10, -2,
    -- layer=1 filter=180 channel=17
    4, -9, 0, 1, 0, -3, -7, -1, 7,
    -- layer=1 filter=180 channel=18
    8, 7, -5, 2, 2, 6, 1, -9, 0,
    -- layer=1 filter=180 channel=19
    7, 0, -8, 5, 0, -3, 5, 3, -1,
    -- layer=1 filter=180 channel=20
    -8, 8, -9, 0, 1, -2, 7, 0, -9,
    -- layer=1 filter=180 channel=21
    6, -2, 0, 4, 4, -12, -6, 2, -4,
    -- layer=1 filter=180 channel=22
    -7, -2, -4, 1, -4, 0, 2, 0, -4,
    -- layer=1 filter=180 channel=23
    6, -3, -4, -1, 1, 4, 1, -9, 2,
    -- layer=1 filter=180 channel=24
    -14, 7, 6, -11, 6, -13, 1, 0, -3,
    -- layer=1 filter=180 channel=25
    -5, 1, -5, -12, -12, -2, 8, 3, -8,
    -- layer=1 filter=180 channel=26
    7, -4, 3, -4, 0, 4, -9, -3, -5,
    -- layer=1 filter=180 channel=27
    -5, -1, 2, -7, -7, 7, -5, -3, 7,
    -- layer=1 filter=180 channel=28
    8, -6, 3, -13, -3, 5, -1, 0, -5,
    -- layer=1 filter=180 channel=29
    9, -7, -7, -1, 0, -10, 0, -10, 1,
    -- layer=1 filter=180 channel=30
    -6, -5, 2, 0, -12, 0, -6, 3, -15,
    -- layer=1 filter=180 channel=31
    -4, 6, 4, -10, 1, 0, 6, 0, 0,
    -- layer=1 filter=180 channel=32
    2, -11, -7, -1, -6, 1, -11, 5, 4,
    -- layer=1 filter=180 channel=33
    7, 0, 7, 0, -10, 7, 7, 5, 10,
    -- layer=1 filter=180 channel=34
    -7, 1, -1, -8, -2, 9, 8, 4, 7,
    -- layer=1 filter=180 channel=35
    0, 2, -4, 0, 7, -5, 2, -3, -11,
    -- layer=1 filter=180 channel=36
    -4, -8, 2, 0, 1, 5, 1, 7, 9,
    -- layer=1 filter=180 channel=37
    0, 0, -8, 0, 6, -3, -5, -7, 0,
    -- layer=1 filter=180 channel=38
    3, -13, 1, 3, -9, 2, -5, 0, -10,
    -- layer=1 filter=180 channel=39
    8, -10, -6, 0, -8, -6, 7, -10, 2,
    -- layer=1 filter=180 channel=40
    8, 5, -3, 6, -4, -6, -3, -6, -5,
    -- layer=1 filter=180 channel=41
    -1, -10, 3, -8, -5, -11, -7, -11, 6,
    -- layer=1 filter=180 channel=42
    -3, -8, -9, 0, 2, 0, 9, 5, 0,
    -- layer=1 filter=180 channel=43
    1, 7, -2, 1, -1, -11, 1, 2, 1,
    -- layer=1 filter=180 channel=44
    0, -5, 3, -7, 5, 4, -4, 0, 8,
    -- layer=1 filter=180 channel=45
    6, 1, -1, -13, 6, -11, -3, 4, -7,
    -- layer=1 filter=180 channel=46
    -4, -11, 3, 2, -6, 8, 7, 1, -9,
    -- layer=1 filter=180 channel=47
    -9, 6, 3, -12, -4, -5, -6, 7, -5,
    -- layer=1 filter=180 channel=48
    2, -4, 7, -10, 5, 4, -12, -10, 0,
    -- layer=1 filter=180 channel=49
    1, -3, -12, -9, -13, -5, -13, 7, 1,
    -- layer=1 filter=180 channel=50
    0, -6, -7, -4, 0, 2, -8, -6, 1,
    -- layer=1 filter=180 channel=51
    2, 0, -8, -6, -8, -5, -4, -5, 0,
    -- layer=1 filter=180 channel=52
    -1, 7, -8, 10, -11, -4, -3, 2, 0,
    -- layer=1 filter=180 channel=53
    -9, -6, -4, -1, 9, 5, 0, -1, 5,
    -- layer=1 filter=180 channel=54
    0, -1, -11, 1, -8, 5, 1, -8, -7,
    -- layer=1 filter=180 channel=55
    5, 1, -2, 10, -1, 3, -4, -1, 8,
    -- layer=1 filter=180 channel=56
    -9, 2, -3, -3, 9, 4, 5, 2, -12,
    -- layer=1 filter=180 channel=57
    -6, -7, -8, 7, -7, -2, -10, -3, 8,
    -- layer=1 filter=180 channel=58
    -16, -1, -4, 0, 7, -12, 6, -2, -4,
    -- layer=1 filter=180 channel=59
    -1, 8, -3, 0, 4, -9, -11, -5, 4,
    -- layer=1 filter=180 channel=60
    -1, 2, -11, -3, 1, -3, 4, 1, 8,
    -- layer=1 filter=180 channel=61
    3, 2, 7, 7, -3, 8, 2, -3, 8,
    -- layer=1 filter=180 channel=62
    -9, -4, -18, -9, -12, 2, -12, 6, -9,
    -- layer=1 filter=180 channel=63
    3, -4, 4, -3, -3, -10, -5, 0, -8,
    -- layer=1 filter=180 channel=64
    -10, 1, -6, -3, 4, 2, -2, 0, -1,
    -- layer=1 filter=180 channel=65
    -8, 8, -5, -11, 0, -9, -5, -11, 2,
    -- layer=1 filter=180 channel=66
    2, 0, -4, 8, 4, -5, -7, -6, -4,
    -- layer=1 filter=180 channel=67
    -4, 4, -3, 11, 0, 8, 11, -9, 4,
    -- layer=1 filter=180 channel=68
    -11, -9, -11, 1, -12, -5, -7, 4, 4,
    -- layer=1 filter=180 channel=69
    3, -14, 3, -8, 5, 5, 2, -10, 2,
    -- layer=1 filter=180 channel=70
    8, 6, 0, 12, 1, -8, -1, 11, 1,
    -- layer=1 filter=180 channel=71
    7, -8, 5, -7, -10, 0, -11, -7, -5,
    -- layer=1 filter=180 channel=72
    -2, 5, 0, -6, -3, -7, 0, -5, 5,
    -- layer=1 filter=180 channel=73
    7, -7, -6, 6, -4, -2, 0, -3, 0,
    -- layer=1 filter=180 channel=74
    4, 7, -11, -5, -3, -2, 1, -7, -9,
    -- layer=1 filter=180 channel=75
    4, -8, -1, 4, -9, -3, -4, -14, 2,
    -- layer=1 filter=180 channel=76
    7, 5, 3, -6, 6, -6, -5, -9, 5,
    -- layer=1 filter=180 channel=77
    3, -2, -11, -4, 6, 4, -3, 0, -3,
    -- layer=1 filter=180 channel=78
    6, -1, -8, -10, 1, 4, 8, 7, 1,
    -- layer=1 filter=180 channel=79
    3, 6, -3, -4, -11, 3, -10, -8, 0,
    -- layer=1 filter=180 channel=80
    -9, -6, -2, 6, -8, -11, 5, -5, -5,
    -- layer=1 filter=180 channel=81
    -1, 5, -11, -9, -5, -8, -2, -2, -2,
    -- layer=1 filter=180 channel=82
    -12, -1, -9, 5, 7, -8, -14, -5, -4,
    -- layer=1 filter=180 channel=83
    -10, 2, -10, 3, -1, -3, -7, 5, -3,
    -- layer=1 filter=180 channel=84
    9, -5, 1, -6, -15, -11, -9, -2, -4,
    -- layer=1 filter=180 channel=85
    -5, -9, -13, -1, -7, -11, 9, -9, -1,
    -- layer=1 filter=180 channel=86
    1, -9, 4, -2, 5, -5, 0, -8, -8,
    -- layer=1 filter=180 channel=87
    -8, 0, -9, -9, 5, -5, 1, -7, -8,
    -- layer=1 filter=180 channel=88
    -14, -4, 8, 2, 0, 3, -3, 4, 4,
    -- layer=1 filter=180 channel=89
    7, -2, -11, 1, -7, -2, -10, 1, 3,
    -- layer=1 filter=180 channel=90
    4, -5, -2, -6, -10, -1, -11, -12, -10,
    -- layer=1 filter=180 channel=91
    6, 4, -8, 5, -4, -5, -3, -11, -5,
    -- layer=1 filter=180 channel=92
    -7, 5, -11, -11, 8, 8, -8, 0, -3,
    -- layer=1 filter=180 channel=93
    0, -6, 0, 3, -8, -9, 0, -10, 5,
    -- layer=1 filter=180 channel=94
    4, -2, 1, -3, -2, 8, -4, -1, 1,
    -- layer=1 filter=180 channel=95
    5, -9, -11, 0, 1, 0, 4, -2, -7,
    -- layer=1 filter=180 channel=96
    -8, 0, 7, -1, 3, 7, -7, -1, 2,
    -- layer=1 filter=180 channel=97
    7, 6, -3, 1, -9, 2, 1, -7, 1,
    -- layer=1 filter=180 channel=98
    3, 1, -4, -7, -9, -9, -8, -4, 0,
    -- layer=1 filter=180 channel=99
    2, -9, 5, -8, 5, -11, -6, 0, -2,
    -- layer=1 filter=180 channel=100
    -9, 1, -6, 4, -1, -8, 8, -9, 5,
    -- layer=1 filter=180 channel=101
    -11, -2, 1, -3, 0, 7, -5, -1, 6,
    -- layer=1 filter=180 channel=102
    1, -2, -11, -2, -3, 2, 8, 0, -2,
    -- layer=1 filter=180 channel=103
    9, 1, 8, 0, 6, -7, 6, 4, -4,
    -- layer=1 filter=180 channel=104
    -4, -8, -5, -10, -8, -5, -4, 4, -8,
    -- layer=1 filter=180 channel=105
    -11, 1, -3, 1, -6, 4, -11, -8, 0,
    -- layer=1 filter=180 channel=106
    -5, 2, -5, 5, -9, 3, 1, 2, 1,
    -- layer=1 filter=180 channel=107
    4, -5, 0, -1, 3, -5, 8, 1, 0,
    -- layer=1 filter=180 channel=108
    1, 8, -4, 0, 10, 0, -5, -12, -2,
    -- layer=1 filter=180 channel=109
    0, -8, -1, 7, -3, 9, 0, 9, -2,
    -- layer=1 filter=180 channel=110
    -8, 6, -11, 5, -11, 2, -2, -2, 4,
    -- layer=1 filter=180 channel=111
    -4, 2, -7, -5, 3, 0, -10, 0, -3,
    -- layer=1 filter=180 channel=112
    -4, -3, 4, -6, 6, -3, 0, 6, 7,
    -- layer=1 filter=180 channel=113
    1, -9, -12, -10, 6, 1, -6, -1, -1,
    -- layer=1 filter=180 channel=114
    -13, -4, 0, 0, 0, -9, -11, 1, 1,
    -- layer=1 filter=180 channel=115
    -5, -1, -4, -3, -1, -2, -2, 0, 8,
    -- layer=1 filter=180 channel=116
    9, 5, 7, 6, 4, -3, 1, 0, -7,
    -- layer=1 filter=180 channel=117
    0, -7, -1, 6, -19, 0, -4, 0, -11,
    -- layer=1 filter=180 channel=118
    0, -9, -11, 4, -12, -6, 4, -5, -11,
    -- layer=1 filter=180 channel=119
    -3, -3, -4, -6, -7, -8, -4, 0, -8,
    -- layer=1 filter=180 channel=120
    6, 7, -4, -3, -6, -7, -6, -9, 4,
    -- layer=1 filter=180 channel=121
    1, -5, 9, 8, 9, -6, -6, 6, -11,
    -- layer=1 filter=180 channel=122
    1, 0, -1, 9, 5, -5, 3, 5, 8,
    -- layer=1 filter=180 channel=123
    7, -1, 2, 7, 6, 4, -5, -5, -1,
    -- layer=1 filter=180 channel=124
    0, 3, 1, -6, -3, 0, -1, -5, 5,
    -- layer=1 filter=180 channel=125
    7, -8, -6, -1, 3, -1, -8, -4, 4,
    -- layer=1 filter=180 channel=126
    -6, 1, -7, -2, 7, 2, 1, 0, -5,
    -- layer=1 filter=180 channel=127
    -7, 4, 5, -9, -11, -10, 2, -12, -13,
    -- layer=1 filter=181 channel=0
    -7, -7, 21, 9, -2, 18, 8, -7, 0,
    -- layer=1 filter=181 channel=1
    -5, -11, -26, -20, 4, 5, -18, 7, -13,
    -- layer=1 filter=181 channel=2
    14, 0, 6, 0, 3, -41, -12, 0, -15,
    -- layer=1 filter=181 channel=3
    -8, -2, 0, 5, -13, 0, -2, 5, -13,
    -- layer=1 filter=181 channel=4
    8, 1, 0, -2, 17, 6, 1, -13, -8,
    -- layer=1 filter=181 channel=5
    10, -41, -27, -13, -5, 1, -22, 16, 1,
    -- layer=1 filter=181 channel=6
    -15, 5, -9, -4, -3, 9, -4, -13, 6,
    -- layer=1 filter=181 channel=7
    -2, 58, 13, 3, 70, 48, 33, 55, 45,
    -- layer=1 filter=181 channel=8
    6, -59, -19, -19, -28, -11, 0, -2, -7,
    -- layer=1 filter=181 channel=9
    11, -29, -47, -4, 38, -28, 10, 3, -42,
    -- layer=1 filter=181 channel=10
    -29, 43, 25, -16, 58, 38, 0, 36, 26,
    -- layer=1 filter=181 channel=11
    -6, -5, 10, -9, -3, -12, 14, 1, -10,
    -- layer=1 filter=181 channel=12
    -25, -11, 26, -43, 6, 28, 32, -40, 43,
    -- layer=1 filter=181 channel=13
    -4, -2, -23, 3, 13, -32, -10, 6, -22,
    -- layer=1 filter=181 channel=14
    -32, 12, 1, -1, 30, 8, 26, 24, 36,
    -- layer=1 filter=181 channel=15
    19, 23, 28, 9, 30, -16, -17, 21, -9,
    -- layer=1 filter=181 channel=16
    -1, -33, -6, -22, -22, -17, -16, 5, -8,
    -- layer=1 filter=181 channel=17
    -3, -15, 20, 4, -15, -4, -10, -18, -8,
    -- layer=1 filter=181 channel=18
    2, 7, 16, -9, -25, 18, 4, -5, 6,
    -- layer=1 filter=181 channel=19
    -2, 0, 19, -10, -14, -18, -4, -19, -8,
    -- layer=1 filter=181 channel=20
    6, -5, -2, -7, -3, -16, -19, -20, -3,
    -- layer=1 filter=181 channel=21
    -8, -3, -3, -22, -35, 8, -10, -17, 12,
    -- layer=1 filter=181 channel=22
    -3, 4, 7, -14, -13, -15, -14, -8, -16,
    -- layer=1 filter=181 channel=23
    -1, 83, -55, 28, 108, 21, 14, 69, 26,
    -- layer=1 filter=181 channel=24
    7, -38, -18, 12, 1, -51, 4, -5, -44,
    -- layer=1 filter=181 channel=25
    0, 39, -10, 3, 46, 20, 5, 27, 17,
    -- layer=1 filter=181 channel=26
    21, 22, -59, 17, 48, -100, 0, 46, -61,
    -- layer=1 filter=181 channel=27
    13, 15, 30, -45, -25, -9, -40, -24, 14,
    -- layer=1 filter=181 channel=28
    -23, 41, 17, -15, 44, 35, 7, 18, 30,
    -- layer=1 filter=181 channel=29
    19, 15, 35, -4, -9, 24, -6, 6, 10,
    -- layer=1 filter=181 channel=30
    -16, 7, 38, -25, -13, -8, -5, -26, -29,
    -- layer=1 filter=181 channel=31
    -17, 16, 5, -6, -13, 0, -12, -10, 0,
    -- layer=1 filter=181 channel=32
    6, 37, -101, 3, 75, -71, 2, 74, -35,
    -- layer=1 filter=181 channel=33
    -6, 0, 1, -6, -30, -20, 0, -4, -9,
    -- layer=1 filter=181 channel=34
    -14, -18, -5, -15, -4, -30, -7, -11, -29,
    -- layer=1 filter=181 channel=35
    -15, 9, 13, -8, 27, 27, 1, 4, -7,
    -- layer=1 filter=181 channel=36
    12, 0, 16, -6, -6, -8, 19, -3, 0,
    -- layer=1 filter=181 channel=37
    6, -46, -2, -29, -21, -8, -16, -10, 0,
    -- layer=1 filter=181 channel=38
    -3, -12, 25, -20, -12, -1, -11, -11, 0,
    -- layer=1 filter=181 channel=39
    1, -10, -6, -7, -19, -19, -16, 0, 0,
    -- layer=1 filter=181 channel=40
    -12, 5, 37, -12, -15, 11, -13, -27, 4,
    -- layer=1 filter=181 channel=41
    -4, 12, -79, -37, 65, -87, 0, 58, -5,
    -- layer=1 filter=181 channel=42
    16, 13, 1, -7, 12, 7, 8, 4, -8,
    -- layer=1 filter=181 channel=43
    -9, -10, -30, -20, -21, 1, -14, 9, 4,
    -- layer=1 filter=181 channel=44
    23, 45, -76, 26, 70, -87, -9, 46, -54,
    -- layer=1 filter=181 channel=45
    16, -11, -8, -1, -9, -13, -1, -9, -22,
    -- layer=1 filter=181 channel=46
    -3, 0, 0, -24, -25, 3, 12, -16, 0,
    -- layer=1 filter=181 channel=47
    18, 77, -89, 18, 75, -47, 0, 44, -24,
    -- layer=1 filter=181 channel=48
    -2, -19, 7, -13, -21, 9, -16, -32, -1,
    -- layer=1 filter=181 channel=49
    -1, -10, -7, -5, 13, -21, -5, -8, -13,
    -- layer=1 filter=181 channel=50
    -28, -8, -19, -10, -10, -22, -19, -13, -26,
    -- layer=1 filter=181 channel=51
    -11, 1, 14, -12, -1, 17, -6, -9, 23,
    -- layer=1 filter=181 channel=52
    25, 16, -3, -8, 11, -2, 2, 7, 0,
    -- layer=1 filter=181 channel=53
    6, 5, 0, 8, 0, 16, -16, 14, 2,
    -- layer=1 filter=181 channel=54
    -9, 21, -7, 6, 40, -7, -8, 11, 7,
    -- layer=1 filter=181 channel=55
    -13, 2, -8, -2, 8, -3, 13, 0, -3,
    -- layer=1 filter=181 channel=56
    9, 11, 6, 0, -1, 11, 6, 13, 5,
    -- layer=1 filter=181 channel=57
    -10, 47, 28, -25, 42, 42, -9, 19, 17,
    -- layer=1 filter=181 channel=58
    39, 104, 2, 55, 110, 53, 49, 58, 50,
    -- layer=1 filter=181 channel=59
    -34, -18, -19, -25, -5, -13, -38, -27, -20,
    -- layer=1 filter=181 channel=60
    -10, 2, 19, 8, 0, -9, -2, 27, -13,
    -- layer=1 filter=181 channel=61
    -15, 18, -9, 1, 0, 1, -1, -7, -16,
    -- layer=1 filter=181 channel=62
    -12, -31, -13, -21, -6, -7, -19, 8, -17,
    -- layer=1 filter=181 channel=63
    10, 10, 0, -4, -10, 0, 21, -3, 0,
    -- layer=1 filter=181 channel=64
    -5, 0, 3, -23, -11, 16, -3, -3, 15,
    -- layer=1 filter=181 channel=65
    -7, -15, 18, -16, -31, 18, -17, -25, 16,
    -- layer=1 filter=181 channel=66
    6, -2, 3, 10, 3, 5, 0, -8, 2,
    -- layer=1 filter=181 channel=67
    -10, -34, -6, -33, -36, 6, 19, -22, 7,
    -- layer=1 filter=181 channel=68
    38, 22, -44, 48, 46, -18, 12, 58, -27,
    -- layer=1 filter=181 channel=69
    4, 14, -7, -14, 15, -28, -16, 7, -31,
    -- layer=1 filter=181 channel=70
    -17, 0, -7, -27, 14, 15, -3, -6, 9,
    -- layer=1 filter=181 channel=71
    4, 3, 4, -18, -9, 13, -27, -1, 13,
    -- layer=1 filter=181 channel=72
    6, 28, 36, -6, 2, 10, -2, -24, -11,
    -- layer=1 filter=181 channel=73
    0, -8, -4, 7, -15, -13, -2, -13, 2,
    -- layer=1 filter=181 channel=74
    0, 6, 24, 28, -20, 35, 10, 34, 25,
    -- layer=1 filter=181 channel=75
    -28, 20, 9, -10, 13, -5, -11, -47, -1,
    -- layer=1 filter=181 channel=76
    6, 1, -11, 10, 2, -15, 16, 16, -19,
    -- layer=1 filter=181 channel=77
    0, -34, 7, 0, -29, 18, -11, -19, -1,
    -- layer=1 filter=181 channel=78
    -31, 4, 12, -20, -5, 9, -16, -14, 4,
    -- layer=1 filter=181 channel=79
    -14, -20, -14, -7, -6, -17, -13, 0, -13,
    -- layer=1 filter=181 channel=80
    1, -13, 3, -4, -4, 18, -4, 14, 1,
    -- layer=1 filter=181 channel=81
    -12, -8, -4, -19, -39, 2, 1, -25, 5,
    -- layer=1 filter=181 channel=82
    -13, -8, -4, -16, -14, 13, -23, -13, 6,
    -- layer=1 filter=181 channel=83
    5, 11, -1, 9, -5, -25, -17, 8, -12,
    -- layer=1 filter=181 channel=84
    13, -4, -26, 14, -5, -35, 14, 15, -16,
    -- layer=1 filter=181 channel=85
    32, 70, -44, 23, 86, -14, 16, 46, 7,
    -- layer=1 filter=181 channel=86
    -11, -9, 2, -8, -9, 0, 3, 0, 10,
    -- layer=1 filter=181 channel=87
    11, 0, -5, 28, 9, 11, 41, -7, -24,
    -- layer=1 filter=181 channel=88
    4, -20, 0, 10, -8, -1, 2, -15, 4,
    -- layer=1 filter=181 channel=89
    0, 0, -1, 0, -26, 1, -17, -26, -18,
    -- layer=1 filter=181 channel=90
    34, 23, -34, 23, 55, -49, 12, 66, -21,
    -- layer=1 filter=181 channel=91
    -9, 9, 12, -28, 1, 15, -4, -12, 8,
    -- layer=1 filter=181 channel=92
    -12, 34, -51, 6, 31, -35, -27, 0, -16,
    -- layer=1 filter=181 channel=93
    -11, -11, 7, -5, -22, -4, -13, -23, -5,
    -- layer=1 filter=181 channel=94
    -6, 13, 25, -8, -2, 3, 9, -5, -6,
    -- layer=1 filter=181 channel=95
    -14, 15, -9, -4, -18, -7, 13, -18, -5,
    -- layer=1 filter=181 channel=96
    5, -7, -19, -2, -6, -22, -1, -17, -14,
    -- layer=1 filter=181 channel=97
    5, -18, 3, 5, -15, -2, -13, -7, -9,
    -- layer=1 filter=181 channel=98
    -2, -27, -7, -29, -23, 13, -20, 9, 5,
    -- layer=1 filter=181 channel=99
    4, 31, 53, 33, 54, 96, 9, 78, 67,
    -- layer=1 filter=181 channel=100
    -11, 12, -6, -9, -7, 4, -17, -5, 8,
    -- layer=1 filter=181 channel=101
    1, 0, 5, -11, -12, 0, -10, -12, 11,
    -- layer=1 filter=181 channel=102
    11, 17, 18, -9, 4, 0, -21, -17, -12,
    -- layer=1 filter=181 channel=103
    -10, -9, 8, -34, -36, 5, 8, 3, 7,
    -- layer=1 filter=181 channel=104
    -1, 28, -46, -6, 51, -27, 9, 32, 4,
    -- layer=1 filter=181 channel=105
    -8, -4, 22, -6, -7, 8, 9, -1, 2,
    -- layer=1 filter=181 channel=106
    7, 0, -48, -2, 14, -31, 2, -5, -27,
    -- layer=1 filter=181 channel=107
    -7, 22, 17, 6, -1, 6, 1, 11, 14,
    -- layer=1 filter=181 channel=108
    10, 39, -98, 20, 81, -68, -1, 66, -32,
    -- layer=1 filter=181 channel=109
    4, 0, 5, 1, -9, -6, 3, -11, -2,
    -- layer=1 filter=181 channel=110
    -1, -10, 7, -18, -9, 5, -15, -4, 9,
    -- layer=1 filter=181 channel=111
    -15, -5, 25, -16, -41, 0, 1, -21, -4,
    -- layer=1 filter=181 channel=112
    -23, -1, -15, -16, -27, -12, 10, -6, -2,
    -- layer=1 filter=181 channel=113
    -11, 19, -9, -4, 4, 15, 7, 12, 21,
    -- layer=1 filter=181 channel=114
    21, -31, 26, -10, 12, 3, 4, 7, 24,
    -- layer=1 filter=181 channel=115
    -32, 16, 15, -27, -6, 15, -14, -8, 20,
    -- layer=1 filter=181 channel=116
    1, 10, -11, -6, 0, 8, -7, 6, 10,
    -- layer=1 filter=181 channel=117
    -19, -19, 12, -54, -35, -4, 6, -23, 7,
    -- layer=1 filter=181 channel=118
    9, 0, 2, 22, -26, -5, 3, -4, -23,
    -- layer=1 filter=181 channel=119
    27, 41, -94, 31, 80, -75, 17, 84, -38,
    -- layer=1 filter=181 channel=120
    -5, -8, -10, -14, -10, 14, -9, -3, 2,
    -- layer=1 filter=181 channel=121
    -14, 7, 29, -26, 1, 15, 6, -13, 19,
    -- layer=1 filter=181 channel=122
    -2, 1, 9, -10, 3, 3, -8, 9, 9,
    -- layer=1 filter=181 channel=123
    0, 24, 28, -33, 0, 12, -13, -13, 20,
    -- layer=1 filter=181 channel=124
    9, 1, 16, 14, 0, 26, 13, 12, 3,
    -- layer=1 filter=181 channel=125
    -9, -2, 15, -25, 2, 29, 0, 15, 23,
    -- layer=1 filter=181 channel=126
    -8, -66, -23, -15, -38, 0, -47, -5, -26,
    -- layer=1 filter=181 channel=127
    1, 7, 5, 14, -24, -2, 17, -6, 5,
    -- layer=1 filter=182 channel=0
    5, -4, 3, 4, -2, -1, -7, -2, -12,
    -- layer=1 filter=182 channel=1
    5, -4, 6, 4, 6, -9, -4, -2, -5,
    -- layer=1 filter=182 channel=2
    2, 3, -4, 7, 1, -5, 3, 7, -6,
    -- layer=1 filter=182 channel=3
    2, 2, 8, -10, 8, -7, 3, -5, 0,
    -- layer=1 filter=182 channel=4
    0, 0, 1, -10, -4, -11, -5, 1, 0,
    -- layer=1 filter=182 channel=5
    -9, 5, 6, 0, -5, -10, 2, -10, 1,
    -- layer=1 filter=182 channel=6
    1, -10, 2, -4, -1, 5, -3, -9, -13,
    -- layer=1 filter=182 channel=7
    0, 9, 1, 2, 7, -10, 1, -12, 6,
    -- layer=1 filter=182 channel=8
    1, -4, 1, -7, 7, -7, -4, 6, 5,
    -- layer=1 filter=182 channel=9
    9, 9, 0, 7, -3, -7, -12, 8, 7,
    -- layer=1 filter=182 channel=10
    5, 7, 2, -9, 0, -3, -1, 0, 11,
    -- layer=1 filter=182 channel=11
    -8, -9, 5, 6, 5, 0, 0, 4, 2,
    -- layer=1 filter=182 channel=12
    -10, 0, -10, 4, 8, 3, -5, -7, -5,
    -- layer=1 filter=182 channel=13
    0, -9, 6, 4, -13, -2, -14, -9, -8,
    -- layer=1 filter=182 channel=14
    -2, -6, 2, -8, 8, 6, 7, -8, -2,
    -- layer=1 filter=182 channel=15
    -1, 0, -4, -9, -1, -8, -8, 5, -3,
    -- layer=1 filter=182 channel=16
    8, 4, -6, 7, -3, -4, 3, -3, 5,
    -- layer=1 filter=182 channel=17
    3, 0, 1, 0, -13, 3, 7, -11, -11,
    -- layer=1 filter=182 channel=18
    -6, -4, 4, -10, 3, -6, 0, 6, 7,
    -- layer=1 filter=182 channel=19
    0, 1, -9, 0, -3, -5, -4, 0, -5,
    -- layer=1 filter=182 channel=20
    0, 6, -1, -6, 2, 1, 3, 6, -11,
    -- layer=1 filter=182 channel=21
    -9, 6, -7, -11, 8, -6, -10, -9, -6,
    -- layer=1 filter=182 channel=22
    -5, 0, -7, -8, 7, -9, 6, -1, -2,
    -- layer=1 filter=182 channel=23
    -2, -10, -4, 4, -6, -1, -8, 2, -8,
    -- layer=1 filter=182 channel=24
    1, -11, 3, 4, 0, -2, -12, 4, -9,
    -- layer=1 filter=182 channel=25
    -11, -3, -4, -9, 6, -8, 4, 0, 13,
    -- layer=1 filter=182 channel=26
    -7, -7, -7, -13, -11, 2, -9, -1, -7,
    -- layer=1 filter=182 channel=27
    -5, -10, 1, 2, 10, -8, 10, -9, -8,
    -- layer=1 filter=182 channel=28
    0, 7, -6, 8, -1, -11, -11, 0, 3,
    -- layer=1 filter=182 channel=29
    -12, 10, -6, 7, 8, -2, -4, -7, 12,
    -- layer=1 filter=182 channel=30
    2, -3, 3, -12, -6, 6, 0, -6, -3,
    -- layer=1 filter=182 channel=31
    -5, -2, -6, -11, 3, 4, -5, 0, -6,
    -- layer=1 filter=182 channel=32
    0, -2, -6, -1, -5, -6, -1, 6, -6,
    -- layer=1 filter=182 channel=33
    5, 4, 0, -10, 8, 3, -13, -6, -8,
    -- layer=1 filter=182 channel=34
    -1, -3, 2, -11, -11, -6, -11, -3, 4,
    -- layer=1 filter=182 channel=35
    8, 8, -2, -1, -9, -1, -2, -12, 0,
    -- layer=1 filter=182 channel=36
    -7, -8, 0, 6, 1, 0, -6, -11, -6,
    -- layer=1 filter=182 channel=37
    -4, 4, -8, 1, 2, -11, -3, -9, 6,
    -- layer=1 filter=182 channel=38
    -12, -12, -4, -10, 1, 9, -1, -4, -9,
    -- layer=1 filter=182 channel=39
    -3, -10, -7, 4, -10, -6, -5, 2, -9,
    -- layer=1 filter=182 channel=40
    -9, 7, -1, 5, 0, -6, 2, 2, -4,
    -- layer=1 filter=182 channel=41
    1, 0, 7, 8, 7, -3, 2, -6, -5,
    -- layer=1 filter=182 channel=42
    6, 3, 6, 2, -1, 8, -3, 4, -10,
    -- layer=1 filter=182 channel=43
    2, 0, -7, 3, 0, 0, -12, -10, -8,
    -- layer=1 filter=182 channel=44
    6, 1, -1, 0, 3, 3, 4, 2, 3,
    -- layer=1 filter=182 channel=45
    -9, -8, -11, -6, -2, -11, -8, 2, -6,
    -- layer=1 filter=182 channel=46
    8, 5, -2, -5, -6, 12, -12, -6, 11,
    -- layer=1 filter=182 channel=47
    -11, -3, 5, -2, -9, 2, 7, -7, -8,
    -- layer=1 filter=182 channel=48
    -3, 0, 3, 0, 7, 3, -8, 5, 0,
    -- layer=1 filter=182 channel=49
    2, 4, 7, -5, 0, -9, -6, -5, -3,
    -- layer=1 filter=182 channel=50
    -11, 7, -10, 6, 7, -8, -10, 8, 1,
    -- layer=1 filter=182 channel=51
    6, 0, -15, 1, 0, 8, -15, -11, -3,
    -- layer=1 filter=182 channel=52
    -8, 0, 8, 7, 6, -4, -9, 6, 5,
    -- layer=1 filter=182 channel=53
    7, 5, 7, -1, -7, 3, -1, -4, -7,
    -- layer=1 filter=182 channel=54
    7, -3, 4, 6, 8, -6, 5, -13, 12,
    -- layer=1 filter=182 channel=55
    -4, -4, 9, 4, -15, -11, -7, -9, -6,
    -- layer=1 filter=182 channel=56
    0, -7, 7, -8, 6, -1, 0, -4, -3,
    -- layer=1 filter=182 channel=57
    0, -5, 1, -4, 1, 7, 7, -1, 2,
    -- layer=1 filter=182 channel=58
    -12, -1, -9, 6, -6, -8, 1, -7, -3,
    -- layer=1 filter=182 channel=59
    7, 1, 1, 7, 7, -5, -3, 6, -11,
    -- layer=1 filter=182 channel=60
    0, 9, -4, 9, 1, -8, -6, 2, 7,
    -- layer=1 filter=182 channel=61
    5, -1, 4, 3, -8, 1, -9, -2, 1,
    -- layer=1 filter=182 channel=62
    7, 0, -11, 5, 6, 0, -6, -5, -12,
    -- layer=1 filter=182 channel=63
    6, -8, 8, -3, -4, 7, -9, -5, -3,
    -- layer=1 filter=182 channel=64
    3, -8, 4, -2, -8, -5, 6, 7, 5,
    -- layer=1 filter=182 channel=65
    -9, 6, 0, -1, 0, 0, -10, 0, -7,
    -- layer=1 filter=182 channel=66
    -3, -6, -9, -4, -1, -8, 8, 0, 5,
    -- layer=1 filter=182 channel=67
    -11, 8, -11, 5, -7, 2, -9, -2, 9,
    -- layer=1 filter=182 channel=68
    7, 0, -5, 0, -12, 2, -2, 4, 4,
    -- layer=1 filter=182 channel=69
    6, 10, 8, -8, 4, 8, -3, -9, -12,
    -- layer=1 filter=182 channel=70
    0, -10, 4, 5, 0, 3, -5, 7, -1,
    -- layer=1 filter=182 channel=71
    -7, -7, -18, 4, 2, 4, -13, 0, 7,
    -- layer=1 filter=182 channel=72
    8, 2, -6, -4, 1, -10, -11, 0, 7,
    -- layer=1 filter=182 channel=73
    3, 0, -9, 1, -7, -4, -9, 6, 0,
    -- layer=1 filter=182 channel=74
    -11, -1, 7, -6, -7, -10, 5, -8, -3,
    -- layer=1 filter=182 channel=75
    5, 4, -12, 0, 3, 7, 3, 1, 10,
    -- layer=1 filter=182 channel=76
    0, 5, 8, 0, -9, 1, -7, -4, -10,
    -- layer=1 filter=182 channel=77
    -2, -6, -11, -1, -9, -7, 4, 0, 0,
    -- layer=1 filter=182 channel=78
    -2, -9, -2, -1, -1, -2, -11, 0, 8,
    -- layer=1 filter=182 channel=79
    -9, 0, 0, -8, -7, -7, 0, -7, 2,
    -- layer=1 filter=182 channel=80
    -2, -4, -4, 0, -10, -9, 4, 4, -3,
    -- layer=1 filter=182 channel=81
    6, -2, -8, -10, -7, 3, 5, -4, 0,
    -- layer=1 filter=182 channel=82
    9, -4, -3, -5, 7, 2, -8, 1, 3,
    -- layer=1 filter=182 channel=83
    7, 7, -4, 0, -11, 0, -11, -2, 3,
    -- layer=1 filter=182 channel=84
    -11, 1, 5, -16, 0, -5, 3, -5, -3,
    -- layer=1 filter=182 channel=85
    -3, 0, 2, 7, 3, -1, 2, 8, -7,
    -- layer=1 filter=182 channel=86
    1, -9, -7, -4, 7, -2, -2, -3, 3,
    -- layer=1 filter=182 channel=87
    -9, -7, -2, -11, 0, -10, -2, -11, -1,
    -- layer=1 filter=182 channel=88
    0, -5, 1, -12, -6, -7, -1, 0, 1,
    -- layer=1 filter=182 channel=89
    1, -17, 0, -5, 7, -13, -10, 0, -12,
    -- layer=1 filter=182 channel=90
    -8, -7, -10, 3, 1, -10, -3, -11, 1,
    -- layer=1 filter=182 channel=91
    0, -8, -2, -8, 5, -5, -9, 0, -1,
    -- layer=1 filter=182 channel=92
    -6, -5, -10, 3, 6, 5, -4, -1, 8,
    -- layer=1 filter=182 channel=93
    3, 1, -5, 3, 0, 3, 3, 0, 0,
    -- layer=1 filter=182 channel=94
    6, 0, -6, 0, -1, -9, 0, 0, 2,
    -- layer=1 filter=182 channel=95
    4, 4, 4, -12, -5, -14, -5, 3, -2,
    -- layer=1 filter=182 channel=96
    -9, -6, 4, 8, 7, 5, -8, -4, 5,
    -- layer=1 filter=182 channel=97
    -7, -7, 5, 0, 3, 0, -10, 3, 5,
    -- layer=1 filter=182 channel=98
    -3, 0, -5, -5, -1, 3, 8, 2, 0,
    -- layer=1 filter=182 channel=99
    -6, 6, -8, 2, -6, 4, -9, 0, -3,
    -- layer=1 filter=182 channel=100
    2, -11, -4, 5, 3, 0, -1, 0, 8,
    -- layer=1 filter=182 channel=101
    -10, -8, -3, 4, 8, -2, 0, 7, -1,
    -- layer=1 filter=182 channel=102
    -3, 1, -3, 5, -5, 6, -4, 0, 3,
    -- layer=1 filter=182 channel=103
    -11, -2, -6, 1, 7, -7, -10, 5, -8,
    -- layer=1 filter=182 channel=104
    4, -2, -9, 0, 0, -3, 3, -7, 1,
    -- layer=1 filter=182 channel=105
    -2, 3, 0, -1, -11, -1, 1, 0, -11,
    -- layer=1 filter=182 channel=106
    -11, -9, 8, -6, -8, -9, 0, -4, -7,
    -- layer=1 filter=182 channel=107
    8, -3, 5, 4, -3, -10, -7, -7, 9,
    -- layer=1 filter=182 channel=108
    -6, -1, 0, -3, -6, -2, -14, -3, -17,
    -- layer=1 filter=182 channel=109
    6, -6, 11, -1, 6, 8, -5, -9, -10,
    -- layer=1 filter=182 channel=110
    -7, -11, -11, -1, -6, 2, -4, -2, -8,
    -- layer=1 filter=182 channel=111
    -4, -4, -9, 0, -3, -8, -9, 0, -6,
    -- layer=1 filter=182 channel=112
    -11, -1, -9, 0, -5, 7, -6, -9, 4,
    -- layer=1 filter=182 channel=113
    -11, -8, 5, -5, -3, -10, -8, -4, -6,
    -- layer=1 filter=182 channel=114
    10, -7, 4, 8, 1, 0, -3, 8, -2,
    -- layer=1 filter=182 channel=115
    1, -7, 5, -10, 0, -9, 1, 0, -9,
    -- layer=1 filter=182 channel=116
    1, -6, -3, -2, -4, -6, 1, -4, -8,
    -- layer=1 filter=182 channel=117
    0, 4, -11, -3, 5, 6, 8, 3, 4,
    -- layer=1 filter=182 channel=118
    2, -12, -12, 3, -10, -1, 2, -1, -2,
    -- layer=1 filter=182 channel=119
    -5, -5, -3, -4, -5, -4, 8, -9, 4,
    -- layer=1 filter=182 channel=120
    1, -3, -9, -2, -7, -2, -3, -17, 1,
    -- layer=1 filter=182 channel=121
    -10, 1, -8, -4, -8, -2, -13, 1, 0,
    -- layer=1 filter=182 channel=122
    5, -2, -2, -7, 3, 1, -10, -8, 2,
    -- layer=1 filter=182 channel=123
    3, -2, 4, 6, 0, 0, -6, -8, 1,
    -- layer=1 filter=182 channel=124
    -4, -2, 8, 2, -11, 1, 4, -3, -6,
    -- layer=1 filter=182 channel=125
    -7, 0, 5, -1, -4, -5, -2, 4, 10,
    -- layer=1 filter=182 channel=126
    -9, 0, 6, -1, -8, 2, -7, 3, 0,
    -- layer=1 filter=182 channel=127
    -9, -3, -2, -8, -9, 4, -4, -2, -4,
    -- layer=1 filter=183 channel=0
    -11, -7, 2, -10, -9, 2, 5, -11, 0,
    -- layer=1 filter=183 channel=1
    7, 8, 23, 19, -17, -32, -7, -15, -34,
    -- layer=1 filter=183 channel=2
    51, 18, 29, 20, 16, 14, 1, -1, 3,
    -- layer=1 filter=183 channel=3
    -6, 8, -4, 1, -12, -7, -7, 2, 3,
    -- layer=1 filter=183 channel=4
    -6, -2, 6, 2, 1, 0, 2, -3, -11,
    -- layer=1 filter=183 channel=5
    -13, 6, 21, 42, -43, -62, -48, -73, -82,
    -- layer=1 filter=183 channel=6
    0, 3, 24, -8, -12, 13, -10, -14, -7,
    -- layer=1 filter=183 channel=7
    18, -11, -15, 5, -72, -82, -22, -88, -68,
    -- layer=1 filter=183 channel=8
    0, 17, 11, 23, -68, -108, -73, -104, -125,
    -- layer=1 filter=183 channel=9
    3, 7, 4, -23, 0, -16, -24, -25, -14,
    -- layer=1 filter=183 channel=10
    25, 7, -24, 16, -67, -66, -13, -82, -48,
    -- layer=1 filter=183 channel=11
    6, 23, 7, -3, 11, 15, 16, 1, 15,
    -- layer=1 filter=183 channel=12
    -20, -27, 0, -30, -20, -32, 9, -98, -83,
    -- layer=1 filter=183 channel=13
    -4, 4, 26, 5, -11, 24, 1, -3, 0,
    -- layer=1 filter=183 channel=14
    -26, -22, 0, 15, -51, -32, -31, -36, -67,
    -- layer=1 filter=183 channel=15
    39, 32, 44, 9, -10, -17, -30, -13, -26,
    -- layer=1 filter=183 channel=16
    -8, 7, 10, 31, -51, -94, -56, -79, -82,
    -- layer=1 filter=183 channel=17
    -8, 14, 21, -8, -1, 0, 3, 12, 17,
    -- layer=1 filter=183 channel=18
    3, -15, 5, -33, -25, -41, -13, -28, -58,
    -- layer=1 filter=183 channel=19
    -3, -33, -33, -73, -119, -99, -118, -131, -173,
    -- layer=1 filter=183 channel=20
    6, 10, 22, 18, 12, 24, 11, 22, 15,
    -- layer=1 filter=183 channel=21
    26, 15, 29, 18, 18, 19, 10, 4, 17,
    -- layer=1 filter=183 channel=22
    10, 30, 27, 18, 0, 14, 17, 11, 7,
    -- layer=1 filter=183 channel=23
    9, -32, -17, -3, -40, -21, -23, 1, -35,
    -- layer=1 filter=183 channel=24
    15, 20, 41, 27, 8, 16, 41, 21, 30,
    -- layer=1 filter=183 channel=25
    46, 15, 0, 33, -51, -87, -30, -94, -52,
    -- layer=1 filter=183 channel=26
    -17, -2, 41, -13, -30, 11, 25, -7, -15,
    -- layer=1 filter=183 channel=27
    -14, -4, 3, 4, 12, 13, 28, 17, 12,
    -- layer=1 filter=183 channel=28
    -10, 11, 7, 47, -34, -34, -4, -34, -18,
    -- layer=1 filter=183 channel=29
    -6, 12, 11, -1, 12, 0, 2, 4, 15,
    -- layer=1 filter=183 channel=30
    -53, -45, -60, -87, -97, -73, -76, -132, -155,
    -- layer=1 filter=183 channel=31
    7, -10, 3, 15, 16, 28, 49, 9, 12,
    -- layer=1 filter=183 channel=32
    -75, -105, -10, -72, -81, -84, -46, -47, -66,
    -- layer=1 filter=183 channel=33
    -8, 0, -4, 1, 8, 15, 0, 12, 0,
    -- layer=1 filter=183 channel=34
    29, 12, 15, 22, 21, 20, 2, 0, 18,
    -- layer=1 filter=183 channel=35
    -1, -13, -12, -17, -16, -10, -1, 0, -18,
    -- layer=1 filter=183 channel=36
    21, 10, 21, 0, 6, 10, 16, 24, 13,
    -- layer=1 filter=183 channel=37
    0, 20, 1, 8, -68, -102, -72, -117, -107,
    -- layer=1 filter=183 channel=38
    19, 24, 28, 2, 16, 12, 12, 13, 14,
    -- layer=1 filter=183 channel=39
    -10, -1, 4, -14, -3, 2, 5, 0, -8,
    -- layer=1 filter=183 channel=40
    2, -6, 25, -13, 3, 20, 23, 1, 5,
    -- layer=1 filter=183 channel=41
    -8, -49, 10, -10, -23, -68, 2, -49, -51,
    -- layer=1 filter=183 channel=42
    38, -5, 7, 8, -6, -1, 17, -11, -27,
    -- layer=1 filter=183 channel=43
    4, 2, 8, 45, -31, -55, -10, -49, -45,
    -- layer=1 filter=183 channel=44
    -54, -60, 4, -65, -84, -47, -35, -60, -67,
    -- layer=1 filter=183 channel=45
    3, 27, 36, -3, -6, 11, 6, -5, 5,
    -- layer=1 filter=183 channel=46
    -8, 25, 15, -47, -59, -47, -102, -95, -89,
    -- layer=1 filter=183 channel=47
    -4, -35, -32, 5, -24, -45, -5, -8, -53,
    -- layer=1 filter=183 channel=48
    4, 0, -4, 5, -1, -4, 2, -1, -3,
    -- layer=1 filter=183 channel=49
    18, 10, -3, -5, 6, -8, -25, -9, -1,
    -- layer=1 filter=183 channel=50
    3, -7, 1, 17, -4, -2, 20, 14, 14,
    -- layer=1 filter=183 channel=51
    21, 12, 24, 3, 14, 14, 9, -8, 1,
    -- layer=1 filter=183 channel=52
    1, -2, 1, 5, -3, 1, 7, -11, -14,
    -- layer=1 filter=183 channel=53
    17, 10, 16, 2, 0, 5, 18, 11, 6,
    -- layer=1 filter=183 channel=54
    69, 23, 0, 36, -45, -56, -35, -55, -54,
    -- layer=1 filter=183 channel=55
    10, 9, 29, 9, 27, 19, 23, 21, 21,
    -- layer=1 filter=183 channel=56
    -2, -10, 7, -1, -8, 6, -1, -4, -4,
    -- layer=1 filter=183 channel=57
    49, 19, 18, 29, -14, 8, 29, -21, 0,
    -- layer=1 filter=183 channel=58
    29, -62, -47, -56, -136, -104, -63, -41, -82,
    -- layer=1 filter=183 channel=59
    -6, -9, -12, 8, -5, 3, -12, -13, -3,
    -- layer=1 filter=183 channel=60
    0, 15, 3, 3, 10, 10, -4, 12, -3,
    -- layer=1 filter=183 channel=61
    -5, -14, 0, -4, -2, -11, -14, -1, -13,
    -- layer=1 filter=183 channel=62
    -11, -1, -2, 0, -82, -103, -76, -108, -98,
    -- layer=1 filter=183 channel=63
    13, 14, 4, -9, 2, 5, 9, 0, 8,
    -- layer=1 filter=183 channel=64
    3, 10, -3, -15, -4, -8, -4, 0, -2,
    -- layer=1 filter=183 channel=65
    -3, 0, 1, 3, 1, 1, 0, -10, 9,
    -- layer=1 filter=183 channel=66
    3, 4, -3, 4, 12, 8, 15, 8, 17,
    -- layer=1 filter=183 channel=67
    29, 17, 14, -18, -7, -2, -16, -35, -8,
    -- layer=1 filter=183 channel=68
    -74, -97, 18, -88, -148, -68, -56, -127, -92,
    -- layer=1 filter=183 channel=69
    0, 1, 46, -11, -59, -48, -34, -31, -69,
    -- layer=1 filter=183 channel=70
    18, 11, 7, 10, 13, 20, 14, -1, 3,
    -- layer=1 filter=183 channel=71
    26, 29, 12, 38, 31, 20, 33, 22, 37,
    -- layer=1 filter=183 channel=72
    -19, -29, -26, -68, -53, -45, -68, -86, -94,
    -- layer=1 filter=183 channel=73
    -1, 9, -4, -1, -8, -5, 13, -7, 6,
    -- layer=1 filter=183 channel=74
    -47, -29, -12, -37, -36, -27, -16, -40, -55,
    -- layer=1 filter=183 channel=75
    6, -9, 3, -34, -46, -53, -29, -89, -100,
    -- layer=1 filter=183 channel=76
    -9, -11, 10, 1, -15, -4, 1, -3, -19,
    -- layer=1 filter=183 channel=77
    10, 10, 17, 11, 10, 15, 4, 5, 1,
    -- layer=1 filter=183 channel=78
    -5, -9, 5, 7, -15, 0, 3, -10, -14,
    -- layer=1 filter=183 channel=79
    15, 13, 31, 5, -62, -78, -31, -51, -70,
    -- layer=1 filter=183 channel=80
    -2, 2, -6, -14, 6, -9, 3, 1, -4,
    -- layer=1 filter=183 channel=81
    16, 13, 7, 25, 22, 11, 26, 33, 26,
    -- layer=1 filter=183 channel=82
    25, 12, 21, 20, 1, 10, 11, 5, 5,
    -- layer=1 filter=183 channel=83
    -19, -2, 16, -25, -36, -26, -28, -18, -26,
    -- layer=1 filter=183 channel=84
    -112, -105, -93, -150, -106, -138, -116, -145, -136,
    -- layer=1 filter=183 channel=85
    48, -23, -10, -25, -67, -42, -25, 1, 0,
    -- layer=1 filter=183 channel=86
    6, 25, 14, 21, 27, 15, 23, 22, 32,
    -- layer=1 filter=183 channel=87
    -11, 6, 0, -74, -42, -52, -27, -81, -81,
    -- layer=1 filter=183 channel=88
    16, 9, 12, 8, 7, 18, 1, 13, 4,
    -- layer=1 filter=183 channel=89
    0, 11, 1, 4, 4, 15, 3, 5, 11,
    -- layer=1 filter=183 channel=90
    -76, -59, 28, -88, -148, -49, -59, -115, -91,
    -- layer=1 filter=183 channel=91
    26, 23, 15, 17, 7, 16, 6, 9, 8,
    -- layer=1 filter=183 channel=92
    7, -27, 3, 12, -8, -54, -29, -6, -59,
    -- layer=1 filter=183 channel=93
    11, 21, 21, 26, 17, 24, 27, 26, 28,
    -- layer=1 filter=183 channel=94
    -3, 13, -5, -14, 10, 2, 6, -9, 10,
    -- layer=1 filter=183 channel=95
    -72, -83, -83, -110, -110, -104, -116, -154, -140,
    -- layer=1 filter=183 channel=96
    -12, 0, -3, -12, -3, -2, -1, -6, -7,
    -- layer=1 filter=183 channel=97
    1, 14, 5, 21, 8, 0, 19, 16, 23,
    -- layer=1 filter=183 channel=98
    17, 34, 29, 18, -40, -52, -17, -60, -48,
    -- layer=1 filter=183 channel=99
    -44, -5, -26, 1, -50, -25, -10, -26, -31,
    -- layer=1 filter=183 channel=100
    2, -6, 1, -7, 3, -18, 3, -2, -13,
    -- layer=1 filter=183 channel=101
    14, 26, 14, 2, 19, 15, -1, 9, 13,
    -- layer=1 filter=183 channel=102
    -22, 8, 6, -5, -14, -11, -20, -9, -3,
    -- layer=1 filter=183 channel=103
    16, 9, 7, -10, 2, 6, 23, 0, -4,
    -- layer=1 filter=183 channel=104
    27, -6, -4, -2, -4, -18, -3, 2, -12,
    -- layer=1 filter=183 channel=105
    0, 13, 10, 5, 17, 1, 7, 19, 14,
    -- layer=1 filter=183 channel=106
    9, 2, 34, 5, 15, 17, 9, 2, -2,
    -- layer=1 filter=183 channel=107
    1, 9, 4, 17, 1, 2, 6, 13, -2,
    -- layer=1 filter=183 channel=108
    -63, -72, 19, -100, -128, -87, -54, -79, -83,
    -- layer=1 filter=183 channel=109
    -7, 0, -8, -3, 8, 5, 0, -9, 2,
    -- layer=1 filter=183 channel=110
    -14, -8, 6, -10, 9, -3, -3, -11, 5,
    -- layer=1 filter=183 channel=111
    -43, -43, -33, -90, -90, -83, -78, -98, -129,
    -- layer=1 filter=183 channel=112
    -42, -49, -26, -66, -61, -77, -80, -83, -93,
    -- layer=1 filter=183 channel=113
    49, 29, 29, 21, 17, 27, 22, 12, 35,
    -- layer=1 filter=183 channel=114
    8, -3, 14, 27, 0, -11, -26, -8, -21,
    -- layer=1 filter=183 channel=115
    24, 12, 18, 30, 24, 24, 17, 17, 33,
    -- layer=1 filter=183 channel=116
    1, 10, 1, -7, -5, -5, -1, 0, -2,
    -- layer=1 filter=183 channel=117
    -63, -102, -62, -145, -132, -120, -90, -103, -137,
    -- layer=1 filter=183 channel=118
    -77, -66, -52, -100, -80, -93, -68, -109, -117,
    -- layer=1 filter=183 channel=119
    -58, -80, 24, -74, -103, -79, -56, -76, -82,
    -- layer=1 filter=183 channel=120
    29, 22, 25, 22, 9, 10, 3, 8, 4,
    -- layer=1 filter=183 channel=121
    -5, 11, -4, -16, -24, -18, 1, -27, -16,
    -- layer=1 filter=183 channel=122
    8, 2, 8, -2, 7, 0, -4, -6, -9,
    -- layer=1 filter=183 channel=123
    17, 14, 6, -7, 10, 1, 6, 1, 10,
    -- layer=1 filter=183 channel=124
    -13, -6, 8, 0, -1, 0, -9, 5, 8,
    -- layer=1 filter=183 channel=125
    4, -3, 10, -5, -15, 7, -8, -36, 4,
    -- layer=1 filter=183 channel=126
    -17, 25, 4, -14, -73, -88, -52, -73, -85,
    -- layer=1 filter=183 channel=127
    -111, -81, -83, -120, -101, -124, -108, -155, -160,
    -- layer=1 filter=184 channel=0
    4, 1, 1, -8, -13, -6, -6, 1, 4,
    -- layer=1 filter=184 channel=1
    -6, -6, 2, 5, -11, 2, -3, -2, -10,
    -- layer=1 filter=184 channel=2
    7, 6, -8, 0, 5, -9, 6, -9, -11,
    -- layer=1 filter=184 channel=3
    3, -10, -4, -4, 3, -2, 6, 9, 7,
    -- layer=1 filter=184 channel=4
    3, -7, -9, -5, -10, -7, 8, -2, -8,
    -- layer=1 filter=184 channel=5
    -5, 1, -1, -1, -5, -7, -11, -13, -17,
    -- layer=1 filter=184 channel=6
    8, 0, 0, 3, -4, 8, -3, -1, 12,
    -- layer=1 filter=184 channel=7
    5, 0, -3, -15, -11, -8, 3, 1, -10,
    -- layer=1 filter=184 channel=8
    3, -1, 0, -8, 0, 3, -7, -5, 1,
    -- layer=1 filter=184 channel=9
    -3, -3, -4, -13, 3, 0, -13, -4, 0,
    -- layer=1 filter=184 channel=10
    3, 0, -18, 0, -3, -11, -15, 6, 7,
    -- layer=1 filter=184 channel=11
    2, -14, -8, -11, -10, -10, -12, -13, -4,
    -- layer=1 filter=184 channel=12
    6, -7, 4, 1, 7, 4, 9, -3, -9,
    -- layer=1 filter=184 channel=13
    -3, 7, 0, -1, 4, -7, -3, 2, 7,
    -- layer=1 filter=184 channel=14
    -16, -12, -8, 1, -15, -2, -8, -10, -6,
    -- layer=1 filter=184 channel=15
    -6, -1, -5, -9, -12, -4, 5, -7, 2,
    -- layer=1 filter=184 channel=16
    -11, -2, 7, 3, -12, 8, 3, 2, -1,
    -- layer=1 filter=184 channel=17
    -1, 2, -12, 0, 7, -5, 5, -10, -8,
    -- layer=1 filter=184 channel=18
    -2, -12, 3, -7, -5, 4, 5, -3, 8,
    -- layer=1 filter=184 channel=19
    7, -10, -7, 3, -11, 4, -8, -2, -4,
    -- layer=1 filter=184 channel=20
    -8, 6, -11, 1, -6, -3, 1, 2, -10,
    -- layer=1 filter=184 channel=21
    -9, 4, 2, 0, -9, 2, -5, 1, -7,
    -- layer=1 filter=184 channel=22
    7, -1, 8, -1, 8, 3, 3, -12, 8,
    -- layer=1 filter=184 channel=23
    -4, 0, 0, -14, -5, 0, 0, -4, -10,
    -- layer=1 filter=184 channel=24
    5, 4, -3, -14, 0, -12, -8, -12, -7,
    -- layer=1 filter=184 channel=25
    -6, -3, -5, 0, 4, -3, -8, 1, -7,
    -- layer=1 filter=184 channel=26
    5, 7, -4, 2, -5, 1, 6, -6, -4,
    -- layer=1 filter=184 channel=27
    0, -2, 8, 8, 0, -11, 0, -9, 3,
    -- layer=1 filter=184 channel=28
    -7, -1, 5, 5, -14, 5, -1, -8, -7,
    -- layer=1 filter=184 channel=29
    1, 6, 4, -10, 0, 8, 0, -3, 8,
    -- layer=1 filter=184 channel=30
    -9, -12, -10, 7, 4, -11, 0, 3, -3,
    -- layer=1 filter=184 channel=31
    5, -8, -1, 6, 6, 3, -2, -6, 5,
    -- layer=1 filter=184 channel=32
    -3, 2, 3, 0, -7, -2, -13, 0, -2,
    -- layer=1 filter=184 channel=33
    0, 3, 8, 8, -4, -2, 11, -12, -4,
    -- layer=1 filter=184 channel=34
    -1, -6, -12, -11, 0, 3, -4, -4, 4,
    -- layer=1 filter=184 channel=35
    -8, -4, -4, 2, 3, 4, 8, -3, 6,
    -- layer=1 filter=184 channel=36
    6, 3, -5, -1, 3, 5, -6, -8, -1,
    -- layer=1 filter=184 channel=37
    0, -4, 6, 0, -8, 4, -1, 1, -11,
    -- layer=1 filter=184 channel=38
    -5, 3, 0, 0, -7, 7, 10, 2, 7,
    -- layer=1 filter=184 channel=39
    7, 6, -10, 6, -8, 2, -3, -6, -11,
    -- layer=1 filter=184 channel=40
    -9, -8, 4, 1, 8, -2, 0, 0, 12,
    -- layer=1 filter=184 channel=41
    0, -4, 4, 5, -7, 0, -11, 4, 6,
    -- layer=1 filter=184 channel=42
    -16, -11, -10, 0, 0, 3, -5, -11, -8,
    -- layer=1 filter=184 channel=43
    7, -8, 6, -9, 1, -13, -10, -3, -7,
    -- layer=1 filter=184 channel=44
    -4, -12, -2, -15, -6, -5, -9, -11, -10,
    -- layer=1 filter=184 channel=45
    0, -10, -12, -5, 4, 7, -3, -2, 7,
    -- layer=1 filter=184 channel=46
    6, -2, -2, -4, -12, 9, 2, 5, 8,
    -- layer=1 filter=184 channel=47
    -7, 4, -4, -6, 1, -2, -5, 3, 2,
    -- layer=1 filter=184 channel=48
    0, -1, 0, 6, -5, -2, -10, -4, 0,
    -- layer=1 filter=184 channel=49
    -2, 10, -9, 0, -4, 2, -9, -4, 0,
    -- layer=1 filter=184 channel=50
    -2, -5, -6, 2, -3, -12, 6, -9, -5,
    -- layer=1 filter=184 channel=51
    -4, 0, -13, -13, -2, -1, 0, 6, 0,
    -- layer=1 filter=184 channel=52
    -3, -6, 8, -7, -9, 10, 5, -5, 0,
    -- layer=1 filter=184 channel=53
    0, -1, -12, 8, 6, -1, 7, 0, 4,
    -- layer=1 filter=184 channel=54
    -1, -10, -7, -9, -2, 0, -14, -1, -10,
    -- layer=1 filter=184 channel=55
    3, 0, -7, -6, -13, 0, -14, -4, 0,
    -- layer=1 filter=184 channel=56
    4, 0, 0, -7, 0, -12, 7, -9, 8,
    -- layer=1 filter=184 channel=57
    6, -11, 3, -8, 3, 0, -10, -9, -5,
    -- layer=1 filter=184 channel=58
    0, 3, -3, 4, 5, -10, -13, 1, -1,
    -- layer=1 filter=184 channel=59
    -1, -10, -4, 6, -2, 7, 7, -6, 6,
    -- layer=1 filter=184 channel=60
    0, -8, -10, 5, 0, -4, -4, -3, -1,
    -- layer=1 filter=184 channel=61
    2, -1, -2, -3, -6, -5, -2, -6, 1,
    -- layer=1 filter=184 channel=62
    -5, 5, -13, 3, -8, -3, -1, -12, -5,
    -- layer=1 filter=184 channel=63
    2, 1, 1, -15, -8, -5, -2, 4, 1,
    -- layer=1 filter=184 channel=64
    -10, 2, -4, -6, -3, -3, 0, -6, 0,
    -- layer=1 filter=184 channel=65
    2, 0, 4, -13, 0, -3, -7, 1, 5,
    -- layer=1 filter=184 channel=66
    4, -3, 0, 3, 4, -15, -14, 0, -5,
    -- layer=1 filter=184 channel=67
    -8, 5, -2, -1, 9, 8, 4, 5, -10,
    -- layer=1 filter=184 channel=68
    0, -10, -10, -3, 3, 1, -6, 1, -1,
    -- layer=1 filter=184 channel=69
    -5, -8, 0, 3, -1, -8, 0, -11, -6,
    -- layer=1 filter=184 channel=70
    -3, 7, 8, 4, -1, 4, 11, -1, -2,
    -- layer=1 filter=184 channel=71
    -10, -7, 0, 6, 1, -12, -3, 3, -7,
    -- layer=1 filter=184 channel=72
    -9, -8, -3, -7, 2, -6, -12, -3, -15,
    -- layer=1 filter=184 channel=73
    0, 0, -3, 0, 5, 6, 4, 0, -10,
    -- layer=1 filter=184 channel=74
    -3, -1, 1, 1, -6, -10, 0, -13, -13,
    -- layer=1 filter=184 channel=75
    -10, 0, -11, -4, -1, -15, 0, -17, -4,
    -- layer=1 filter=184 channel=76
    -3, -1, -5, 5, -11, -6, -3, 0, -1,
    -- layer=1 filter=184 channel=77
    -10, 4, 6, -4, -13, -9, 0, -3, -13,
    -- layer=1 filter=184 channel=78
    -7, -10, -13, -2, 2, 0, -8, -4, -8,
    -- layer=1 filter=184 channel=79
    5, -4, -9, 9, -4, -7, 4, 8, -9,
    -- layer=1 filter=184 channel=80
    6, 3, -4, -6, -1, -2, 4, 7, 6,
    -- layer=1 filter=184 channel=81
    -10, -13, 8, -2, -1, 2, -9, -4, 6,
    -- layer=1 filter=184 channel=82
    3, -8, -8, -7, -7, 7, 1, -7, -4,
    -- layer=1 filter=184 channel=83
    -1, 3, -13, -12, -13, -5, 4, -8, 4,
    -- layer=1 filter=184 channel=84
    1, -4, 4, 0, -10, 2, -7, 4, 0,
    -- layer=1 filter=184 channel=85
    -15, -4, -13, 0, -6, -9, 1, -6, -7,
    -- layer=1 filter=184 channel=86
    -9, 3, -8, -1, 1, 2, 6, -10, 5,
    -- layer=1 filter=184 channel=87
    -10, -1, 3, 5, 5, -5, -1, -7, -6,
    -- layer=1 filter=184 channel=88
    -4, -10, 0, 4, 11, -5, -6, 0, 0,
    -- layer=1 filter=184 channel=89
    -6, -11, -3, -7, 1, -6, 6, -1, -7,
    -- layer=1 filter=184 channel=90
    -2, -9, 0, -10, 0, 4, -12, 3, -1,
    -- layer=1 filter=184 channel=91
    0, -7, 8, 8, 2, 9, 9, 0, -1,
    -- layer=1 filter=184 channel=92
    0, 2, 2, 4, 0, 1, 6, -4, 6,
    -- layer=1 filter=184 channel=93
    -1, -5, -13, -8, 2, 1, -7, -4, -3,
    -- layer=1 filter=184 channel=94
    -4, 1, 5, -10, -9, -4, -11, -9, -6,
    -- layer=1 filter=184 channel=95
    -13, -13, -2, -4, -2, -4, -4, -13, 2,
    -- layer=1 filter=184 channel=96
    1, 3, -1, -5, 4, -7, -10, -8, -4,
    -- layer=1 filter=184 channel=97
    -2, 4, -2, -13, -9, -3, -6, -9, 1,
    -- layer=1 filter=184 channel=98
    3, 10, 7, 7, -5, -1, -6, -9, 9,
    -- layer=1 filter=184 channel=99
    -1, 1, 5, -5, -7, -8, 0, 5, 4,
    -- layer=1 filter=184 channel=100
    2, -8, -6, -10, 6, 0, -9, 0, 5,
    -- layer=1 filter=184 channel=101
    -10, 1, -4, 6, 0, 5, 4, -12, 6,
    -- layer=1 filter=184 channel=102
    -1, -5, -15, -9, 3, -5, -1, -7, 5,
    -- layer=1 filter=184 channel=103
    -7, -12, -14, -14, -15, -10, -10, -5, -8,
    -- layer=1 filter=184 channel=104
    -7, -3, 4, 4, -6, -6, -5, -3, -3,
    -- layer=1 filter=184 channel=105
    -8, -6, -4, 1, -11, -4, -9, -5, -15,
    -- layer=1 filter=184 channel=106
    -6, -8, -9, -2, 4, -7, 4, -9, 8,
    -- layer=1 filter=184 channel=107
    -10, -2, 2, -10, 0, -4, -9, 0, 3,
    -- layer=1 filter=184 channel=108
    -5, -2, -12, 3, 6, -1, 0, -17, -16,
    -- layer=1 filter=184 channel=109
    3, 1, -4, 6, -2, 3, 4, -9, -3,
    -- layer=1 filter=184 channel=110
    3, -11, -4, -12, 1, -11, -3, -1, -9,
    -- layer=1 filter=184 channel=111
    2, -2, 0, -2, -2, -14, -6, -4, 6,
    -- layer=1 filter=184 channel=112
    6, -4, -2, 0, -13, -8, 4, -12, 1,
    -- layer=1 filter=184 channel=113
    3, 3, 8, -5, 4, -3, -8, -9, 0,
    -- layer=1 filter=184 channel=114
    0, -11, -2, 2, -2, 1, -10, 0, -13,
    -- layer=1 filter=184 channel=115
    -7, 1, -14, 0, -8, 0, 2, 2, -8,
    -- layer=1 filter=184 channel=116
    -9, 0, 1, 0, -4, -8, 4, 5, 6,
    -- layer=1 filter=184 channel=117
    -14, 0, -15, 0, -4, -2, -15, -2, -16,
    -- layer=1 filter=184 channel=118
    -5, -10, -2, -1, -5, -11, -8, -1, -8,
    -- layer=1 filter=184 channel=119
    -15, -12, -10, 0, -11, -5, -8, -2, -11,
    -- layer=1 filter=184 channel=120
    -3, 0, 3, 3, 2, 7, 4, -8, 12,
    -- layer=1 filter=184 channel=121
    0, -3, -18, -8, -11, -1, -10, -3, -11,
    -- layer=1 filter=184 channel=122
    -7, 0, 2, 10, -5, 10, -3, -5, 0,
    -- layer=1 filter=184 channel=123
    -4, -2, -14, 0, -4, -4, -10, 5, 0,
    -- layer=1 filter=184 channel=124
    -8, -5, -6, -2, 4, 9, 6, -8, -6,
    -- layer=1 filter=184 channel=125
    -7, -8, -1, -4, 4, -13, 7, 11, 10,
    -- layer=1 filter=184 channel=126
    -3, -13, -4, -13, 4, -15, -5, -4, 1,
    -- layer=1 filter=184 channel=127
    -3, 0, -11, 4, -10, -12, -13, 6, -1,
    -- layer=1 filter=185 channel=0
    -8, -2, -11, 2, -2, 0, -5, 5, 6,
    -- layer=1 filter=185 channel=1
    2, 5, 6, -10, -2, 4, -4, 0, -7,
    -- layer=1 filter=185 channel=2
    -8, 4, 0, 5, 8, -10, 9, -3, -14,
    -- layer=1 filter=185 channel=3
    6, 7, 6, 3, 7, 3, -1, 3, 5,
    -- layer=1 filter=185 channel=4
    8, -7, 0, -4, -5, 7, -7, 8, 0,
    -- layer=1 filter=185 channel=5
    -9, -11, 4, -1, 9, 7, -10, -3, 9,
    -- layer=1 filter=185 channel=6
    9, -1, -5, 3, 0, 5, -9, 7, -1,
    -- layer=1 filter=185 channel=7
    4, -5, -1, -13, 1, 3, -4, 3, 0,
    -- layer=1 filter=185 channel=8
    -3, 7, 7, 8, -1, 9, 0, 9, 2,
    -- layer=1 filter=185 channel=9
    2, 6, 5, 10, -6, 3, -4, -2, -1,
    -- layer=1 filter=185 channel=10
    -4, -10, 6, -8, -4, -1, -9, 0, -3,
    -- layer=1 filter=185 channel=11
    -8, -11, -10, 7, 7, -2, -10, -3, 0,
    -- layer=1 filter=185 channel=12
    -10, 3, -6, 0, -3, 4, 7, 9, -1,
    -- layer=1 filter=185 channel=13
    0, -9, -1, -2, -9, -11, -11, 1, 1,
    -- layer=1 filter=185 channel=14
    6, 9, 0, 6, 9, 4, -1, 8, 1,
    -- layer=1 filter=185 channel=15
    9, 4, 2, 2, 6, 8, -6, 0, -9,
    -- layer=1 filter=185 channel=16
    5, 6, -3, 7, 4, -7, 2, -8, -10,
    -- layer=1 filter=185 channel=17
    2, -3, 3, 5, -6, 4, -1, 3, -8,
    -- layer=1 filter=185 channel=18
    -4, 5, -5, -2, 2, -6, 7, -8, 0,
    -- layer=1 filter=185 channel=19
    3, 0, 1, -2, 0, 2, -11, 0, 0,
    -- layer=1 filter=185 channel=20
    -1, -8, 2, -1, -11, 0, 4, -4, -7,
    -- layer=1 filter=185 channel=21
    -6, 6, 3, 0, 4, 10, 8, 1, 0,
    -- layer=1 filter=185 channel=22
    1, -5, 0, 7, -7, -10, -4, 5, -9,
    -- layer=1 filter=185 channel=23
    5, -3, 6, -1, -11, -1, -8, 6, -4,
    -- layer=1 filter=185 channel=24
    -7, -2, -3, 2, 0, 0, -10, 7, -4,
    -- layer=1 filter=185 channel=25
    0, 8, 1, 3, 3, -3, -5, 11, -5,
    -- layer=1 filter=185 channel=26
    -9, 4, 1, -1, 1, 2, -8, -7, 1,
    -- layer=1 filter=185 channel=27
    -3, -10, 6, 0, 0, 2, -7, 2, 6,
    -- layer=1 filter=185 channel=28
    -4, -4, -10, -3, -9, 5, -11, 9, 3,
    -- layer=1 filter=185 channel=29
    -11, -6, 0, 10, -8, 7, 11, 4, 9,
    -- layer=1 filter=185 channel=30
    -1, -10, -8, -10, -8, 10, -3, -7, 5,
    -- layer=1 filter=185 channel=31
    0, 0, 8, 5, -4, -1, -7, -11, -4,
    -- layer=1 filter=185 channel=32
    5, -1, 4, 2, 5, -7, 2, 7, -10,
    -- layer=1 filter=185 channel=33
    -5, -8, -5, 8, 2, 0, -1, 0, 0,
    -- layer=1 filter=185 channel=34
    8, 1, 4, 2, -7, 1, -8, 0, -3,
    -- layer=1 filter=185 channel=35
    6, -4, 6, 0, 8, -6, -3, 5, -6,
    -- layer=1 filter=185 channel=36
    -1, -2, 0, -8, 5, 3, -11, 6, -6,
    -- layer=1 filter=185 channel=37
    -5, 4, 9, -5, -7, -7, -3, -10, -3,
    -- layer=1 filter=185 channel=38
    -5, -2, 2, 0, -11, -11, 8, -10, -7,
    -- layer=1 filter=185 channel=39
    8, -2, -3, 8, 0, 2, 0, 8, 9,
    -- layer=1 filter=185 channel=40
    -3, -3, -10, 8, -9, -5, 3, 4, -2,
    -- layer=1 filter=185 channel=41
    5, 0, -6, 0, -2, 7, 5, 9, 2,
    -- layer=1 filter=185 channel=42
    4, 6, -9, -9, 2, -2, -10, 2, 3,
    -- layer=1 filter=185 channel=43
    4, -12, -8, -3, 9, 6, 6, -1, -2,
    -- layer=1 filter=185 channel=44
    -11, 5, -5, -10, 2, -2, 5, 6, 1,
    -- layer=1 filter=185 channel=45
    -10, -9, 8, 2, -6, 3, 6, -8, 0,
    -- layer=1 filter=185 channel=46
    3, -1, -7, 3, -6, 4, -10, -10, 9,
    -- layer=1 filter=185 channel=47
    -5, 11, -5, -4, -9, -6, -1, -4, -5,
    -- layer=1 filter=185 channel=48
    3, -1, 6, 7, -3, 1, -4, -7, -1,
    -- layer=1 filter=185 channel=49
    -5, 1, -8, 8, -8, 4, 8, -5, -7,
    -- layer=1 filter=185 channel=50
    -5, 4, -2, -11, 1, -6, 8, 4, 0,
    -- layer=1 filter=185 channel=51
    6, 1, -9, -7, -10, 2, 1, 7, -4,
    -- layer=1 filter=185 channel=52
    2, 0, -9, -3, 4, -1, -7, -5, 6,
    -- layer=1 filter=185 channel=53
    -4, -8, 5, -5, -11, 5, -5, 6, -2,
    -- layer=1 filter=185 channel=54
    -6, -4, 2, 0, -1, -9, 9, -5, -9,
    -- layer=1 filter=185 channel=55
    -2, 0, -6, 7, -4, 1, 2, -3, -6,
    -- layer=1 filter=185 channel=56
    0, 0, 1, 4, 6, 4, 0, 0, -3,
    -- layer=1 filter=185 channel=57
    0, -9, -8, 8, -9, -11, 0, -6, 6,
    -- layer=1 filter=185 channel=58
    -3, 5, 0, 0, -5, -3, -10, 0, -2,
    -- layer=1 filter=185 channel=59
    4, 0, 4, -3, -5, -5, 5, 8, 6,
    -- layer=1 filter=185 channel=60
    5, 8, 3, 0, -8, -3, -10, 6, 0,
    -- layer=1 filter=185 channel=61
    -11, 0, -8, -1, 3, 2, -7, 8, 3,
    -- layer=1 filter=185 channel=62
    -5, 3, -10, -3, 11, 9, 7, 7, -1,
    -- layer=1 filter=185 channel=63
    6, 4, 0, 0, -1, -3, 5, 5, -2,
    -- layer=1 filter=185 channel=64
    1, -2, -3, 6, 6, -8, 0, 2, 2,
    -- layer=1 filter=185 channel=65
    -3, -3, 3, 4, -8, 6, -5, -11, -10,
    -- layer=1 filter=185 channel=66
    -4, 1, -9, -9, 0, 8, -1, -1, -5,
    -- layer=1 filter=185 channel=67
    -6, 6, 3, -8, 4, -3, -1, 2, -4,
    -- layer=1 filter=185 channel=68
    8, -3, 4, -6, -7, 1, -8, -4, -4,
    -- layer=1 filter=185 channel=69
    9, 2, -10, -5, -8, -9, 3, -9, 2,
    -- layer=1 filter=185 channel=70
    -3, 2, -8, -7, 2, -11, -6, 2, 0,
    -- layer=1 filter=185 channel=71
    -4, 1, -10, -3, 2, 9, 3, -10, 3,
    -- layer=1 filter=185 channel=72
    -7, -1, -6, -2, 0, 7, -11, 3, 3,
    -- layer=1 filter=185 channel=73
    -8, 5, -12, -5, 4, -6, 7, 0, 0,
    -- layer=1 filter=185 channel=74
    -10, 7, -6, -10, -3, 1, -3, 4, -7,
    -- layer=1 filter=185 channel=75
    -3, -8, -1, 3, -4, 7, -6, -5, -8,
    -- layer=1 filter=185 channel=76
    -9, -4, 4, -10, -2, 0, -8, 4, -9,
    -- layer=1 filter=185 channel=77
    -6, 4, 0, -9, -6, -4, 5, -6, 2,
    -- layer=1 filter=185 channel=78
    -11, -8, 7, 8, 1, 7, -7, -11, 6,
    -- layer=1 filter=185 channel=79
    0, 3, 0, -2, -5, -6, -3, 2, -5,
    -- layer=1 filter=185 channel=80
    -8, 3, -10, -5, 0, 9, 0, 9, -4,
    -- layer=1 filter=185 channel=81
    2, -11, 3, -6, -7, -7, -7, 4, 0,
    -- layer=1 filter=185 channel=82
    -8, 7, -7, 8, -6, -9, -7, -2, -8,
    -- layer=1 filter=185 channel=83
    -7, 4, -10, 0, 5, 3, -5, -1, -8,
    -- layer=1 filter=185 channel=84
    0, 1, -11, -3, -6, -5, -3, 4, 0,
    -- layer=1 filter=185 channel=85
    5, -11, 4, 5, 7, -9, 1, -8, -7,
    -- layer=1 filter=185 channel=86
    -7, 0, -3, 5, 5, -10, 5, -4, 0,
    -- layer=1 filter=185 channel=87
    -1, -2, -6, 3, 8, -11, 2, 2, -4,
    -- layer=1 filter=185 channel=88
    3, -6, -11, 7, -1, -12, -8, -5, 3,
    -- layer=1 filter=185 channel=89
    -2, -3, 0, 3, 1, -10, -7, -3, -9,
    -- layer=1 filter=185 channel=90
    5, -7, -2, -9, -2, 7, -9, -2, 8,
    -- layer=1 filter=185 channel=91
    -9, -7, 7, 8, -10, 5, 0, -8, 0,
    -- layer=1 filter=185 channel=92
    0, 0, -1, -5, -1, 0, 1, -2, 8,
    -- layer=1 filter=185 channel=93
    6, 6, 0, 5, -5, 3, 5, -1, 0,
    -- layer=1 filter=185 channel=94
    -2, -5, -9, -5, 2, 0, 8, 3, 0,
    -- layer=1 filter=185 channel=95
    0, -5, -7, -10, -6, -8, -10, 0, 4,
    -- layer=1 filter=185 channel=96
    -8, -8, -9, -5, 7, 0, -11, -4, -3,
    -- layer=1 filter=185 channel=97
    3, -2, -2, -3, -10, -10, -7, -11, -3,
    -- layer=1 filter=185 channel=98
    4, 6, 5, 4, -10, 11, -5, 8, -7,
    -- layer=1 filter=185 channel=99
    7, -10, -5, 3, -4, 3, -7, -7, -1,
    -- layer=1 filter=185 channel=100
    -11, 8, 1, 0, 0, -10, 4, -3, 0,
    -- layer=1 filter=185 channel=101
    -8, 7, -1, -1, -8, -3, -1, -10, -4,
    -- layer=1 filter=185 channel=102
    -3, -1, -4, -2, 4, 0, -6, 0, -3,
    -- layer=1 filter=185 channel=103
    8, -5, -4, 0, -5, 2, 3, 2, 5,
    -- layer=1 filter=185 channel=104
    -3, 7, -1, -5, -9, 4, -8, -3, -9,
    -- layer=1 filter=185 channel=105
    7, 1, -2, 6, -1, -10, 0, 1, -4,
    -- layer=1 filter=185 channel=106
    8, 1, -11, 8, -7, -4, 2, 4, -1,
    -- layer=1 filter=185 channel=107
    11, 9, 11, -1, -2, 9, -10, -2, -8,
    -- layer=1 filter=185 channel=108
    9, -7, 5, -5, -7, 0, -11, -14, 0,
    -- layer=1 filter=185 channel=109
    4, 7, -1, -9, 2, 6, 0, 0, -8,
    -- layer=1 filter=185 channel=110
    -3, 3, 0, -1, 8, -10, 0, -8, -11,
    -- layer=1 filter=185 channel=111
    6, -2, -4, 5, 0, -5, 4, -2, -11,
    -- layer=1 filter=185 channel=112
    5, 1, 4, 0, -7, 6, -2, -6, 3,
    -- layer=1 filter=185 channel=113
    4, -4, -1, -4, 0, -11, -8, 5, -3,
    -- layer=1 filter=185 channel=114
    1, -5, -3, -6, -1, 1, 1, 1, -9,
    -- layer=1 filter=185 channel=115
    -5, 8, -3, 5, -1, -10, 5, -7, 1,
    -- layer=1 filter=185 channel=116
    -2, -10, -1, -2, -8, 7, -5, 2, -5,
    -- layer=1 filter=185 channel=117
    -7, 6, -2, -5, 2, 0, 5, 0, -5,
    -- layer=1 filter=185 channel=118
    -7, -3, -3, 0, 2, -12, -2, 4, 8,
    -- layer=1 filter=185 channel=119
    -9, -11, 7, 5, 2, 9, -2, 4, -4,
    -- layer=1 filter=185 channel=120
    3, 4, -1, -8, 8, 0, 10, -7, -6,
    -- layer=1 filter=185 channel=121
    -11, -4, 2, -7, -4, -5, -4, 2, 2,
    -- layer=1 filter=185 channel=122
    10, 3, 4, -7, -3, 0, -5, 7, -1,
    -- layer=1 filter=185 channel=123
    -5, -5, -2, -4, -5, 4, -9, 1, 3,
    -- layer=1 filter=185 channel=124
    -5, 11, 0, 1, 10, -2, -8, -10, 4,
    -- layer=1 filter=185 channel=125
    -8, -8, 0, -6, 0, -8, 8, -6, -3,
    -- layer=1 filter=185 channel=126
    -3, -2, -5, -12, -4, 5, 8, 3, 7,
    -- layer=1 filter=185 channel=127
    8, 4, 8, -3, 2, 8, 1, -1, 0,
    -- layer=1 filter=186 channel=0
    -3, -5, -11, -2, 1, 7, -5, 0, -1,
    -- layer=1 filter=186 channel=1
    1, -5, 5, -11, -2, 0, 4, -10, 7,
    -- layer=1 filter=186 channel=2
    5, -5, -4, -7, -11, -9, 9, -11, -3,
    -- layer=1 filter=186 channel=3
    -1, -7, 5, 8, -10, -9, 10, 6, 5,
    -- layer=1 filter=186 channel=4
    -4, 7, 1, 4, -3, 1, 5, -5, -10,
    -- layer=1 filter=186 channel=5
    -6, -2, 2, 6, 3, -10, -12, -5, -9,
    -- layer=1 filter=186 channel=6
    -2, -7, -2, 0, 8, -3, -4, 0, 8,
    -- layer=1 filter=186 channel=7
    8, -2, -4, -9, -6, 8, 0, 11, -8,
    -- layer=1 filter=186 channel=8
    -8, -6, 4, 6, 1, -1, 0, -11, -10,
    -- layer=1 filter=186 channel=9
    6, -6, -6, -6, -4, -12, 0, 8, 2,
    -- layer=1 filter=186 channel=10
    -3, -2, -2, -2, -3, 2, 8, -6, -1,
    -- layer=1 filter=186 channel=11
    -9, -7, -3, -2, -7, -12, 8, 1, -3,
    -- layer=1 filter=186 channel=12
    0, -1, 5, 0, -4, -1, -4, 1, 5,
    -- layer=1 filter=186 channel=13
    4, -7, -10, 7, -4, -1, -5, -6, -2,
    -- layer=1 filter=186 channel=14
    4, 5, 1, -9, -4, -11, 10, -12, 3,
    -- layer=1 filter=186 channel=15
    8, -2, -3, -2, 4, -12, -2, 6, -12,
    -- layer=1 filter=186 channel=16
    2, 0, 4, 2, 6, -2, -6, 6, -9,
    -- layer=1 filter=186 channel=17
    -6, 0, -5, 7, -3, 7, -1, -9, -2,
    -- layer=1 filter=186 channel=18
    -2, -4, -9, -10, -4, 0, 6, -9, 1,
    -- layer=1 filter=186 channel=19
    -7, 2, 5, -9, 7, -1, -12, -4, -11,
    -- layer=1 filter=186 channel=20
    1, -9, 6, 5, -9, -2, -11, -4, 3,
    -- layer=1 filter=186 channel=21
    7, 8, -2, 3, 0, 1, -10, -8, -9,
    -- layer=1 filter=186 channel=22
    5, -4, 3, 0, 2, 1, -2, -1, -5,
    -- layer=1 filter=186 channel=23
    5, -7, 0, -11, -12, 6, -8, -3, -4,
    -- layer=1 filter=186 channel=24
    -7, 0, 1, -6, -6, -5, -12, -5, -5,
    -- layer=1 filter=186 channel=25
    8, 7, 8, 2, -7, 8, 2, 8, -4,
    -- layer=1 filter=186 channel=26
    2, 8, 5, -7, 2, 6, 3, -1, -9,
    -- layer=1 filter=186 channel=27
    0, -6, 6, 8, -8, -5, -12, 5, 0,
    -- layer=1 filter=186 channel=28
    4, 8, -8, 4, -8, -4, 7, 5, -3,
    -- layer=1 filter=186 channel=29
    -8, -1, 0, 7, 3, -4, -7, 2, -12,
    -- layer=1 filter=186 channel=30
    0, 1, 0, -2, -3, -6, 7, -1, -11,
    -- layer=1 filter=186 channel=31
    4, -8, -1, -1, -11, 0, 0, -6, 8,
    -- layer=1 filter=186 channel=32
    0, -6, -10, 6, 2, 6, -4, -4, -8,
    -- layer=1 filter=186 channel=33
    -2, -7, 10, 8, 3, -9, -7, -6, -4,
    -- layer=1 filter=186 channel=34
    -9, 0, -8, 5, -6, -10, -7, 0, 4,
    -- layer=1 filter=186 channel=35
    -1, 0, 7, 0, -8, 0, 0, -10, -5,
    -- layer=1 filter=186 channel=36
    -9, 7, -8, 7, -6, -4, 5, -12, 4,
    -- layer=1 filter=186 channel=37
    5, 2, -1, -3, 2, 9, -2, 3, -6,
    -- layer=1 filter=186 channel=38
    -2, -6, 5, 4, -4, -9, -5, -1, -7,
    -- layer=1 filter=186 channel=39
    -10, -2, -10, 4, -3, 6, 3, -8, 8,
    -- layer=1 filter=186 channel=40
    8, 0, 10, -7, 0, -8, -7, -7, -6,
    -- layer=1 filter=186 channel=41
    6, 1, 2, -9, 1, -7, -3, 6, 7,
    -- layer=1 filter=186 channel=42
    4, -5, -10, 2, 8, 5, -6, -1, 2,
    -- layer=1 filter=186 channel=43
    7, 5, -7, -5, 3, 4, -4, -2, 4,
    -- layer=1 filter=186 channel=44
    7, 6, 4, -12, -5, -3, 0, 4, -10,
    -- layer=1 filter=186 channel=45
    -5, -3, 1, 0, -10, 2, -1, 1, 5,
    -- layer=1 filter=186 channel=46
    0, 3, 2, -8, 7, 4, -4, -8, -5,
    -- layer=1 filter=186 channel=47
    2, -4, 0, 0, -11, 7, -1, -13, 6,
    -- layer=1 filter=186 channel=48
    3, 1, 7, 5, 2, 2, -11, -4, 5,
    -- layer=1 filter=186 channel=49
    4, -7, 6, -3, 5, 6, 4, -5, 4,
    -- layer=1 filter=186 channel=50
    -6, 3, 1, 6, 7, 2, -9, -10, -5,
    -- layer=1 filter=186 channel=51
    7, 1, -1, -12, -8, 1, 6, -5, -2,
    -- layer=1 filter=186 channel=52
    4, -6, 1, 4, 3, 2, 6, -1, -6,
    -- layer=1 filter=186 channel=53
    7, -12, 2, -2, -1, -10, 4, -11, 8,
    -- layer=1 filter=186 channel=54
    -10, 7, 4, -5, -6, -4, 0, -1, 8,
    -- layer=1 filter=186 channel=55
    -3, 1, -6, -10, -2, 3, -11, 0, 0,
    -- layer=1 filter=186 channel=56
    3, 7, -13, -12, -6, 6, 8, 5, 0,
    -- layer=1 filter=186 channel=57
    4, 0, 3, 2, 5, -1, -6, 3, -12,
    -- layer=1 filter=186 channel=58
    2, 6, -1, 2, -5, 5, 5, -3, 3,
    -- layer=1 filter=186 channel=59
    2, 4, 0, 4, 2, -1, -7, -7, 7,
    -- layer=1 filter=186 channel=60
    0, -2, 0, -3, 9, 6, -10, 1, -1,
    -- layer=1 filter=186 channel=61
    0, 5, -8, 3, -2, -2, -2, -5, -1,
    -- layer=1 filter=186 channel=62
    -6, 2, -9, 8, -7, 11, 1, -5, 1,
    -- layer=1 filter=186 channel=63
    2, -12, 4, 1, -9, 0, -8, 4, -6,
    -- layer=1 filter=186 channel=64
    -1, -5, 2, -2, -10, 2, -12, -4, 4,
    -- layer=1 filter=186 channel=65
    -7, -5, -2, 6, 0, 1, 6, 6, 4,
    -- layer=1 filter=186 channel=66
    2, -11, -5, -1, 6, -6, 0, -4, -2,
    -- layer=1 filter=186 channel=67
    -8, -6, 4, -10, 3, -8, 2, 1, 3,
    -- layer=1 filter=186 channel=68
    0, -6, -12, 2, 0, -9, -9, -3, -10,
    -- layer=1 filter=186 channel=69
    -3, 1, -7, -13, -8, 4, 5, 7, 0,
    -- layer=1 filter=186 channel=70
    -8, -10, 6, -7, -8, 6, 9, 1, -13,
    -- layer=1 filter=186 channel=71
    5, 0, -5, -10, -12, 1, -5, 6, -12,
    -- layer=1 filter=186 channel=72
    -2, 2, 3, 3, 6, -13, -5, -3, 0,
    -- layer=1 filter=186 channel=73
    -9, -10, -3, -7, -12, 5, 0, -10, 0,
    -- layer=1 filter=186 channel=74
    0, -5, -11, 6, -4, 3, -11, 8, 0,
    -- layer=1 filter=186 channel=75
    -4, -7, 6, -1, 7, 6, 8, -11, 2,
    -- layer=1 filter=186 channel=76
    -12, -6, -12, -3, 8, 6, -6, -3, -7,
    -- layer=1 filter=186 channel=77
    4, 5, 2, 0, -3, 2, -6, 7, -3,
    -- layer=1 filter=186 channel=78
    5, -1, -1, 3, -2, -9, -11, -5, -2,
    -- layer=1 filter=186 channel=79
    -4, -8, 1, -6, -5, -5, -7, 3, 7,
    -- layer=1 filter=186 channel=80
    0, -3, 5, -7, 3, 0, 1, 5, -8,
    -- layer=1 filter=186 channel=81
    -2, -6, -2, 4, -9, 4, -5, -5, 4,
    -- layer=1 filter=186 channel=82
    0, -2, 4, -11, 1, 6, -9, 4, 3,
    -- layer=1 filter=186 channel=83
    6, -8, -2, -11, 5, -8, 0, -1, -8,
    -- layer=1 filter=186 channel=84
    -3, -4, -2, -2, -9, -11, 4, 2, 2,
    -- layer=1 filter=186 channel=85
    0, -3, 1, -4, -10, -7, 8, -1, -3,
    -- layer=1 filter=186 channel=86
    -3, -9, 0, -2, -6, -11, -3, 6, -9,
    -- layer=1 filter=186 channel=87
    5, -1, -12, 0, -2, 3, -5, 3, -11,
    -- layer=1 filter=186 channel=88
    7, -1, 0, 1, -10, 2, 7, -4, 8,
    -- layer=1 filter=186 channel=89
    0, 8, 4, -11, -10, -3, -7, 1, -5,
    -- layer=1 filter=186 channel=90
    -3, -9, -2, 5, -1, 0, -4, -8, 2,
    -- layer=1 filter=186 channel=91
    5, -9, 10, -4, -3, -10, 1, 3, -5,
    -- layer=1 filter=186 channel=92
    -12, -1, -1, -2, 0, -2, -12, -8, -3,
    -- layer=1 filter=186 channel=93
    -12, -2, -4, 7, -2, -2, -2, -5, 0,
    -- layer=1 filter=186 channel=94
    7, -8, 4, 5, -2, -2, 4, 4, -6,
    -- layer=1 filter=186 channel=95
    -11, 2, 0, 1, -1, -5, 7, -4, 7,
    -- layer=1 filter=186 channel=96
    -9, 7, -5, 3, 6, 3, 6, -5, -5,
    -- layer=1 filter=186 channel=97
    -10, 0, -5, -5, -5, -2, -4, -7, -7,
    -- layer=1 filter=186 channel=98
    0, -1, -2, 2, 10, 6, -11, -5, 2,
    -- layer=1 filter=186 channel=99
    2, -7, 5, -12, -4, 8, 0, -5, -6,
    -- layer=1 filter=186 channel=100
    -4, 0, 1, 5, 6, 1, 5, 3, -6,
    -- layer=1 filter=186 channel=101
    -9, 5, 7, -10, -2, 6, 2, 0, 6,
    -- layer=1 filter=186 channel=102
    -11, 2, 5, 6, 5, -5, 0, -10, -10,
    -- layer=1 filter=186 channel=103
    5, 0, -8, -10, 1, -12, -8, 0, -11,
    -- layer=1 filter=186 channel=104
    5, -4, -8, 2, 5, 0, 8, -10, 8,
    -- layer=1 filter=186 channel=105
    -6, 5, -8, -4, -5, -5, 0, -12, 4,
    -- layer=1 filter=186 channel=106
    -7, -2, -10, -8, 9, 7, 1, -6, 9,
    -- layer=1 filter=186 channel=107
    0, 1, -5, -3, 5, 4, -4, -8, 1,
    -- layer=1 filter=186 channel=108
    -9, -4, 3, 0, -10, -7, 3, -7, 2,
    -- layer=1 filter=186 channel=109
    0, -5, -10, 4, -4, -7, 5, 3, 2,
    -- layer=1 filter=186 channel=110
    -1, -8, -5, 5, 0, 7, -5, -4, 6,
    -- layer=1 filter=186 channel=111
    0, 11, 6, 4, -10, -10, 0, -8, -4,
    -- layer=1 filter=186 channel=112
    2, 6, -12, -7, -6, 0, 0, 7, -4,
    -- layer=1 filter=186 channel=113
    7, 0, 9, 6, 10, -3, -2, -7, 6,
    -- layer=1 filter=186 channel=114
    8, 5, -2, -7, -8, -1, -4, -10, -9,
    -- layer=1 filter=186 channel=115
    5, -1, 6, 3, -5, -1, -1, 5, -12,
    -- layer=1 filter=186 channel=116
    -1, -4, 8, 3, 4, -10, 2, -2, 6,
    -- layer=1 filter=186 channel=117
    -2, -9, -4, 6, -11, -9, -4, -9, 8,
    -- layer=1 filter=186 channel=118
    -1, -5, -7, -6, 3, -7, -3, -4, -3,
    -- layer=1 filter=186 channel=119
    6, 3, 1, 3, 3, -12, 5, 0, -5,
    -- layer=1 filter=186 channel=120
    -8, 3, -1, -11, 6, 4, 5, -3, 8,
    -- layer=1 filter=186 channel=121
    -6, 7, 6, -6, 5, -5, -8, -12, 0,
    -- layer=1 filter=186 channel=122
    4, -5, 0, -4, -10, 4, -7, 4, 10,
    -- layer=1 filter=186 channel=123
    0, 2, -5, -3, 4, 3, -11, -9, 5,
    -- layer=1 filter=186 channel=124
    5, 5, 8, -8, -5, 5, 7, 2, 0,
    -- layer=1 filter=186 channel=125
    -6, 2, -6, 5, -5, 7, -8, -8, -8,
    -- layer=1 filter=186 channel=126
    -4, -3, 7, 0, 1, -2, 4, -1, -5,
    -- layer=1 filter=186 channel=127
    9, 7, -1, 7, 0, 4, 0, -2, 6,
    -- layer=1 filter=187 channel=0
    -4, -6, 8, -8, -1, -19, -9, 2, -17,
    -- layer=1 filter=187 channel=1
    -28, 5, -11, 1, 0, 32, 6, -7, 20,
    -- layer=1 filter=187 channel=2
    -9, 0, -3, -6, -19, -3, -13, 12, 45,
    -- layer=1 filter=187 channel=3
    5, 8, 11, 0, -2, 0, -9, 0, 3,
    -- layer=1 filter=187 channel=4
    -2, -9, -10, 3, 5, -7, -1, -8, 4,
    -- layer=1 filter=187 channel=5
    -13, -12, 17, -26, 0, 23, 26, -7, 27,
    -- layer=1 filter=187 channel=6
    -31, -37, -23, -10, -47, -63, 0, -13, -4,
    -- layer=1 filter=187 channel=7
    -75, -76, -22, -83, -82, -77, -60, -59, -50,
    -- layer=1 filter=187 channel=8
    -47, -21, -4, 7, 18, 23, 22, 4, 34,
    -- layer=1 filter=187 channel=9
    6, -20, -27, -12, 10, 14, -9, -43, 15,
    -- layer=1 filter=187 channel=10
    -72, -77, -12, -80, -76, -59, -48, -45, -37,
    -- layer=1 filter=187 channel=11
    5, -3, 14, 14, 18, 10, -6, 1, 4,
    -- layer=1 filter=187 channel=12
    -28, -52, -26, -42, -23, 3, -19, 12, 12,
    -- layer=1 filter=187 channel=13
    5, -11, -31, 6, 12, -5, 1, 8, 15,
    -- layer=1 filter=187 channel=14
    -85, -27, 0, -18, 5, -35, -60, -27, -84,
    -- layer=1 filter=187 channel=15
    -61, 8, -41, 0, -20, 21, 22, -14, -22,
    -- layer=1 filter=187 channel=16
    -35, -23, 3, -4, 34, 31, 22, 15, 44,
    -- layer=1 filter=187 channel=17
    21, 11, 1, 0, -6, 4, 11, 16, -6,
    -- layer=1 filter=187 channel=18
    -37, -34, 41, 19, 14, 2, -27, -23, -4,
    -- layer=1 filter=187 channel=19
    -11, -16, -41, 3, 39, 50, -31, 10, 7,
    -- layer=1 filter=187 channel=20
    -5, -11, -17, -8, -9, -22, 1, 19, 8,
    -- layer=1 filter=187 channel=21
    -16, -21, -28, -1, -8, -11, 3, -1, 10,
    -- layer=1 filter=187 channel=22
    -14, -13, -17, 13, 15, -4, 18, 7, 26,
    -- layer=1 filter=187 channel=23
    -29, -33, -11, -23, -49, -43, -13, 1, -9,
    -- layer=1 filter=187 channel=24
    -4, -21, -53, -32, 15, 26, 6, 0, 17,
    -- layer=1 filter=187 channel=25
    -30, -39, -6, -26, -23, -8, -32, -22, 17,
    -- layer=1 filter=187 channel=26
    0, -9, -25, -19, 22, 14, 16, -11, 15,
    -- layer=1 filter=187 channel=27
    -20, -16, -20, -18, -36, -22, -18, -27, -20,
    -- layer=1 filter=187 channel=28
    -43, -54, -9, -43, -45, -47, -43, -34, -17,
    -- layer=1 filter=187 channel=29
    -24, -21, -14, -34, -15, -20, -39, -13, -16,
    -- layer=1 filter=187 channel=30
    -12, -54, 12, -9, 26, 26, -15, -19, -10,
    -- layer=1 filter=187 channel=31
    -37, -42, -14, -3, -4, -32, -41, -31, -11,
    -- layer=1 filter=187 channel=32
    -31, -32, -14, -9, 14, -2, -14, -42, 22,
    -- layer=1 filter=187 channel=33
    4, 7, -1, -7, 9, -1, -5, -7, 3,
    -- layer=1 filter=187 channel=34
    1, -3, -4, -9, 4, 5, -15, -12, -17,
    -- layer=1 filter=187 channel=35
    -5, -2, -9, -7, 0, 0, 0, -14, -17,
    -- layer=1 filter=187 channel=36
    23, 11, 17, 22, 20, 19, 12, 7, -4,
    -- layer=1 filter=187 channel=37
    -8, -12, 12, -22, 11, 36, 12, 8, 9,
    -- layer=1 filter=187 channel=38
    -15, -12, -38, -16, -21, -26, -5, -10, -11,
    -- layer=1 filter=187 channel=39
    4, -2, -16, 5, -11, -15, 7, -11, -14,
    -- layer=1 filter=187 channel=40
    -69, -82, -36, -21, -25, -43, -38, -45, -21,
    -- layer=1 filter=187 channel=41
    -1, -35, -31, 22, 40, 27, -12, -13, 18,
    -- layer=1 filter=187 channel=42
    -15, -16, -9, -28, -12, -20, -31, -40, 1,
    -- layer=1 filter=187 channel=43
    -50, -25, -16, 15, 14, 37, 6, -4, 39,
    -- layer=1 filter=187 channel=44
    -44, -12, 0, -25, 12, 19, 13, -25, 32,
    -- layer=1 filter=187 channel=45
    -36, -22, -48, -18, 1, 15, -4, -8, -2,
    -- layer=1 filter=187 channel=46
    -53, -45, -21, -31, 16, 32, -25, -15, -9,
    -- layer=1 filter=187 channel=47
    -17, -20, -41, -14, -58, -27, -16, -3, 11,
    -- layer=1 filter=187 channel=48
    -16, -4, -14, 6, -17, -9, -1, 7, -14,
    -- layer=1 filter=187 channel=49
    -15, -3, -21, -7, -22, -21, -8, -3, -3,
    -- layer=1 filter=187 channel=50
    -3, -6, 0, -25, -13, 5, -18, -16, -18,
    -- layer=1 filter=187 channel=51
    -33, -24, -29, -27, -40, -37, -5, -32, -25,
    -- layer=1 filter=187 channel=52
    4, -3, -1, -3, 3, -3, 7, 18, 11,
    -- layer=1 filter=187 channel=53
    -2, 0, -8, -10, -14, 2, 0, 2, -5,
    -- layer=1 filter=187 channel=54
    -18, -36, -20, -37, -34, 0, -33, 9, 13,
    -- layer=1 filter=187 channel=55
    6, 6, 0, 7, 0, 18, -3, 3, -8,
    -- layer=1 filter=187 channel=56
    -12, 7, 4, 1, -12, -4, -2, -7, 7,
    -- layer=1 filter=187 channel=57
    -68, -78, -44, -53, -63, -56, -33, -43, -45,
    -- layer=1 filter=187 channel=58
    -98, -93, -61, -31, -118, -71, -49, 6, -16,
    -- layer=1 filter=187 channel=59
    -1, -5, 4, -9, 4, -12, -9, -12, 0,
    -- layer=1 filter=187 channel=60
    -17, -11, -3, 0, 7, -13, -5, -8, -6,
    -- layer=1 filter=187 channel=61
    -1, -1, -1, 6, 1, 5, -5, 0, 1,
    -- layer=1 filter=187 channel=62
    -37, -28, -1, -6, 18, 37, 17, 6, 31,
    -- layer=1 filter=187 channel=63
    2, 8, 15, 17, 16, 14, 0, -12, -2,
    -- layer=1 filter=187 channel=64
    -3, 13, -1, 11, 0, 4, -1, -2, 2,
    -- layer=1 filter=187 channel=65
    0, -17, -24, 0, -12, -11, 4, -3, -1,
    -- layer=1 filter=187 channel=66
    10, 0, 4, 4, -1, 8, -9, -1, -5,
    -- layer=1 filter=187 channel=67
    10, -24, -48, 1, -10, -29, 33, -28, -6,
    -- layer=1 filter=187 channel=68
    -34, -26, -16, -37, 17, 14, 18, -25, 40,
    -- layer=1 filter=187 channel=69
    -8, -9, -34, 12, 25, 47, 37, 13, 25,
    -- layer=1 filter=187 channel=70
    6, 21, -36, -13, -31, -12, 8, -7, -31,
    -- layer=1 filter=187 channel=71
    4, -5, 0, 8, 7, 9, 0, 15, -1,
    -- layer=1 filter=187 channel=72
    -11, -51, -27, 30, 47, 6, -26, -24, 13,
    -- layer=1 filter=187 channel=73
    0, 3, 5, 10, 0, 0, 4, -3, 11,
    -- layer=1 filter=187 channel=74
    -19, -20, 18, -9, -3, 16, -36, -31, 18,
    -- layer=1 filter=187 channel=75
    -61, -38, 18, 12, 16, 7, -57, 0, -9,
    -- layer=1 filter=187 channel=76
    -14, -24, -3, -5, 9, -4, 4, -11, 5,
    -- layer=1 filter=187 channel=77
    -3, -17, -15, -5, 3, -5, 3, 9, 4,
    -- layer=1 filter=187 channel=78
    17, 8, 13, -3, 5, 12, -8, -2, 12,
    -- layer=1 filter=187 channel=79
    -14, -25, 4, 18, 31, 22, 11, 17, 23,
    -- layer=1 filter=187 channel=80
    4, -4, -7, -4, 6, -3, -4, 8, -6,
    -- layer=1 filter=187 channel=81
    -21, -24, -39, -9, 0, 1, -5, 8, 19,
    -- layer=1 filter=187 channel=82
    -31, -21, -45, 3, -26, -29, 9, -2, -1,
    -- layer=1 filter=187 channel=83
    -24, -8, -28, -18, 9, 7, 17, -11, 8,
    -- layer=1 filter=187 channel=84
    -34, -35, 51, -7, 0, 15, -12, -27, 30,
    -- layer=1 filter=187 channel=85
    -41, -54, -38, -17, -54, -52, -47, -16, -7,
    -- layer=1 filter=187 channel=86
    13, 10, 9, 12, 14, 3, 6, 0, 5,
    -- layer=1 filter=187 channel=87
    -23, -53, -32, -4, 31, 17, -39, -12, 9,
    -- layer=1 filter=187 channel=88
    -4, 3, -12, -17, -24, -16, 6, -10, -8,
    -- layer=1 filter=187 channel=89
    -32, -9, -14, -5, -29, -26, 10, 1, 13,
    -- layer=1 filter=187 channel=90
    -22, -30, -38, -38, 20, 19, 3, -28, 14,
    -- layer=1 filter=187 channel=91
    -7, -8, -13, -1, -21, -34, -6, 2, -14,
    -- layer=1 filter=187 channel=92
    -58, 20, -74, -16, -18, -7, -19, -35, -25,
    -- layer=1 filter=187 channel=93
    -2, -2, 0, 2, -8, -6, 8, 1, 4,
    -- layer=1 filter=187 channel=94
    7, -2, 18, 0, 5, 5, 1, 10, -7,
    -- layer=1 filter=187 channel=95
    -45, -37, 45, 5, 18, 21, -30, -21, 17,
    -- layer=1 filter=187 channel=96
    9, 5, -9, 3, 8, -7, 4, 5, -1,
    -- layer=1 filter=187 channel=97
    5, 1, 10, 0, 4, 2, 11, 9, 14,
    -- layer=1 filter=187 channel=98
    -31, -21, -10, 1, 25, 23, 9, 0, 38,
    -- layer=1 filter=187 channel=99
    -42, -78, -60, -76, -82, -55, -26, -40, -26,
    -- layer=1 filter=187 channel=100
    -19, -2, -10, 12, 13, 5, -21, -11, -5,
    -- layer=1 filter=187 channel=101
    -6, 0, -11, -15, -25, -19, 15, 7, 3,
    -- layer=1 filter=187 channel=102
    13, -3, -3, 14, 8, -6, 3, 9, -7,
    -- layer=1 filter=187 channel=103
    -18, -11, -1, -6, -3, -21, -15, -38, -27,
    -- layer=1 filter=187 channel=104
    -31, -9, -1, -4, -33, -7, -26, -9, -4,
    -- layer=1 filter=187 channel=105
    10, -1, -1, 4, -6, -12, -4, -2, 3,
    -- layer=1 filter=187 channel=106
    -1, -14, 0, -23, -24, -32, -14, -20, 1,
    -- layer=1 filter=187 channel=107
    -6, 2, 0, 16, -3, 2, -1, 5, 1,
    -- layer=1 filter=187 channel=108
    -31, -52, -32, -28, 11, 9, 11, -24, 20,
    -- layer=1 filter=187 channel=109
    3, 7, 1, 9, -2, 6, -6, 1, 6,
    -- layer=1 filter=187 channel=110
    -4, 0, 0, -9, -11, 8, 8, -5, 5,
    -- layer=1 filter=187 channel=111
    -22, -30, 52, -4, 2, 14, -12, -19, 11,
    -- layer=1 filter=187 channel=112
    1, 15, 59, -2, 5, 11, -17, -11, 16,
    -- layer=1 filter=187 channel=113
    -25, -29, -26, -9, -26, -25, -29, -46, -18,
    -- layer=1 filter=187 channel=114
    -40, -19, -27, -7, -7, 35, 31, -7, 14,
    -- layer=1 filter=187 channel=115
    7, 7, -6, 13, 1, 0, 7, 0, -9,
    -- layer=1 filter=187 channel=116
    2, -3, 0, -9, 2, 4, -11, 7, -4,
    -- layer=1 filter=187 channel=117
    -4, -17, 71, -10, -24, -6, 15, -4, 3,
    -- layer=1 filter=187 channel=118
    -18, -28, 38, 7, 8, 17, -14, -40, 27,
    -- layer=1 filter=187 channel=119
    -11, -47, -33, -49, 12, 0, -7, -25, 21,
    -- layer=1 filter=187 channel=120
    -9, -29, -32, -13, -15, -9, -10, -2, 2,
    -- layer=1 filter=187 channel=121
    -22, -28, -25, -4, 29, 17, -43, -34, -55,
    -- layer=1 filter=187 channel=122
    -5, 7, 0, 3, -2, 9, 5, 4, -2,
    -- layer=1 filter=187 channel=123
    -14, -1, -15, 10, 7, 4, -19, -3, -32,
    -- layer=1 filter=187 channel=124
    -7, 7, -4, 5, -2, 0, 3, -4, -10,
    -- layer=1 filter=187 channel=125
    -10, 2, -24, 14, -13, -17, 4, -31, -25,
    -- layer=1 filter=187 channel=126
    -42, -24, -3, -11, -9, -13, 3, -14, 23,
    -- layer=1 filter=187 channel=127
    -11, -36, 47, 16, 18, 19, -24, -36, 8,
    -- layer=1 filter=188 channel=0
    1, 0, 1, -2, -4, 1, 0, -11, -2,
    -- layer=1 filter=188 channel=1
    -2, -12, -12, 1, 6, -4, -13, -3, 3,
    -- layer=1 filter=188 channel=2
    -7, 0, -8, 0, -14, 2, 0, -14, -1,
    -- layer=1 filter=188 channel=3
    -8, 4, -8, -6, 2, 5, 6, 0, 2,
    -- layer=1 filter=188 channel=4
    -13, -10, -1, 5, 0, -4, -10, 6, -10,
    -- layer=1 filter=188 channel=5
    2, 5, 0, -13, 4, 5, -2, -1, 2,
    -- layer=1 filter=188 channel=6
    5, -11, -5, -2, 6, 1, -2, -10, -6,
    -- layer=1 filter=188 channel=7
    9, 0, -12, -1, 1, -1, 12, -12, -11,
    -- layer=1 filter=188 channel=8
    -2, -5, -10, 2, -1, 0, -4, 8, -11,
    -- layer=1 filter=188 channel=9
    1, -15, -3, 1, -4, -2, -12, 4, -1,
    -- layer=1 filter=188 channel=10
    -3, -11, -13, 3, -2, 5, -5, -7, -11,
    -- layer=1 filter=188 channel=11
    -11, -7, -1, 2, 1, 3, 0, 1, -1,
    -- layer=1 filter=188 channel=12
    -7, 0, 5, -4, 6, -9, -8, 5, 2,
    -- layer=1 filter=188 channel=13
    5, -5, -5, 4, 2, -6, -6, 2, 0,
    -- layer=1 filter=188 channel=14
    -9, -9, -9, -2, 7, -5, 7, -3, 3,
    -- layer=1 filter=188 channel=15
    4, 9, -4, 6, -3, 6, -9, -7, 8,
    -- layer=1 filter=188 channel=16
    10, -5, 2, -6, 5, 3, -4, -5, -13,
    -- layer=1 filter=188 channel=17
    -2, 5, -12, 2, -7, 1, 0, -11, -2,
    -- layer=1 filter=188 channel=18
    -15, -12, -3, -5, 0, 2, 3, 3, 6,
    -- layer=1 filter=188 channel=19
    -1, 2, -9, -11, 2, -1, 2, -4, 4,
    -- layer=1 filter=188 channel=20
    -8, -1, 4, -1, -3, 3, 5, -4, 1,
    -- layer=1 filter=188 channel=21
    -6, 0, 1, -12, 1, -10, -7, -3, -8,
    -- layer=1 filter=188 channel=22
    5, -1, -8, 10, 5, 3, 0, -1, 6,
    -- layer=1 filter=188 channel=23
    -6, 1, -7, 1, -7, -6, 0, -1, -5,
    -- layer=1 filter=188 channel=24
    8, 5, -6, -10, 2, -12, -9, -1, 0,
    -- layer=1 filter=188 channel=25
    -5, 1, 6, -11, 3, -1, -7, 6, -11,
    -- layer=1 filter=188 channel=26
    -3, -4, -3, 3, -9, -2, -11, -9, -2,
    -- layer=1 filter=188 channel=27
    8, -4, -4, 2, 2, 3, -1, 10, 10,
    -- layer=1 filter=188 channel=28
    0, 4, 7, 2, -1, 4, -7, -7, -8,
    -- layer=1 filter=188 channel=29
    -4, -10, -11, 0, 1, -3, 4, -7, -2,
    -- layer=1 filter=188 channel=30
    4, -5, 3, 7, -8, 4, -3, 7, -8,
    -- layer=1 filter=188 channel=31
    -2, -13, 0, -4, 2, 6, -8, -9, -10,
    -- layer=1 filter=188 channel=32
    0, -7, -12, -6, -4, -1, -4, -10, -10,
    -- layer=1 filter=188 channel=33
    -6, -1, -7, 4, 11, -1, 1, 5, 4,
    -- layer=1 filter=188 channel=34
    -6, 2, 5, 2, 1, -9, -6, -11, 6,
    -- layer=1 filter=188 channel=35
    0, 5, 3, 0, 1, 0, -5, 3, 2,
    -- layer=1 filter=188 channel=36
    -12, 7, -4, 4, -8, -11, -1, -5, 8,
    -- layer=1 filter=188 channel=37
    7, -5, -6, -13, -11, 0, 8, -8, -1,
    -- layer=1 filter=188 channel=38
    -3, -7, 6, 2, 3, -9, -4, -2, 1,
    -- layer=1 filter=188 channel=39
    -12, -10, 3, 0, 7, -3, -13, 8, -12,
    -- layer=1 filter=188 channel=40
    -9, 4, -8, -8, 1, 6, 8, 1, -7,
    -- layer=1 filter=188 channel=41
    -5, 6, -8, -4, 0, -7, -5, 1, -7,
    -- layer=1 filter=188 channel=42
    10, -13, 0, -8, 0, 0, 2, -4, -12,
    -- layer=1 filter=188 channel=43
    -10, -5, 1, -9, 1, -9, 4, -12, 1,
    -- layer=1 filter=188 channel=44
    0, -5, 6, -9, 6, 0, -10, -9, 6,
    -- layer=1 filter=188 channel=45
    -1, 5, -5, 6, 8, -12, 0, 5, 8,
    -- layer=1 filter=188 channel=46
    -14, -13, -13, 10, -2, 0, 4, -6, 6,
    -- layer=1 filter=188 channel=47
    2, -7, 2, -10, 5, -1, -5, 0, -5,
    -- layer=1 filter=188 channel=48
    -5, -4, 4, 0, -1, -2, -5, 4, 1,
    -- layer=1 filter=188 channel=49
    -1, -1, -9, 6, 7, 4, -4, -7, -10,
    -- layer=1 filter=188 channel=50
    -13, -12, 5, -3, 0, -8, 4, 8, 7,
    -- layer=1 filter=188 channel=51
    -10, 7, 1, -1, 6, 8, -1, 0, -7,
    -- layer=1 filter=188 channel=52
    5, -6, 0, -10, 2, -11, 0, 4, 2,
    -- layer=1 filter=188 channel=53
    -3, -1, 7, 4, 9, 0, -11, -4, -10,
    -- layer=1 filter=188 channel=54
    1, -11, 0, -12, 1, 0, -6, -3, 5,
    -- layer=1 filter=188 channel=55
    -4, -8, 7, 2, 6, -4, -12, -8, 2,
    -- layer=1 filter=188 channel=56
    -9, -12, -7, 4, -9, -4, 0, 4, 4,
    -- layer=1 filter=188 channel=57
    2, 3, -1, 5, -2, -3, 0, 0, 0,
    -- layer=1 filter=188 channel=58
    -1, -8, -11, -5, -13, -6, 5, 5, 0,
    -- layer=1 filter=188 channel=59
    -10, -8, -2, 7, -2, 0, -9, -4, 3,
    -- layer=1 filter=188 channel=60
    -6, -11, 3, 8, 8, 3, -1, 4, 10,
    -- layer=1 filter=188 channel=61
    -5, 0, -3, 0, -1, -3, -1, -7, -3,
    -- layer=1 filter=188 channel=62
    -1, 1, 10, 4, 5, -12, -9, -5, -12,
    -- layer=1 filter=188 channel=63
    4, 5, -12, 0, 1, 8, 9, -9, -7,
    -- layer=1 filter=188 channel=64
    -1, -12, -5, -11, 3, 5, 5, 6, 2,
    -- layer=1 filter=188 channel=65
    0, -2, -6, 2, -8, 7, 5, 3, -9,
    -- layer=1 filter=188 channel=66
    0, -7, 5, 8, 0, -3, -7, -11, -4,
    -- layer=1 filter=188 channel=67
    5, -5, 0, 5, 0, -11, 7, -6, 3,
    -- layer=1 filter=188 channel=68
    6, 7, 2, -6, -9, -2, -10, 3, 5,
    -- layer=1 filter=188 channel=69
    -4, 3, 9, -10, 0, -8, -8, -15, 5,
    -- layer=1 filter=188 channel=70
    5, -10, 0, 0, -2, -9, 4, -1, -9,
    -- layer=1 filter=188 channel=71
    -8, 0, -7, -7, -10, -9, -13, 7, -3,
    -- layer=1 filter=188 channel=72
    -6, -6, -7, 6, -9, -9, 3, -2, -3,
    -- layer=1 filter=188 channel=73
    -12, 2, -5, 0, -1, -11, -12, -9, 0,
    -- layer=1 filter=188 channel=74
    6, -9, -7, 1, 0, -9, -2, 0, -1,
    -- layer=1 filter=188 channel=75
    -5, -4, -3, -3, 8, -10, -6, -6, 2,
    -- layer=1 filter=188 channel=76
    3, 4, 1, -5, 5, -2, 6, -12, 1,
    -- layer=1 filter=188 channel=77
    -11, -3, 5, -8, 0, 0, -9, -3, 4,
    -- layer=1 filter=188 channel=78
    -9, 6, -5, 4, 4, -7, 6, -1, -12,
    -- layer=1 filter=188 channel=79
    -6, -3, 0, -8, 2, -4, 8, 2, -7,
    -- layer=1 filter=188 channel=80
    7, 3, 8, -10, 0, -4, 0, -4, 8,
    -- layer=1 filter=188 channel=81
    7, -2, 4, 4, 1, 0, -14, -11, -2,
    -- layer=1 filter=188 channel=82
    -10, -7, 0, 1, 7, -10, 0, -3, -5,
    -- layer=1 filter=188 channel=83
    -1, -12, 1, -2, -7, -7, 3, 0, 5,
    -- layer=1 filter=188 channel=84
    0, 4, -4, -9, -6, 5, 0, 10, 2,
    -- layer=1 filter=188 channel=85
    0, -3, 0, -8, -6, -7, -5, -2, 7,
    -- layer=1 filter=188 channel=86
    1, 10, 9, 3, -2, -3, 7, -11, 0,
    -- layer=1 filter=188 channel=87
    -3, -14, -2, -5, 1, 5, -8, 6, 0,
    -- layer=1 filter=188 channel=88
    2, 8, 2, -1, -5, 0, -9, 5, 0,
    -- layer=1 filter=188 channel=89
    -5, -2, 3, -9, 1, 6, -6, -4, -9,
    -- layer=1 filter=188 channel=90
    6, -10, -8, 3, -3, 5, 3, -2, 6,
    -- layer=1 filter=188 channel=91
    -1, -10, 4, 4, 1, 0, 4, -3, -9,
    -- layer=1 filter=188 channel=92
    5, 0, -4, 6, -8, -8, 1, 3, -5,
    -- layer=1 filter=188 channel=93
    -9, 0, -6, 2, 0, -5, 0, -1, -3,
    -- layer=1 filter=188 channel=94
    1, -8, -5, 2, 5, 0, -6, 0, -4,
    -- layer=1 filter=188 channel=95
    -14, 1, 3, 4, -1, -2, 0, 6, -3,
    -- layer=1 filter=188 channel=96
    4, -13, -3, 2, 4, 6, 7, 8, -1,
    -- layer=1 filter=188 channel=97
    0, -13, -2, 0, -9, -3, 2, 0, 2,
    -- layer=1 filter=188 channel=98
    5, 1, 10, -1, -10, 2, 3, -8, 4,
    -- layer=1 filter=188 channel=99
    6, -12, 5, 6, -3, -12, 5, 1, 6,
    -- layer=1 filter=188 channel=100
    -8, 2, -12, 4, -8, 5, -1, -11, 7,
    -- layer=1 filter=188 channel=101
    7, 1, 3, -4, -6, -10, -5, 0, -7,
    -- layer=1 filter=188 channel=102
    -6, -7, -12, 0, 5, 4, 4, 2, -11,
    -- layer=1 filter=188 channel=103
    -5, 6, 1, -6, -6, -11, 0, -6, 0,
    -- layer=1 filter=188 channel=104
    6, 5, -1, -2, 5, -3, 2, 7, -10,
    -- layer=1 filter=188 channel=105
    3, 0, 5, 2, -11, -11, -11, -10, 5,
    -- layer=1 filter=188 channel=106
    -12, 7, -12, -11, 0, -6, 7, 1, 7,
    -- layer=1 filter=188 channel=107
    -4, -4, 1, 1, 8, 7, 1, 2, 0,
    -- layer=1 filter=188 channel=108
    0, 3, -9, -18, 10, 2, 2, 1, 5,
    -- layer=1 filter=188 channel=109
    2, 5, -11, -10, 0, -8, -2, 9, -4,
    -- layer=1 filter=188 channel=110
    -5, -7, 3, -1, -8, 3, -10, -10, 2,
    -- layer=1 filter=188 channel=111
    4, 0, 4, -8, 0, -4, 7, 2, 8,
    -- layer=1 filter=188 channel=112
    -7, -5, 0, -6, -8, -11, 2, 4, -1,
    -- layer=1 filter=188 channel=113
    -1, -1, -4, 3, 7, -6, 0, -8, -3,
    -- layer=1 filter=188 channel=114
    -5, 1, -8, -3, -5, -8, 3, 1, -5,
    -- layer=1 filter=188 channel=115
    -9, -10, 5, 8, 5, -3, 7, 10, 7,
    -- layer=1 filter=188 channel=116
    0, 0, 5, 2, -2, -2, -6, 4, -6,
    -- layer=1 filter=188 channel=117
    3, 6, 6, -6, 4, -8, -3, -2, 6,
    -- layer=1 filter=188 channel=118
    -8, -4, -3, -7, 0, 3, 2, 7, 3,
    -- layer=1 filter=188 channel=119
    0, 0, -2, -11, 2, -8, -2, 0, 3,
    -- layer=1 filter=188 channel=120
    0, -3, -6, -8, 3, 0, -12, 6, 0,
    -- layer=1 filter=188 channel=121
    1, -2, 3, 7, 10, -6, 10, 3, -4,
    -- layer=1 filter=188 channel=122
    7, -4, -10, -5, -4, -4, -3, -5, 6,
    -- layer=1 filter=188 channel=123
    -13, 4, -5, -9, 3, -8, 7, -7, -1,
    -- layer=1 filter=188 channel=124
    -5, 3, 0, 1, 3, -12, 0, 2, -12,
    -- layer=1 filter=188 channel=125
    1, 7, 2, -3, -9, -4, 1, -5, -5,
    -- layer=1 filter=188 channel=126
    -5, 7, 3, -5, 6, 5, 0, 0, 2,
    -- layer=1 filter=188 channel=127
    4, 3, 5, 6, 2, 10, -5, -8, 9,
    -- layer=1 filter=189 channel=0
    4, -9, -10, -7, -2, 8, -6, 8, -9,
    -- layer=1 filter=189 channel=1
    1, -2, -13, -12, 7, 5, -6, -2, -8,
    -- layer=1 filter=189 channel=2
    0, -1, -8, -15, -4, -6, -12, 6, -6,
    -- layer=1 filter=189 channel=3
    1, 4, 0, -2, -3, 0, -1, 0, 0,
    -- layer=1 filter=189 channel=4
    -8, -5, 0, 0, 5, -4, 6, -7, 4,
    -- layer=1 filter=189 channel=5
    -17, -10, -5, -15, 2, 3, -12, -2, -1,
    -- layer=1 filter=189 channel=6
    -15, -4, 1, -10, 6, -17, -2, -7, -1,
    -- layer=1 filter=189 channel=7
    -11, -1, -7, 6, -2, -19, -23, -6, -13,
    -- layer=1 filter=189 channel=8
    -18, -3, -2, -11, 3, 10, 12, -9, 3,
    -- layer=1 filter=189 channel=9
    8, -2, -10, 3, -18, -12, 3, 1, 6,
    -- layer=1 filter=189 channel=10
    -9, -3, -12, 4, 1, -27, -10, -5, 1,
    -- layer=1 filter=189 channel=11
    6, -8, -8, 8, -6, 1, 7, 3, -2,
    -- layer=1 filter=189 channel=12
    -7, -16, 2, 1, 11, 6, -11, -1, 1,
    -- layer=1 filter=189 channel=13
    -15, -17, -15, -10, -1, -7, 0, -1, -12,
    -- layer=1 filter=189 channel=14
    -26, -16, 3, -6, -2, 3, -12, -4, -9,
    -- layer=1 filter=189 channel=15
    2, 7, 12, -7, 0, -14, -1, 0, -5,
    -- layer=1 filter=189 channel=16
    -17, -3, 2, 0, -9, -6, -12, -6, -11,
    -- layer=1 filter=189 channel=17
    0, 0, -3, 0, -8, -9, -6, -2, -8,
    -- layer=1 filter=189 channel=18
    -1, 1, -2, 0, -11, 1, -4, -6, -11,
    -- layer=1 filter=189 channel=19
    0, -7, -1, -10, 0, -14, -12, 1, -1,
    -- layer=1 filter=189 channel=20
    -16, -12, 2, 0, -7, -7, -7, -7, -9,
    -- layer=1 filter=189 channel=21
    -9, -16, -18, -11, -9, -18, -3, -5, -22,
    -- layer=1 filter=189 channel=22
    -10, -6, -12, 4, -6, 3, -8, -1, -18,
    -- layer=1 filter=189 channel=23
    1, 2, 11, 1, -2, 5, -8, 0, 2,
    -- layer=1 filter=189 channel=24
    1, -13, 3, -5, -11, -8, -2, -4, -2,
    -- layer=1 filter=189 channel=25
    -5, -11, -10, 9, -5, -12, -6, -14, -9,
    -- layer=1 filter=189 channel=26
    6, 4, -3, -15, -12, 0, 8, 4, 3,
    -- layer=1 filter=189 channel=27
    3, 0, -5, 7, -9, 4, -5, -5, -6,
    -- layer=1 filter=189 channel=28
    -17, -4, -10, 0, -2, -6, 0, 0, -2,
    -- layer=1 filter=189 channel=29
    -8, 5, 0, 3, 7, 0, 0, -11, 0,
    -- layer=1 filter=189 channel=30
    -8, -13, -12, 0, 2, -2, -7, -7, -2,
    -- layer=1 filter=189 channel=31
    -14, 0, -4, 0, 8, 12, -7, 6, 2,
    -- layer=1 filter=189 channel=32
    6, 2, 13, -8, -10, -6, 3, 11, -9,
    -- layer=1 filter=189 channel=33
    -5, -8, -7, -8, 0, 7, -6, 10, 1,
    -- layer=1 filter=189 channel=34
    3, -2, 6, -8, 7, -12, -12, -4, 5,
    -- layer=1 filter=189 channel=35
    4, 0, -6, 0, -4, -7, -5, 2, -3,
    -- layer=1 filter=189 channel=36
    1, -6, -9, -4, -7, -4, -11, -8, 2,
    -- layer=1 filter=189 channel=37
    -5, 6, -12, -8, 0, 3, -18, 3, -6,
    -- layer=1 filter=189 channel=38
    -2, -13, -11, -8, -1, -2, -17, -8, -15,
    -- layer=1 filter=189 channel=39
    7, -4, -7, 4, 4, -3, -5, -8, -2,
    -- layer=1 filter=189 channel=40
    -3, -15, 2, 0, 3, -12, 0, -10, 3,
    -- layer=1 filter=189 channel=41
    -4, 2, 5, -6, -3, -1, -2, 3, -13,
    -- layer=1 filter=189 channel=42
    -8, -2, 1, -5, -19, -8, -15, -19, -9,
    -- layer=1 filter=189 channel=43
    -14, -12, -15, -5, -10, -8, -6, -9, 2,
    -- layer=1 filter=189 channel=44
    3, 0, 2, -10, -1, 5, 11, 8, 1,
    -- layer=1 filter=189 channel=45
    -6, -2, -1, 0, 3, -2, 9, 10, -13,
    -- layer=1 filter=189 channel=46
    -1, -3, -2, 0, 3, -25, -13, 6, 5,
    -- layer=1 filter=189 channel=47
    -11, -1, 4, -8, 0, -3, -17, -4, 1,
    -- layer=1 filter=189 channel=48
    5, -3, 3, 2, -3, -13, -6, -1, -5,
    -- layer=1 filter=189 channel=49
    -13, 3, -9, 0, 0, -9, -13, -3, -1,
    -- layer=1 filter=189 channel=50
    -1, 4, -4, 2, 8, 0, 0, 5, 4,
    -- layer=1 filter=189 channel=51
    -4, -2, 0, -8, -2, -16, -7, -2, -14,
    -- layer=1 filter=189 channel=52
    3, 8, -1, 3, 7, -1, 11, 3, 2,
    -- layer=1 filter=189 channel=53
    0, -1, -8, -2, -8, -4, 9, -5, 6,
    -- layer=1 filter=189 channel=54
    -14, -3, -5, 7, -2, -5, -18, -8, 2,
    -- layer=1 filter=189 channel=55
    -9, -3, -2, -8, 5, -4, 0, 8, -1,
    -- layer=1 filter=189 channel=56
    0, 0, 4, -10, -10, -9, 8, 3, -2,
    -- layer=1 filter=189 channel=57
    -10, -9, -10, -6, 2, 0, 1, -11, -7,
    -- layer=1 filter=189 channel=58
    -4, 3, 9, 3, 0, -4, -6, 7, -16,
    -- layer=1 filter=189 channel=59
    9, 1, 0, -9, 0, 6, 3, -2, 6,
    -- layer=1 filter=189 channel=60
    -8, -7, 7, 0, -4, -6, -8, 10, 1,
    -- layer=1 filter=189 channel=61
    0, 5, 7, 5, -4, -7, -1, 0, 8,
    -- layer=1 filter=189 channel=62
    -15, 0, -15, -14, -2, 5, -5, -11, -3,
    -- layer=1 filter=189 channel=63
    -11, -7, 2, 0, 9, 0, -11, 7, -11,
    -- layer=1 filter=189 channel=64
    0, -3, -10, -4, -2, -2, 5, -5, -11,
    -- layer=1 filter=189 channel=65
    1, -3, -4, -2, -7, -14, -10, -1, 3,
    -- layer=1 filter=189 channel=66
    -10, -7, -12, -9, 5, -15, -1, -2, -2,
    -- layer=1 filter=189 channel=67
    0, 0, 7, -8, -16, -14, -7, -4, -9,
    -- layer=1 filter=189 channel=68
    -10, 2, 8, -11, -9, 7, 4, -4, -13,
    -- layer=1 filter=189 channel=69
    -12, 7, 12, -17, -22, -3, 4, 3, -10,
    -- layer=1 filter=189 channel=70
    -27, -8, -5, -5, -14, -8, -9, -7, -12,
    -- layer=1 filter=189 channel=71
    -2, -6, -6, 3, 0, -13, 0, -19, -12,
    -- layer=1 filter=189 channel=72
    0, -11, -17, -12, -2, 0, -14, -8, 6,
    -- layer=1 filter=189 channel=73
    6, -8, -10, 7, 6, 6, 9, -8, 3,
    -- layer=1 filter=189 channel=74
    5, 5, 0, -13, 1, -9, 2, 3, 3,
    -- layer=1 filter=189 channel=75
    -20, -3, -15, -12, -9, 6, -13, -11, 3,
    -- layer=1 filter=189 channel=76
    3, -12, 1, -15, 5, -7, -9, -2, 7,
    -- layer=1 filter=189 channel=77
    -14, -10, -5, -6, -15, -14, -8, 6, -10,
    -- layer=1 filter=189 channel=78
    -4, -2, -10, -8, -1, 0, -8, -7, 0,
    -- layer=1 filter=189 channel=79
    -3, -4, -15, -12, -12, -9, -4, 3, 0,
    -- layer=1 filter=189 channel=80
    -6, -5, -1, 3, 3, 0, -2, 8, 5,
    -- layer=1 filter=189 channel=81
    1, -6, -5, 1, 0, -6, 1, 4, -10,
    -- layer=1 filter=189 channel=82
    -15, -10, -9, -2, -1, -14, -5, 4, -5,
    -- layer=1 filter=189 channel=83
    -13, -5, -10, -5, 6, 10, -1, -10, -7,
    -- layer=1 filter=189 channel=84
    6, -3, -14, -3, 0, 4, -5, -1, -5,
    -- layer=1 filter=189 channel=85
    -8, 13, -13, -6, 7, -7, 8, 16, -9,
    -- layer=1 filter=189 channel=86
    5, 0, 0, -1, 3, -7, -8, 2, -5,
    -- layer=1 filter=189 channel=87
    -6, 1, 1, 10, 7, -4, 0, -8, 3,
    -- layer=1 filter=189 channel=88
    -4, 4, -13, 1, -17, -2, -21, -19, -12,
    -- layer=1 filter=189 channel=89
    2, -17, -15, -5, -10, -3, -12, -4, -4,
    -- layer=1 filter=189 channel=90
    -6, -8, 6, -17, -6, 6, 8, -12, 0,
    -- layer=1 filter=189 channel=91
    -1, -13, -7, -6, -9, 2, -9, -6, -3,
    -- layer=1 filter=189 channel=92
    -5, 4, -4, -15, -10, -10, 7, 4, -14,
    -- layer=1 filter=189 channel=93
    -10, 3, -11, -6, -15, -4, -3, 1, 1,
    -- layer=1 filter=189 channel=94
    1, -12, -1, -3, 2, -14, 2, 2, -5,
    -- layer=1 filter=189 channel=95
    3, -5, 4, -2, -3, 2, 0, 1, -2,
    -- layer=1 filter=189 channel=96
    4, -11, -6, -5, -3, 3, 5, 4, 2,
    -- layer=1 filter=189 channel=97
    2, -3, -3, 2, -10, -15, -1, -9, -15,
    -- layer=1 filter=189 channel=98
    -13, -11, -11, -8, 2, -3, 0, -25, -9,
    -- layer=1 filter=189 channel=99
    4, -13, 2, -11, -12, -14, -2, 4, 0,
    -- layer=1 filter=189 channel=100
    0, 2, 4, -12, -3, -7, -10, -9, -2,
    -- layer=1 filter=189 channel=101
    -10, -15, -8, -12, -9, -16, 0, -16, -17,
    -- layer=1 filter=189 channel=102
    3, -14, -12, 2, 3, -2, -13, -11, -11,
    -- layer=1 filter=189 channel=103
    11, -7, -10, 7, -2, -8, 7, -4, 0,
    -- layer=1 filter=189 channel=104
    0, 0, 3, 5, 1, -5, -3, -10, -10,
    -- layer=1 filter=189 channel=105
    -1, 4, -16, 0, -6, 0, 6, -10, 6,
    -- layer=1 filter=189 channel=106
    -11, -16, -12, -13, 4, -3, 6, -3, -20,
    -- layer=1 filter=189 channel=107
    -5, 12, -10, -3, -4, -8, -4, 4, 6,
    -- layer=1 filter=189 channel=108
    -1, -14, 9, -8, -10, -3, -3, 6, -17,
    -- layer=1 filter=189 channel=109
    10, 4, 8, 4, 2, -1, -8, 2, -7,
    -- layer=1 filter=189 channel=110
    -9, 3, -4, 2, -7, 7, 8, -1, -10,
    -- layer=1 filter=189 channel=111
    -8, -3, -13, -1, 7, 0, -2, -1, 2,
    -- layer=1 filter=189 channel=112
    -1, -12, -3, -15, 4, -14, 1, -3, 0,
    -- layer=1 filter=189 channel=113
    -8, 2, -10, -4, 3, -6, -15, -11, -9,
    -- layer=1 filter=189 channel=114
    -18, -4, 11, -7, 2, 5, 3, -14, -4,
    -- layer=1 filter=189 channel=115
    -11, 1, 0, -5, -8, 2, -1, -15, 1,
    -- layer=1 filter=189 channel=116
    8, 3, 11, 3, 0, -2, 9, 3, 8,
    -- layer=1 filter=189 channel=117
    5, -8, -8, -15, -6, -2, 10, 11, -9,
    -- layer=1 filter=189 channel=118
    0, -5, -5, -18, -13, -13, 5, 0, -2,
    -- layer=1 filter=189 channel=119
    -4, -1, -2, -7, -8, 5, -8, 1, -13,
    -- layer=1 filter=189 channel=120
    -8, 1, -7, 1, -7, 0, -5, -12, -14,
    -- layer=1 filter=189 channel=121
    -2, -7, -12, 5, 5, -3, -14, -14, 7,
    -- layer=1 filter=189 channel=122
    5, 6, -3, 8, -3, 0, -6, -8, -8,
    -- layer=1 filter=189 channel=123
    -8, 3, -6, 4, -11, 0, -8, 1, -13,
    -- layer=1 filter=189 channel=124
    -1, -5, 1, -3, -11, -1, 3, 3, -7,
    -- layer=1 filter=189 channel=125
    -2, -7, -11, -4, -10, 2, -7, -10, -12,
    -- layer=1 filter=189 channel=126
    1, -3, 1, -4, -10, 13, 12, -15, 0,
    -- layer=1 filter=189 channel=127
    -3, -9, -4, 0, 8, -7, -12, -7, 6,
    -- layer=1 filter=190 channel=0
    -17, -14, -4, -13, -17, -9, -8, -23, -11,
    -- layer=1 filter=190 channel=1
    -7, -28, -59, -54, -34, -83, 27, 39, 36,
    -- layer=1 filter=190 channel=2
    -49, -73, -65, -24, -39, -7, -18, -31, -23,
    -- layer=1 filter=190 channel=3
    1, 0, 2, -1, -7, -7, -7, 2, 2,
    -- layer=1 filter=190 channel=4
    0, 3, 1, -13, 0, -9, 13, 0, 7,
    -- layer=1 filter=190 channel=5
    -67, -123, -151, -57, -60, -65, 52, 52, 45,
    -- layer=1 filter=190 channel=6
    -75, -47, -39, -3, -36, -17, 2, -9, -33,
    -- layer=1 filter=190 channel=7
    -72, -22, -16, -89, -61, -2, 24, 28, -9,
    -- layer=1 filter=190 channel=8
    -19, -82, -115, -53, -79, -108, 28, 43, 45,
    -- layer=1 filter=190 channel=9
    7, -43, 3, -64, -24, -7, -28, -54, -12,
    -- layer=1 filter=190 channel=10
    -55, -33, 7, -36, -72, -29, 61, 36, 14,
    -- layer=1 filter=190 channel=11
    -5, -1, 0, 2, -24, -3, 5, -15, -21,
    -- layer=1 filter=190 channel=12
    -90, -22, 16, -81, -51, -29, 26, -14, 11,
    -- layer=1 filter=190 channel=13
    -26, -34, -13, 2, -19, -32, 32, 21, 25,
    -- layer=1 filter=190 channel=14
    -62, 9, 11, -59, -50, -41, 52, -4, -21,
    -- layer=1 filter=190 channel=15
    1, -73, -101, -54, -88, -31, -23, -23, 6,
    -- layer=1 filter=190 channel=16
    -48, -108, -116, -43, -61, -87, 35, 64, 46,
    -- layer=1 filter=190 channel=17
    -26, -51, -12, -20, -23, -36, 11, 2, 9,
    -- layer=1 filter=190 channel=18
    -55, -14, -13, -68, -91, -97, -24, -28, 3,
    -- layer=1 filter=190 channel=19
    -36, -99, -65, -18, -41, -17, 109, 83, 101,
    -- layer=1 filter=190 channel=20
    -15, -17, -29, -4, -26, -24, 31, 25, 17,
    -- layer=1 filter=190 channel=21
    5, 16, 24, 0, 17, 13, -3, -2, -1,
    -- layer=1 filter=190 channel=22
    23, -10, -6, -34, -36, -52, 18, 7, 28,
    -- layer=1 filter=190 channel=23
    -30, 0, -83, -57, -77, -16, -32, 1, 6,
    -- layer=1 filter=190 channel=24
    12, 9, 36, 25, 28, 29, 12, 19, 38,
    -- layer=1 filter=190 channel=25
    -65, -52, -42, -71, -81, -45, 61, 64, 24,
    -- layer=1 filter=190 channel=26
    -11, -18, 3, -37, -50, -29, 24, 1, 27,
    -- layer=1 filter=190 channel=27
    32, 30, 42, 36, 50, 43, 16, 8, 16,
    -- layer=1 filter=190 channel=28
    -5, -15, -4, 2, -49, -26, 73, 26, 9,
    -- layer=1 filter=190 channel=29
    53, 60, 51, 21, 21, 35, 22, 17, 2,
    -- layer=1 filter=190 channel=30
    -18, -54, 14, -33, -54, -54, 2, -41, -5,
    -- layer=1 filter=190 channel=31
    -66, 2, -13, -19, -29, -22, 24, 7, 39,
    -- layer=1 filter=190 channel=32
    8, -66, 13, -18, -66, -34, 32, 5, -22,
    -- layer=1 filter=190 channel=33
    21, 44, -1, 14, 3, -11, 16, 5, -12,
    -- layer=1 filter=190 channel=34
    -37, -5, -7, 23, -2, -24, 42, -25, -46,
    -- layer=1 filter=190 channel=35
    15, -5, 3, 5, 13, 4, 0, 7, 11,
    -- layer=1 filter=190 channel=36
    -9, -28, -16, -4, -27, -21, -8, -9, -8,
    -- layer=1 filter=190 channel=37
    -87, -142, -131, -64, -59, -78, 58, 64, 54,
    -- layer=1 filter=190 channel=38
    -6, -12, 0, 21, 15, 10, 24, 23, 5,
    -- layer=1 filter=190 channel=39
    10, 0, -7, 26, 2, 9, 13, 5, 12,
    -- layer=1 filter=190 channel=40
    -78, -37, -26, 3, -22, -36, 27, -4, 0,
    -- layer=1 filter=190 channel=41
    29, -31, 48, 5, -18, -30, 50, -1, 5,
    -- layer=1 filter=190 channel=42
    -51, -63, -56, -33, -36, -33, 4, 2, -3,
    -- layer=1 filter=190 channel=43
    -20, -46, -73, -34, -44, -56, 39, 47, 31,
    -- layer=1 filter=190 channel=44
    -47, -67, 0, -33, -92, -41, 8, 10, 19,
    -- layer=1 filter=190 channel=45
    -18, -8, -6, -23, -20, -6, 15, 1, 34,
    -- layer=1 filter=190 channel=46
    -75, -87, -97, -54, -70, -13, 73, 102, 101,
    -- layer=1 filter=190 channel=47
    -36, -80, -46, -58, -33, -21, 1, 23, 35,
    -- layer=1 filter=190 channel=48
    -10, 6, 10, 0, 20, 11, 0, -10, 2,
    -- layer=1 filter=190 channel=49
    -18, -29, -8, 8, -1, -3, 8, -4, -7,
    -- layer=1 filter=190 channel=50
    -13, -15, -14, -23, -22, 2, -14, -14, -12,
    -- layer=1 filter=190 channel=51
    -9, 19, -7, 13, 9, 11, 25, -6, 0,
    -- layer=1 filter=190 channel=52
    2, 7, -3, -24, -26, -12, -9, -16, 3,
    -- layer=1 filter=190 channel=53
    10, 7, 1, 0, 16, 6, 13, 10, 1,
    -- layer=1 filter=190 channel=54
    -70, -90, -55, -40, -73, -43, 75, 70, 50,
    -- layer=1 filter=190 channel=55
    14, -3, -1, 14, 2, 5, -4, -11, -16,
    -- layer=1 filter=190 channel=56
    -3, -10, -9, -9, 0, -1, 3, 1, -2,
    -- layer=1 filter=190 channel=57
    -58, -45, -7, -50, -49, -20, 69, 30, 35,
    -- layer=1 filter=190 channel=58
    -84, -43, -35, -74, -80, -17, 10, 34, 43,
    -- layer=1 filter=190 channel=59
    -21, -9, -1, -19, 0, -8, -3, -15, -3,
    -- layer=1 filter=190 channel=60
    -2, -11, -16, 7, -19, -6, -14, -19, -13,
    -- layer=1 filter=190 channel=61
    0, 5, 4, -4, -6, 2, 0, -5, 2,
    -- layer=1 filter=190 channel=62
    -67, -109, -124, -33, -72, -84, 41, 55, 57,
    -- layer=1 filter=190 channel=63
    -4, 8, 3, -7, -4, -1, -24, -25, -22,
    -- layer=1 filter=190 channel=64
    -1, -3, -3, -2, -19, -13, 4, 4, 1,
    -- layer=1 filter=190 channel=65
    5, 10, 6, 13, 7, 11, -9, -3, -18,
    -- layer=1 filter=190 channel=66
    9, 19, 8, -11, -13, 5, -19, -1, -15,
    -- layer=1 filter=190 channel=67
    -55, -37, -25, -44, -40, -22, -35, -20, -32,
    -- layer=1 filter=190 channel=68
    -51, -55, 14, -65, -93, -54, -4, -27, 14,
    -- layer=1 filter=190 channel=69
    -37, -93, -97, -30, -56, -55, 42, 63, 58,
    -- layer=1 filter=190 channel=70
    -109, -69, -75, -8, 3, -5, 35, -23, -21,
    -- layer=1 filter=190 channel=71
    22, 34, 15, 33, 35, 32, 24, 37, 35,
    -- layer=1 filter=190 channel=72
    -24, -46, 6, -47, -89, -71, 58, -50, 31,
    -- layer=1 filter=190 channel=73
    -3, 0, -2, 5, -8, -9, -6, -7, 10,
    -- layer=1 filter=190 channel=74
    -53, -13, 9, -42, -70, -68, -61, 1, -4,
    -- layer=1 filter=190 channel=75
    -31, -2, 30, -79, -90, -33, -17, -13, 39,
    -- layer=1 filter=190 channel=76
    -37, -33, 6, -39, -42, -46, -10, -19, -14,
    -- layer=1 filter=190 channel=77
    12, 21, 18, -2, 8, 14, -13, 0, -1,
    -- layer=1 filter=190 channel=78
    -22, -8, 6, 2, -9, -22, 47, 45, 3,
    -- layer=1 filter=190 channel=79
    -18, -69, -83, -9, -46, -59, 47, 60, 56,
    -- layer=1 filter=190 channel=80
    1, 16, 22, 0, -2, 9, 21, 8, 7,
    -- layer=1 filter=190 channel=81
    25, 27, 25, 16, 27, 23, 12, 18, 29,
    -- layer=1 filter=190 channel=82
    23, 18, 20, 25, 30, 13, -11, 3, 7,
    -- layer=1 filter=190 channel=83
    -41, -97, -47, -53, -87, -87, -18, -14, 23,
    -- layer=1 filter=190 channel=84
    -53, -62, -5, -68, -96, -131, -36, -29, -30,
    -- layer=1 filter=190 channel=85
    -65, -52, -46, -36, -85, -12, 16, 20, 25,
    -- layer=1 filter=190 channel=86
    -2, -8, -10, -10, -21, 6, 34, 19, 10,
    -- layer=1 filter=190 channel=87
    -46, -112, -42, -42, 1, -50, 56, 50, 25,
    -- layer=1 filter=190 channel=88
    3, 6, 1, -7, -6, 1, -25, -18, -32,
    -- layer=1 filter=190 channel=89
    0, 21, 28, 14, 25, 24, -5, -5, -9,
    -- layer=1 filter=190 channel=90
    -44, -90, -22, -49, -94, -29, 9, 17, 36,
    -- layer=1 filter=190 channel=91
    -21, -12, -11, 0, 6, 0, 11, 18, 0,
    -- layer=1 filter=190 channel=92
    4, -72, -22, -29, -76, 8, 21, -17, 56,
    -- layer=1 filter=190 channel=93
    19, 30, 27, 5, 26, 25, 14, 8, 12,
    -- layer=1 filter=190 channel=94
    -42, -25, -23, -28, -23, -11, 8, -21, -13,
    -- layer=1 filter=190 channel=95
    -54, -38, -8, -82, -86, -87, -37, -35, -6,
    -- layer=1 filter=190 channel=96
    4, 12, 11, -1, -13, -7, 6, -3, 9,
    -- layer=1 filter=190 channel=97
    17, 21, 0, -4, -3, -3, -3, 14, 11,
    -- layer=1 filter=190 channel=98
    4, -36, -44, -57, -77, -89, 29, 32, 34,
    -- layer=1 filter=190 channel=99
    -12, -33, 27, -2, -57, -64, 40, -5, -12,
    -- layer=1 filter=190 channel=100
    12, 15, 31, 20, -1, 0, 39, 3, 17,
    -- layer=1 filter=190 channel=101
    3, 2, 2, 7, 3, 1, 7, 4, 10,
    -- layer=1 filter=190 channel=102
    -52, -39, -44, -34, -39, -27, -22, -33, -15,
    -- layer=1 filter=190 channel=103
    29, 24, 28, 19, 0, 3, -2, 10, -1,
    -- layer=1 filter=190 channel=104
    1, -18, -13, -11, -42, -14, -25, 21, -7,
    -- layer=1 filter=190 channel=105
    11, 11, 20, 9, 6, -10, -7, -7, 7,
    -- layer=1 filter=190 channel=106
    -14, -32, -4, -8, -27, -27, -10, -13, -14,
    -- layer=1 filter=190 channel=107
    15, 3, 5, 17, 0, 9, 9, 0, 4,
    -- layer=1 filter=190 channel=108
    -14, -71, -27, -11, -54, -14, 20, 32, 21,
    -- layer=1 filter=190 channel=109
    -10, -10, -3, -2, 6, -3, -5, 0, 0,
    -- layer=1 filter=190 channel=110
    -14, 6, 13, 1, 0, -14, -12, -6, 0,
    -- layer=1 filter=190 channel=111
    -29, -52, 20, -47, -57, -89, -11, -18, 16,
    -- layer=1 filter=190 channel=112
    -35, -31, -14, -106, -90, -120, -55, -20, 4,
    -- layer=1 filter=190 channel=113
    -47, -26, -41, -34, -11, -1, 19, 23, -16,
    -- layer=1 filter=190 channel=114
    8, -35, -54, -29, -2, -34, 36, 57, 60,
    -- layer=1 filter=190 channel=115
    -19, -21, -4, -6, -29, 0, 50, -3, 15,
    -- layer=1 filter=190 channel=116
    8, -7, -8, -1, -5, 4, -7, 0, 8,
    -- layer=1 filter=190 channel=117
    -68, -53, -17, -77, -108, -138, -30, 0, 48,
    -- layer=1 filter=190 channel=118
    -52, -53, 7, -31, -46, -69, -13, -5, -1,
    -- layer=1 filter=190 channel=119
    0, -69, 12, -18, -66, -25, -8, -29, -3,
    -- layer=1 filter=190 channel=120
    -6, 9, -6, 5, 2, 7, 5, 35, 10,
    -- layer=1 filter=190 channel=121
    44, -6, 22, -28, -15, -2, 13, 22, 23,
    -- layer=1 filter=190 channel=122
    3, 0, 2, 9, 0, -6, -5, 5, 6,
    -- layer=1 filter=190 channel=123
    15, 14, 27, -8, -21, -6, 0, -2, 2,
    -- layer=1 filter=190 channel=124
    -10, 2, 22, 3, 28, 9, 8, -4, 8,
    -- layer=1 filter=190 channel=125
    -135, -67, -70, -25, 16, -9, -19, -9, -70,
    -- layer=1 filter=190 channel=126
    16, -11, 3, -48, -45, -105, 14, 10, 30,
    -- layer=1 filter=190 channel=127
    -67, -42, -25, -64, -91, -85, -35, -2, -5,
    -- layer=1 filter=191 channel=0
    1, 1, 8, 0, 0, -6, -8, 1, 3,
    -- layer=1 filter=191 channel=1
    7, -5, -12, -2, -5, -7, -6, -8, 1,
    -- layer=1 filter=191 channel=2
    -8, -4, -18, -9, -5, -12, -7, -17, -16,
    -- layer=1 filter=191 channel=3
    0, 9, 6, -1, -4, 1, 0, -2, -8,
    -- layer=1 filter=191 channel=4
    -6, -10, -1, 0, 7, 0, 7, 0, 0,
    -- layer=1 filter=191 channel=5
    -3, -4, -1, 4, 7, -10, -6, -10, 7,
    -- layer=1 filter=191 channel=6
    0, -13, 3, -14, -5, 2, -10, -6, -3,
    -- layer=1 filter=191 channel=7
    -22, 0, -12, 3, -7, -9, -6, -2, -13,
    -- layer=1 filter=191 channel=8
    -2, 6, -2, 3, -2, -10, -3, -9, 0,
    -- layer=1 filter=191 channel=9
    7, -17, -7, -1, -3, -1, -18, -17, -20,
    -- layer=1 filter=191 channel=10
    -13, 0, -7, 1, 0, -17, -9, -7, -17,
    -- layer=1 filter=191 channel=11
    -8, -1, 9, 0, 1, 10, 3, -7, -8,
    -- layer=1 filter=191 channel=12
    -11, -7, -8, 4, -14, 11, 6, -6, -8,
    -- layer=1 filter=191 channel=13
    -6, -2, -11, 0, -1, 4, -2, 7, 0,
    -- layer=1 filter=191 channel=14
    2, -13, -10, -7, -3, 0, -11, -7, -4,
    -- layer=1 filter=191 channel=15
    -3, 0, -2, -10, -4, 0, -2, -14, -6,
    -- layer=1 filter=191 channel=16
    -15, -2, -8, 5, -4, 0, -8, 0, 1,
    -- layer=1 filter=191 channel=17
    -4, 0, 3, 7, -7, -4, 6, 2, 3,
    -- layer=1 filter=191 channel=18
    -7, -7, 9, -11, -12, 5, -1, 0, -10,
    -- layer=1 filter=191 channel=19
    -7, 0, 2, -5, -6, -10, -7, -5, -6,
    -- layer=1 filter=191 channel=20
    0, 0, -9, -3, -8, 7, -2, 0, 8,
    -- layer=1 filter=191 channel=21
    -17, 6, -9, -4, -4, 1, -1, 0, -4,
    -- layer=1 filter=191 channel=22
    -7, 8, -2, -5, -7, -8, 8, 4, -5,
    -- layer=1 filter=191 channel=23
    4, -5, -12, -7, -8, 1, -5, -6, 8,
    -- layer=1 filter=191 channel=24
    -11, -2, 0, -1, -2, -2, 1, -12, 3,
    -- layer=1 filter=191 channel=25
    -11, 1, -18, 13, -5, -10, 1, -10, -2,
    -- layer=1 filter=191 channel=26
    -15, 0, 7, 1, -1, -4, -12, -13, -14,
    -- layer=1 filter=191 channel=27
    2, -6, -10, 0, -14, -14, 1, -12, -15,
    -- layer=1 filter=191 channel=28
    -16, -9, -2, -6, -2, -3, 9, -10, 0,
    -- layer=1 filter=191 channel=29
    -11, 0, 8, -8, 9, -10, -5, 5, -8,
    -- layer=1 filter=191 channel=30
    0, -12, -1, 7, -3, 9, -10, -4, -11,
    -- layer=1 filter=191 channel=31
    0, -9, 5, 1, 5, 6, 4, 0, -9,
    -- layer=1 filter=191 channel=32
    -7, 0, 6, -14, -9, -8, -7, -15, -3,
    -- layer=1 filter=191 channel=33
    4, 2, 2, -6, -9, 6, 3, 10, -1,
    -- layer=1 filter=191 channel=34
    1, -8, 5, -4, -6, 7, -4, 2, -10,
    -- layer=1 filter=191 channel=35
    0, 8, 0, -1, -6, 1, -4, 0, 7,
    -- layer=1 filter=191 channel=36
    -10, -2, -4, 2, 1, 0, 8, -5, 2,
    -- layer=1 filter=191 channel=37
    -1, 12, -8, -4, 4, -15, -19, -2, 9,
    -- layer=1 filter=191 channel=38
    -11, 4, 3, -2, -8, 2, -5, 1, -2,
    -- layer=1 filter=191 channel=39
    -4, -7, -10, -10, -1, 1, -2, 2, 1,
    -- layer=1 filter=191 channel=40
    -13, 5, -1, -4, -3, -7, -4, -17, -9,
    -- layer=1 filter=191 channel=41
    8, -2, 9, -8, 2, 0, -5, -9, 3,
    -- layer=1 filter=191 channel=42
    5, 6, -9, -10, -16, -10, -15, 1, -7,
    -- layer=1 filter=191 channel=43
    0, -11, 3, -4, -8, 7, 5, -3, 1,
    -- layer=1 filter=191 channel=44
    0, -15, 0, -3, -11, -4, 2, -6, -9,
    -- layer=1 filter=191 channel=45
    -7, -10, -1, 5, -8, 4, -10, 0, -10,
    -- layer=1 filter=191 channel=46
    7, 3, -5, 2, -2, -3, -9, -14, -12,
    -- layer=1 filter=191 channel=47
    -9, -21, -1, -1, -11, -5, -8, -9, -10,
    -- layer=1 filter=191 channel=48
    0, 1, -1, -4, -12, -8, 9, 4, 0,
    -- layer=1 filter=191 channel=49
    -9, -5, 6, 1, -13, -2, -7, -5, -7,
    -- layer=1 filter=191 channel=50
    -10, -4, -9, 6, 6, -8, -1, -4, -6,
    -- layer=1 filter=191 channel=51
    -12, 3, 4, 4, -9, -5, -9, 5, 1,
    -- layer=1 filter=191 channel=52
    -9, -8, -10, 0, -6, -5, -10, 2, -1,
    -- layer=1 filter=191 channel=53
    4, -1, 4, -3, 0, -3, 0, 0, -9,
    -- layer=1 filter=191 channel=54
    -11, -5, -18, -9, -14, -18, 1, -11, -10,
    -- layer=1 filter=191 channel=55
    -12, -9, -8, -4, -14, -6, -6, 3, -6,
    -- layer=1 filter=191 channel=56
    -2, 4, -6, 4, 2, 6, 4, 6, 5,
    -- layer=1 filter=191 channel=57
    -5, -10, 5, 7, 3, -11, 7, 4, -13,
    -- layer=1 filter=191 channel=58
    -18, -3, 4, 10, -12, -10, -4, -8, -13,
    -- layer=1 filter=191 channel=59
    7, -2, 4, -10, -6, 0, -8, 0, -9,
    -- layer=1 filter=191 channel=60
    -5, 1, -3, 7, 8, 5, 7, -4, 10,
    -- layer=1 filter=191 channel=61
    -1, -6, 9, -4, -5, -6, -7, 0, 5,
    -- layer=1 filter=191 channel=62
    -4, 6, 1, -5, 7, -7, -14, -9, 8,
    -- layer=1 filter=191 channel=63
    6, 0, 0, -11, -5, 7, -14, -11, -10,
    -- layer=1 filter=191 channel=64
    7, 3, -7, -8, -6, 2, -11, 6, -7,
    -- layer=1 filter=191 channel=65
    -10, 7, 9, 6, -3, -8, 8, 3, -8,
    -- layer=1 filter=191 channel=66
    -10, 1, -5, -10, -1, -1, 0, 2, -10,
    -- layer=1 filter=191 channel=67
    0, 1, 3, -15, -6, -9, 6, 0, 8,
    -- layer=1 filter=191 channel=68
    7, -13, -7, -16, 5, -13, -10, 4, 0,
    -- layer=1 filter=191 channel=69
    -1, -13, -14, -6, -16, -14, -15, -6, -6,
    -- layer=1 filter=191 channel=70
    5, -2, -9, 0, -16, 2, -2, -11, 6,
    -- layer=1 filter=191 channel=71
    -1, 8, 0, -9, -3, 2, -5, -12, -14,
    -- layer=1 filter=191 channel=72
    -3, -1, -8, -1, -3, 1, 3, -1, -12,
    -- layer=1 filter=191 channel=73
    8, -4, -10, 4, 8, 0, 1, 8, 3,
    -- layer=1 filter=191 channel=74
    -1, 4, -11, -4, 0, -9, 7, 0, 6,
    -- layer=1 filter=191 channel=75
    -3, 6, -8, -1, -4, 11, -1, -21, -13,
    -- layer=1 filter=191 channel=76
    1, 0, 2, 4, 6, -3, 0, 0, 0,
    -- layer=1 filter=191 channel=77
    7, 0, 7, 6, -6, 7, -5, 9, -3,
    -- layer=1 filter=191 channel=78
    -1, 1, 0, -8, -1, -9, 0, -4, -7,
    -- layer=1 filter=191 channel=79
    -12, -6, -13, 5, 1, 2, 3, 5, -3,
    -- layer=1 filter=191 channel=80
    3, 6, 6, 0, 8, 7, -6, -1, -10,
    -- layer=1 filter=191 channel=81
    -4, -13, -13, 0, -1, -11, -12, -1, -4,
    -- layer=1 filter=191 channel=82
    -8, 2, -6, -16, -10, -12, 6, 0, -8,
    -- layer=1 filter=191 channel=83
    0, -1, -3, -6, 3, -4, 6, -11, -10,
    -- layer=1 filter=191 channel=84
    -3, -16, -3, -4, 0, -14, -9, -13, -1,
    -- layer=1 filter=191 channel=85
    5, -3, -7, 7, -2, -6, 3, 1, 3,
    -- layer=1 filter=191 channel=86
    0, 9, -2, -2, 15, 10, 13, 8, 16,
    -- layer=1 filter=191 channel=87
    9, 4, 3, 0, -5, -7, -11, 2, -3,
    -- layer=1 filter=191 channel=88
    0, -13, 0, -5, 4, -3, 1, 0, -3,
    -- layer=1 filter=191 channel=89
    2, 2, 3, -2, 5, 7, -7, 0, 5,
    -- layer=1 filter=191 channel=90
    -5, -15, 8, 8, -3, 1, -8, 2, 6,
    -- layer=1 filter=191 channel=91
    -1, -3, -5, 1, 0, -6, 3, -6, -3,
    -- layer=1 filter=191 channel=92
    -7, -6, 3, -8, -10, -7, 2, 0, 2,
    -- layer=1 filter=191 channel=93
    -8, -12, -10, 2, 1, -10, 0, -5, -1,
    -- layer=1 filter=191 channel=94
    -5, 3, 1, 1, 2, -4, -8, 4, -11,
    -- layer=1 filter=191 channel=95
    4, -15, -1, 2, 0, 2, 2, 4, -1,
    -- layer=1 filter=191 channel=96
    -1, 3, 0, 0, 1, 8, -12, 8, -8,
    -- layer=1 filter=191 channel=97
    -1, 9, -7, -9, -9, 2, -7, 5, -10,
    -- layer=1 filter=191 channel=98
    -12, 9, -17, 4, -2, 0, 3, -1, -5,
    -- layer=1 filter=191 channel=99
    -3, 0, -6, 5, -2, -12, 5, 0, -6,
    -- layer=1 filter=191 channel=100
    7, -10, -5, 7, -5, -10, 0, 8, -11,
    -- layer=1 filter=191 channel=101
    4, -12, -6, 4, -7, -12, -11, 3, -1,
    -- layer=1 filter=191 channel=102
    -7, 0, 5, 0, -10, -10, 2, -6, -11,
    -- layer=1 filter=191 channel=103
    -7, -6, -2, 8, -9, -8, 3, 10, -5,
    -- layer=1 filter=191 channel=104
    -1, 3, -1, -10, 0, -3, -3, 0, 6,
    -- layer=1 filter=191 channel=105
    -4, -7, 7, 2, 1, -5, -10, -8, 5,
    -- layer=1 filter=191 channel=106
    -10, -7, 0, -16, 0, -7, -4, -9, -11,
    -- layer=1 filter=191 channel=107
    -6, 1, -6, 5, -3, -4, 3, 6, -7,
    -- layer=1 filter=191 channel=108
    4, -9, -1, -15, -6, -4, -17, -11, -16,
    -- layer=1 filter=191 channel=109
    -7, 4, 2, -7, 9, -2, 0, 6, -9,
    -- layer=1 filter=191 channel=110
    -6, -1, -1, 0, -10, 0, 2, 9, -5,
    -- layer=1 filter=191 channel=111
    8, -4, 12, 6, -11, -4, -3, -4, -7,
    -- layer=1 filter=191 channel=112
    -3, -4, 3, 1, -8, 1, -10, 7, -2,
    -- layer=1 filter=191 channel=113
    5, 3, -7, 8, 1, -3, -7, 0, -6,
    -- layer=1 filter=191 channel=114
    -8, -7, -5, 7, -7, 2, -10, -18, 1,
    -- layer=1 filter=191 channel=115
    7, 8, -7, 8, 11, 1, 5, -2, 2,
    -- layer=1 filter=191 channel=116
    1, 2, 4, -10, 0, 3, -4, 8, 2,
    -- layer=1 filter=191 channel=117
    4, -12, 11, -9, -3, -5, -7, -2, -2,
    -- layer=1 filter=191 channel=118
    -6, -3, 10, 0, -3, 1, -6, -4, -2,
    -- layer=1 filter=191 channel=119
    1, 3, -5, -9, -14, -5, -4, -14, 0,
    -- layer=1 filter=191 channel=120
    -7, 5, -2, -4, 5, 5, -4, -10, -11,
    -- layer=1 filter=191 channel=121
    1, 10, -10, -5, 3, 5, -6, 0, -1,
    -- layer=1 filter=191 channel=122
    7, -4, -2, -1, 2, -4, -7, 5, 2,
    -- layer=1 filter=191 channel=123
    3, 4, 0, -1, -11, 0, -8, -14, -9,
    -- layer=1 filter=191 channel=124
    7, 8, 8, -11, 2, 1, 0, 3, 0,
    -- layer=1 filter=191 channel=125
    -8, -7, -2, 0, -3, 2, 0, -8, -9,
    -- layer=1 filter=191 channel=126
    4, -9, -12, 4, 3, -3, -8, -9, -6,
    -- layer=1 filter=191 channel=127
    4, -2, 9, 2, -9, -7, -12, -3, -13,
    -- layer=1 filter=192 channel=0
    10, 1, 11, 0, -5, 0, -24, -16, -1,
    -- layer=1 filter=192 channel=1
    32, 2, 29, -30, 6, -13, -21, -19, -40,
    -- layer=1 filter=192 channel=2
    26, 41, 21, 0, 21, 15, 22, 17, 12,
    -- layer=1 filter=192 channel=3
    2, 0, -3, 0, 4, 5, 10, 3, -2,
    -- layer=1 filter=192 channel=4
    5, -10, -6, -4, 13, -1, 4, 0, 12,
    -- layer=1 filter=192 channel=5
    43, 31, 53, -62, -9, -75, -40, -51, -80,
    -- layer=1 filter=192 channel=6
    -67, -72, -22, -66, -88, -66, -20, -116, -80,
    -- layer=1 filter=192 channel=7
    19, 8, 26, 70, 11, 28, 62, 75, 15,
    -- layer=1 filter=192 channel=8
    21, 15, 35, -51, 12, -45, -76, -32, -46,
    -- layer=1 filter=192 channel=9
    3, 12, -52, -34, -26, 52, 36, -26, -31,
    -- layer=1 filter=192 channel=10
    14, 0, 30, 62, 39, 10, 54, 54, 20,
    -- layer=1 filter=192 channel=11
    24, 33, 12, 16, 14, 26, -19, -11, 5,
    -- layer=1 filter=192 channel=12
    -11, 26, 3, 10, -13, -5, -41, -52, -82,
    -- layer=1 filter=192 channel=13
    -4, -33, -40, 10, -62, -53, 6, -21, -31,
    -- layer=1 filter=192 channel=14
    7, -17, 14, 61, -2, -16, 15, 55, -12,
    -- layer=1 filter=192 channel=15
    -24, -18, 7, -26, -33, -19, -17, -62, -16,
    -- layer=1 filter=192 channel=16
    14, 20, 33, -20, -30, -66, -44, -28, -60,
    -- layer=1 filter=192 channel=17
    11, 14, 20, -12, -18, -5, -28, -26, -27,
    -- layer=1 filter=192 channel=18
    76, 51, 9, 9, 20, 5, -1, 5, -16,
    -- layer=1 filter=192 channel=19
    -13, -4, -27, -59, -21, -59, -23, -37, -31,
    -- layer=1 filter=192 channel=20
    -24, -14, -11, -27, -64, -36, -32, -39, -40,
    -- layer=1 filter=192 channel=21
    -11, -25, 12, 3, -26, 0, -14, -3, -11,
    -- layer=1 filter=192 channel=22
    -27, -39, -11, -42, -35, -22, -22, -27, -31,
    -- layer=1 filter=192 channel=23
    9, 27, 12, 49, 66, 28, 60, 60, 34,
    -- layer=1 filter=192 channel=24
    0, 19, 7, 1, -4, 7, 22, -2, 17,
    -- layer=1 filter=192 channel=25
    6, -13, -8, 34, -19, -41, 27, 36, -37,
    -- layer=1 filter=192 channel=26
    7, 8, -12, 18, -15, -21, 27, -11, -17,
    -- layer=1 filter=192 channel=27
    -32, -33, -1, -21, -24, 3, -10, -9, 1,
    -- layer=1 filter=192 channel=28
    -28, -21, 9, 38, 1, 1, 42, 48, 12,
    -- layer=1 filter=192 channel=29
    -55, -24, -28, -38, -23, 3, -22, -14, -19,
    -- layer=1 filter=192 channel=30
    56, 46, 8, -18, 25, -14, -5, -18, -21,
    -- layer=1 filter=192 channel=31
    5, -8, -13, -6, -25, -40, -52, -60, -60,
    -- layer=1 filter=192 channel=32
    -1, 19, -15, 22, 0, -20, 64, 23, -7,
    -- layer=1 filter=192 channel=33
    -10, -7, 0, 9, -10, 4, 7, -19, 10,
    -- layer=1 filter=192 channel=34
    0, -8, -13, 8, -14, -9, -12, -17, -16,
    -- layer=1 filter=192 channel=35
    -12, 1, -7, -19, -10, -8, -9, -15, -17,
    -- layer=1 filter=192 channel=36
    43, 39, 32, 18, 26, 21, -9, 3, 10,
    -- layer=1 filter=192 channel=37
    28, 30, 36, -21, -36, -80, -34, -49, -84,
    -- layer=1 filter=192 channel=38
    -24, -35, 12, -19, -59, -29, -14, -37, -11,
    -- layer=1 filter=192 channel=39
    12, 4, 20, -21, 13, -9, -17, -27, -19,
    -- layer=1 filter=192 channel=40
    -25, -42, -47, -31, -32, -50, -31, -41, -41,
    -- layer=1 filter=192 channel=41
    -21, 67, 4, 12, -22, -3, 80, -23, -1,
    -- layer=1 filter=192 channel=42
    33, 40, 17, 22, 19, -23, -3, -8, -26,
    -- layer=1 filter=192 channel=43
    0, 7, 34, -30, -38, -59, -26, -16, -55,
    -- layer=1 filter=192 channel=44
    0, 4, -18, 53, 11, 4, 60, 26, 0,
    -- layer=1 filter=192 channel=45
    2, 9, 8, -27, 3, -18, 10, -26, -1,
    -- layer=1 filter=192 channel=46
    -50, -45, 19, -57, -70, -66, -62, -89, -103,
    -- layer=1 filter=192 channel=47
    -20, 44, 12, 51, 8, 3, 65, 15, 13,
    -- layer=1 filter=192 channel=48
    -17, -25, 2, -26, -11, -7, -6, -18, -7,
    -- layer=1 filter=192 channel=49
    -28, 5, 6, -27, -31, 6, 23, -14, -4,
    -- layer=1 filter=192 channel=50
    11, -16, -11, 2, -2, 15, 6, -35, -14,
    -- layer=1 filter=192 channel=51
    1, -30, 4, 20, 0, -5, 7, 0, -6,
    -- layer=1 filter=192 channel=52
    26, 19, 21, 14, 24, -2, 19, 6, 11,
    -- layer=1 filter=192 channel=53
    -1, 20, 2, 13, 15, -11, -8, 1, 6,
    -- layer=1 filter=192 channel=54
    -6, -12, -4, 35, -22, -57, 23, 36, -39,
    -- layer=1 filter=192 channel=55
    20, 30, 13, 12, 15, 18, 0, 11, 9,
    -- layer=1 filter=192 channel=56
    2, 8, 2, -7, -7, 5, -5, 5, 14,
    -- layer=1 filter=192 channel=57
    0, -34, -10, 35, -7, -4, 38, 15, 7,
    -- layer=1 filter=192 channel=58
    47, 32, 24, 83, 59, 12, 106, 77, 56,
    -- layer=1 filter=192 channel=59
    -1, 3, -15, -5, -1, -5, -6, -10, -9,
    -- layer=1 filter=192 channel=60
    -14, -15, -13, 1, -17, -2, -13, -21, 6,
    -- layer=1 filter=192 channel=61
    -9, -2, 8, -10, -8, -10, -10, -1, 7,
    -- layer=1 filter=192 channel=62
    20, 0, 28, -41, -33, -87, -59, -34, -68,
    -- layer=1 filter=192 channel=63
    48, 32, 26, 20, 22, 34, 6, 1, 5,
    -- layer=1 filter=192 channel=64
    -5, -5, 6, -6, -8, 9, 0, -14, -3,
    -- layer=1 filter=192 channel=65
    -29, -13, 10, -18, -21, -1, -24, -18, 3,
    -- layer=1 filter=192 channel=66
    5, 4, 25, -6, 13, 6, -11, -12, 2,
    -- layer=1 filter=192 channel=67
    -1, 10, 29, 7, -19, 15, -25, -20, 17,
    -- layer=1 filter=192 channel=68
    37, 21, -16, 61, -8, 13, 60, 48, 11,
    -- layer=1 filter=192 channel=69
    0, 4, -9, -24, -13, -65, -24, -52, -43,
    -- layer=1 filter=192 channel=70
    -57, -11, 40, -63, -25, 14, -48, -93, -60,
    -- layer=1 filter=192 channel=71
    -22, 1, 8, -14, -7, -1, -7, 30, -4,
    -- layer=1 filter=192 channel=72
    18, 32, 6, -17, 1, -27, -1, -54, -31,
    -- layer=1 filter=192 channel=73
    -5, -4, -6, 0, -3, -8, -6, -2, 6,
    -- layer=1 filter=192 channel=74
    12, -19, -34, 20, -23, -12, 26, -18, -15,
    -- layer=1 filter=192 channel=75
    32, -2, 21, 2, 8, -35, 6, 2, -47,
    -- layer=1 filter=192 channel=76
    37, 33, 2, 17, -4, 6, 16, 4, -11,
    -- layer=1 filter=192 channel=77
    -5, -31, -1, -12, -8, -2, -21, -9, 0,
    -- layer=1 filter=192 channel=78
    -12, -15, 0, 16, -13, 0, 12, 2, 4,
    -- layer=1 filter=192 channel=79
    4, 11, 11, -30, -13, -67, -57, -51, -59,
    -- layer=1 filter=192 channel=80
    1, -11, -2, -2, -5, -9, -5, -5, -5,
    -- layer=1 filter=192 channel=81
    -20, 6, -2, -10, -9, 1, -6, 8, 6,
    -- layer=1 filter=192 channel=82
    -29, -28, 1, -28, -24, 0, -2, -24, -12,
    -- layer=1 filter=192 channel=83
    12, 6, -3, -24, 9, -45, 3, -21, -9,
    -- layer=1 filter=192 channel=84
    49, 44, 4, 18, -8, -9, 36, -1, -30,
    -- layer=1 filter=192 channel=85
    -3, 31, 18, 44, 58, -3, 70, 53, 14,
    -- layer=1 filter=192 channel=86
    18, 16, 24, -19, -3, 12, -28, -26, -25,
    -- layer=1 filter=192 channel=87
    -28, -8, -43, -78, -61, -40, -35, -58, -46,
    -- layer=1 filter=192 channel=88
    -7, 5, 16, -20, 0, 23, -25, 1, 4,
    -- layer=1 filter=192 channel=89
    -17, -25, 3, -2, -30, -11, 8, -21, -10,
    -- layer=1 filter=192 channel=90
    19, 3, -15, 34, 8, -11, 55, 29, -2,
    -- layer=1 filter=192 channel=91
    -3, -16, -13, 2, -45, -31, 7, -32, -29,
    -- layer=1 filter=192 channel=92
    -17, -23, -6, 0, -30, 15, 34, -7, -17,
    -- layer=1 filter=192 channel=93
    -12, 12, 2, -9, 8, 1, -3, -8, -3,
    -- layer=1 filter=192 channel=94
    10, 21, 12, 6, 5, 5, -24, -7, -5,
    -- layer=1 filter=192 channel=95
    49, 40, 3, 40, 3, -4, 25, 11, -16,
    -- layer=1 filter=192 channel=96
    2, 3, -4, 1, 8, -3, 0, 3, 8,
    -- layer=1 filter=192 channel=97
    21, 0, 22, -7, 0, 15, -13, 4, 1,
    -- layer=1 filter=192 channel=98
    -3, -11, 14, -39, -26, -67, -42, -17, -39,
    -- layer=1 filter=192 channel=99
    -19, -21, 5, 35, 64, 28, 33, 86, 52,
    -- layer=1 filter=192 channel=100
    25, 16, 24, 6, 0, 5, -10, -7, 3,
    -- layer=1 filter=192 channel=101
    -10, -31, -13, -5, -46, -10, -15, -26, -22,
    -- layer=1 filter=192 channel=102
    20, 1, 19, 2, -3, -3, -31, -25, -2,
    -- layer=1 filter=192 channel=103
    20, 15, 9, -10, -5, 9, -10, -12, -12,
    -- layer=1 filter=192 channel=104
    -19, 28, -4, 5, 31, -2, 38, 21, 13,
    -- layer=1 filter=192 channel=105
    14, 13, 20, -3, 9, 24, -5, 11, 8,
    -- layer=1 filter=192 channel=106
    -7, -14, -46, -2, -30, -39, 23, -17, -25,
    -- layer=1 filter=192 channel=107
    -4, 3, 3, -10, 2, 0, -5, -10, -11,
    -- layer=1 filter=192 channel=108
    -13, 13, -20, 44, 10, 1, 62, 29, 17,
    -- layer=1 filter=192 channel=109
    2, -5, 0, 6, 2, -7, 8, 0, -3,
    -- layer=1 filter=192 channel=110
    1, -7, 5, -6, -1, -13, -6, 8, -16,
    -- layer=1 filter=192 channel=111
    54, 43, 6, 3, 19, 7, -9, -2, -17,
    -- layer=1 filter=192 channel=112
    33, 6, -2, 13, -2, -3, -13, -30, -12,
    -- layer=1 filter=192 channel=113
    3, 0, 7, -1, -36, -25, -8, -35, -18,
    -- layer=1 filter=192 channel=114
    8, 5, 4, -55, 0, -61, -34, -91, -58,
    -- layer=1 filter=192 channel=115
    2, -1, 22, -17, -6, 8, -24, -9, -12,
    -- layer=1 filter=192 channel=116
    4, -10, 1, 4, -6, 0, 4, -8, 1,
    -- layer=1 filter=192 channel=117
    28, -13, -24, -29, -8, -24, -33, -24, -7,
    -- layer=1 filter=192 channel=118
    50, 43, -7, -10, -6, -10, 7, -20, -25,
    -- layer=1 filter=192 channel=119
    4, 37, -14, 21, 1, 1, 70, 16, 22,
    -- layer=1 filter=192 channel=120
    -1, 0, -16, 21, -17, -22, 15, 5, -35,
    -- layer=1 filter=192 channel=121
    9, 11, 10, -25, -13, -25, -18, 10, -11,
    -- layer=1 filter=192 channel=122
    -9, -4, 0, -2, -10, -10, 3, 8, -10,
    -- layer=1 filter=192 channel=123
    27, 10, 0, 14, 20, 2, 2, 25, 14,
    -- layer=1 filter=192 channel=124
    -12, -7, 1, -16, -7, 0, -10, 2, 1,
    -- layer=1 filter=192 channel=125
    -15, 12, 57, -84, -47, 16, -47, -122, -46,
    -- layer=1 filter=192 channel=126
    12, -11, 11, -45, -28, -57, -51, -36, -34,
    -- layer=1 filter=192 channel=127
    50, 34, 7, 14, 11, -5, 0, -20, -28,
    -- layer=1 filter=193 channel=0
    -1, 3, -12, -6, -11, 1, 7, 0, 6,
    -- layer=1 filter=193 channel=1
    -3, -9, -9, 4, 3, 1, 5, -11, -2,
    -- layer=1 filter=193 channel=2
    -5, -9, 2, -5, -6, -11, 4, -7, 2,
    -- layer=1 filter=193 channel=3
    2, -4, -10, -3, -9, -7, -8, 5, 3,
    -- layer=1 filter=193 channel=4
    -10, 8, 9, 4, -1, -8, 1, -2, 2,
    -- layer=1 filter=193 channel=5
    7, 4, 6, -7, 4, -14, -9, 0, -3,
    -- layer=1 filter=193 channel=6
    3, -13, -2, -8, 6, -4, -10, -4, -4,
    -- layer=1 filter=193 channel=7
    1, -4, 0, -9, -9, -6, 3, -2, -6,
    -- layer=1 filter=193 channel=8
    0, -10, -9, -5, 0, 4, 3, -4, -10,
    -- layer=1 filter=193 channel=9
    2, -3, -10, 2, -1, 1, 1, -2, -10,
    -- layer=1 filter=193 channel=10
    -13, -7, 4, 0, -8, -3, -7, -13, -10,
    -- layer=1 filter=193 channel=11
    -11, 3, 0, -11, -2, -2, 0, 5, 0,
    -- layer=1 filter=193 channel=12
    -3, 7, -2, 0, 2, 1, 4, -4, -4,
    -- layer=1 filter=193 channel=13
    1, -6, -14, -8, -9, -8, 0, -5, -2,
    -- layer=1 filter=193 channel=14
    -5, -10, 5, 2, 0, -3, 0, -5, -6,
    -- layer=1 filter=193 channel=15
    5, 1, -2, -1, 0, 0, 8, 2, 3,
    -- layer=1 filter=193 channel=16
    0, -9, 1, 8, 8, -5, -3, -5, -4,
    -- layer=1 filter=193 channel=17
    4, -5, -11, -11, -3, -8, -8, 0, -1,
    -- layer=1 filter=193 channel=18
    0, -13, -15, -4, -8, -7, 2, 2, 4,
    -- layer=1 filter=193 channel=19
    7, -11, -3, -1, -4, 6, 0, 1, 3,
    -- layer=1 filter=193 channel=20
    2, -4, -2, -5, 2, -1, 0, -10, -8,
    -- layer=1 filter=193 channel=21
    -2, -12, -10, 4, 2, -10, -9, -3, 8,
    -- layer=1 filter=193 channel=22
    -8, 4, -3, 7, 0, 0, 6, 0, -5,
    -- layer=1 filter=193 channel=23
    0, 9, -7, 8, -1, -13, 5, -1, -10,
    -- layer=1 filter=193 channel=24
    0, -4, -14, -11, 6, -10, -3, -5, -3,
    -- layer=1 filter=193 channel=25
    -2, 3, 6, -6, -7, -9, 6, 2, 3,
    -- layer=1 filter=193 channel=26
    -11, -6, 5, -6, 0, -4, 4, -7, -8,
    -- layer=1 filter=193 channel=27
    4, 2, 10, -2, 0, 0, 7, 3, 6,
    -- layer=1 filter=193 channel=28
    -14, -13, -6, 6, -3, -8, 2, -10, -7,
    -- layer=1 filter=193 channel=29
    1, 4, 1, -2, -10, -1, -1, -1, -6,
    -- layer=1 filter=193 channel=30
    -7, -11, -16, 0, -5, -10, 7, 4, -10,
    -- layer=1 filter=193 channel=31
    -4, 2, 0, 0, -10, 2, -8, -3, -7,
    -- layer=1 filter=193 channel=32
    2, -5, 3, -9, -10, 0, -4, 7, 1,
    -- layer=1 filter=193 channel=33
    -7, 2, 3, -6, 3, -5, -10, 6, 1,
    -- layer=1 filter=193 channel=34
    -4, 7, -9, -7, -4, 8, 1, 3, 0,
    -- layer=1 filter=193 channel=35
    7, 2, 9, -3, 2, -3, 7, 6, -5,
    -- layer=1 filter=193 channel=36
    -8, -6, 0, 3, -6, -7, -10, -1, 1,
    -- layer=1 filter=193 channel=37
    2, 4, 3, -5, -11, 0, 0, 1, 2,
    -- layer=1 filter=193 channel=38
    -6, 4, -7, -4, 5, 0, 4, -8, 5,
    -- layer=1 filter=193 channel=39
    -5, -1, 1, -4, -7, -7, 6, 0, -6,
    -- layer=1 filter=193 channel=40
    3, 5, 6, -1, -1, -5, 6, -2, -2,
    -- layer=1 filter=193 channel=41
    -3, 6, -8, 0, 3, 1, 5, 7, -14,
    -- layer=1 filter=193 channel=42
    3, 0, 10, 4, -3, -7, 0, 1, 9,
    -- layer=1 filter=193 channel=43
    1, -5, 7, -7, -7, -1, 0, -3, 1,
    -- layer=1 filter=193 channel=44
    -8, 5, 1, 7, -3, 6, -3, -7, 0,
    -- layer=1 filter=193 channel=45
    -3, -4, 3, -10, -9, -1, -5, 6, 6,
    -- layer=1 filter=193 channel=46
    7, -9, 6, 7, -5, -8, -5, -3, 0,
    -- layer=1 filter=193 channel=47
    7, 1, -5, -1, 4, -3, -12, 9, -6,
    -- layer=1 filter=193 channel=48
    -5, 5, 6, 2, -3, -1, 2, -1, -5,
    -- layer=1 filter=193 channel=49
    3, -3, -12, 2, -5, 0, 0, -3, -7,
    -- layer=1 filter=193 channel=50
    9, -3, 5, 9, -9, 3, 3, -7, -6,
    -- layer=1 filter=193 channel=51
    5, -5, -10, 3, -4, 2, 10, -1, 7,
    -- layer=1 filter=193 channel=52
    8, 9, -2, -8, -3, 2, -7, -9, -4,
    -- layer=1 filter=193 channel=53
    -2, -3, 2, -1, 4, 4, -7, 2, 7,
    -- layer=1 filter=193 channel=54
    -14, -9, 1, 2, -4, 9, 6, 0, 1,
    -- layer=1 filter=193 channel=55
    5, 0, 0, 6, -4, 3, 6, -7, 2,
    -- layer=1 filter=193 channel=56
    -3, 3, 3, -2, -9, -9, 6, -9, -4,
    -- layer=1 filter=193 channel=57
    -10, 1, 8, -13, 5, -8, -4, -7, 7,
    -- layer=1 filter=193 channel=58
    4, -4, -2, -2, 2, -7, -8, 5, 4,
    -- layer=1 filter=193 channel=59
    -7, -10, -2, -11, -1, 4, 10, -1, 6,
    -- layer=1 filter=193 channel=60
    -5, -3, 3, 1, 5, -8, -2, -6, -6,
    -- layer=1 filter=193 channel=61
    4, 9, -5, 8, 7, -9, 6, 0, -8,
    -- layer=1 filter=193 channel=62
    -1, 0, -9, 4, 6, -7, -1, 4, -7,
    -- layer=1 filter=193 channel=63
    -6, -9, -6, -8, -6, 3, 4, 0, 6,
    -- layer=1 filter=193 channel=64
    -8, 2, 7, -10, -5, 0, -7, -9, 2,
    -- layer=1 filter=193 channel=65
    0, -11, -5, -10, 2, -8, 3, -7, 0,
    -- layer=1 filter=193 channel=66
    -1, -11, -1, 0, 4, 7, 0, 2, -3,
    -- layer=1 filter=193 channel=67
    7, -7, 7, -5, 0, 7, -8, 5, 6,
    -- layer=1 filter=193 channel=68
    8, 8, 0, -1, -8, -5, -6, 0, -7,
    -- layer=1 filter=193 channel=69
    -2, 3, 6, -5, 9, -12, -6, -6, 1,
    -- layer=1 filter=193 channel=70
    -6, 5, 9, -11, -7, 1, 1, 0, 1,
    -- layer=1 filter=193 channel=71
    0, 6, -1, -3, -1, -5, -10, 3, 1,
    -- layer=1 filter=193 channel=72
    -3, 6, -1, 10, 6, -6, -3, -7, 0,
    -- layer=1 filter=193 channel=73
    -10, -4, -6, -10, -5, -3, 7, 10, -10,
    -- layer=1 filter=193 channel=74
    5, -4, -7, -4, -9, -8, -7, -1, -6,
    -- layer=1 filter=193 channel=75
    4, -8, -5, -6, -9, 5, -11, -5, 8,
    -- layer=1 filter=193 channel=76
    -3, 2, 4, 9, 2, -4, -5, 8, 1,
    -- layer=1 filter=193 channel=77
    -8, 5, 6, -3, -4, -3, 5, 0, -3,
    -- layer=1 filter=193 channel=78
    10, -1, 6, -6, -6, 3, 1, -11, 0,
    -- layer=1 filter=193 channel=79
    -3, 7, -7, -10, -2, 1, -8, 0, -7,
    -- layer=1 filter=193 channel=80
    -8, -4, 2, 9, -6, -2, -2, 8, -2,
    -- layer=1 filter=193 channel=81
    -2, 0, 2, -1, 1, -9, 2, 4, 2,
    -- layer=1 filter=193 channel=82
    3, 5, -3, 2, 6, 2, -12, -3, -8,
    -- layer=1 filter=193 channel=83
    -8, 3, -2, -5, -10, 1, 8, 1, -8,
    -- layer=1 filter=193 channel=84
    -2, -6, -12, 7, -10, 2, 1, -11, -8,
    -- layer=1 filter=193 channel=85
    -6, -10, -4, 2, -4, -6, 5, -5, -8,
    -- layer=1 filter=193 channel=86
    -3, -9, -8, 3, -4, -11, -5, -5, -11,
    -- layer=1 filter=193 channel=87
    7, 0, -9, -1, -5, 6, 1, -7, -8,
    -- layer=1 filter=193 channel=88
    -4, -7, 6, 7, -7, 2, 9, 4, -9,
    -- layer=1 filter=193 channel=89
    -7, 6, 1, -3, -2, -2, -5, 10, -6,
    -- layer=1 filter=193 channel=90
    7, 0, -10, -3, 4, 0, 4, -1, 2,
    -- layer=1 filter=193 channel=91
    -8, -11, -8, -1, 5, -12, 4, 6, -9,
    -- layer=1 filter=193 channel=92
    7, -2, -7, 5, -10, 0, -6, 2, -7,
    -- layer=1 filter=193 channel=93
    -14, -10, 4, -4, 0, -5, -6, -7, -8,
    -- layer=1 filter=193 channel=94
    0, 0, 0, -3, -6, -11, -6, -8, -4,
    -- layer=1 filter=193 channel=95
    -1, 4, 4, -6, -6, 5, 3, 5, -6,
    -- layer=1 filter=193 channel=96
    -3, 8, -4, -1, -10, -3, 3, 6, 2,
    -- layer=1 filter=193 channel=97
    -11, 0, -4, 0, -7, -3, 9, 8, -5,
    -- layer=1 filter=193 channel=98
    -1, 0, -2, 5, 4, 7, 5, 2, 9,
    -- layer=1 filter=193 channel=99
    -2, -4, 9, 1, -16, 0, 4, -3, -7,
    -- layer=1 filter=193 channel=100
    -4, -6, 0, -10, 5, -1, -10, 5, 6,
    -- layer=1 filter=193 channel=101
    6, -7, -1, 0, 6, -11, -9, 6, -9,
    -- layer=1 filter=193 channel=102
    -3, -6, 4, -3, -8, -9, -3, -1, 8,
    -- layer=1 filter=193 channel=103
    -4, 8, -7, -3, 2, 5, -3, 0, 2,
    -- layer=1 filter=193 channel=104
    4, -3, 0, -11, -9, 4, 2, -2, 5,
    -- layer=1 filter=193 channel=105
    -2, -5, -8, 6, 5, 8, -7, -11, -12,
    -- layer=1 filter=193 channel=106
    0, 1, -11, -9, 8, -1, 0, -2, -4,
    -- layer=1 filter=193 channel=107
    3, 5, 0, 1, 0, 0, 5, 9, 0,
    -- layer=1 filter=193 channel=108
    -10, -9, -1, 2, 0, -3, 8, 0, 1,
    -- layer=1 filter=193 channel=109
    3, -6, -9, 4, -7, 6, 1, 1, -9,
    -- layer=1 filter=193 channel=110
    7, 2, -5, -3, -5, 0, -7, 0, 3,
    -- layer=1 filter=193 channel=111
    -11, 2, 2, 0, 6, -9, 0, 2, 6,
    -- layer=1 filter=193 channel=112
    -8, 0, -5, -2, -7, 0, -11, -4, -13,
    -- layer=1 filter=193 channel=113
    5, 3, 2, 5, -5, -4, -4, 7, 0,
    -- layer=1 filter=193 channel=114
    0, -3, 8, -7, 5, -5, 0, -6, -3,
    -- layer=1 filter=193 channel=115
    -6, -7, 9, -3, -1, -8, 1, -5, -2,
    -- layer=1 filter=193 channel=116
    9, 1, -1, 0, 6, -2, 9, -8, -2,
    -- layer=1 filter=193 channel=117
    6, 3, -10, 2, 6, -1, 4, 4, 6,
    -- layer=1 filter=193 channel=118
    0, 1, 6, -7, 0, -4, 3, 4, 5,
    -- layer=1 filter=193 channel=119
    0, -8, 3, 6, 10, 4, -8, 2, -3,
    -- layer=1 filter=193 channel=120
    -3, 7, -4, 1, -5, -13, -8, -11, -12,
    -- layer=1 filter=193 channel=121
    -5, -9, -10, -13, 0, 5, -9, -13, -7,
    -- layer=1 filter=193 channel=122
    6, 1, -4, -5, 1, -5, -5, -9, -5,
    -- layer=1 filter=193 channel=123
    -6, 2, 3, 5, 8, -6, -2, 0, -1,
    -- layer=1 filter=193 channel=124
    6, 3, -10, 5, 5, 3, 4, 6, -7,
    -- layer=1 filter=193 channel=125
    0, 1, -11, -12, -2, 4, 8, 1, 5,
    -- layer=1 filter=193 channel=126
    6, -1, 9, 1, 6, -1, -3, -1, -5,
    -- layer=1 filter=193 channel=127
    6, -11, -2, -5, 4, -7, -4, -10, -6,
    -- layer=1 filter=194 channel=0
    0, 5, -11, 6, -6, 1, -8, 8, -5,
    -- layer=1 filter=194 channel=1
    -10, 3, 5, -4, -4, -8, -8, 3, -4,
    -- layer=1 filter=194 channel=2
    -1, -4, 2, 6, 1, 2, 3, -2, 11,
    -- layer=1 filter=194 channel=3
    -7, 0, -5, 5, -2, 3, -2, -8, -6,
    -- layer=1 filter=194 channel=4
    -2, -2, 0, -6, 1, -3, 5, 7, -4,
    -- layer=1 filter=194 channel=5
    -6, 3, -7, -20, -9, -22, -12, -9, -6,
    -- layer=1 filter=194 channel=6
    8, -2, 2, 8, 6, -7, -10, -11, -15,
    -- layer=1 filter=194 channel=7
    -3, -1, -3, -13, -17, 1, 0, -13, -8,
    -- layer=1 filter=194 channel=8
    -7, -2, -10, -16, -6, -17, -3, -13, -1,
    -- layer=1 filter=194 channel=9
    -11, 10, -2, -5, -1, -1, -9, -8, 3,
    -- layer=1 filter=194 channel=10
    -1, -14, 9, 4, -7, -8, 6, -9, 0,
    -- layer=1 filter=194 channel=11
    -12, -6, 3, -3, -9, -1, -4, -14, -14,
    -- layer=1 filter=194 channel=12
    1, -12, 9, 18, 8, 1, 2, -7, 2,
    -- layer=1 filter=194 channel=13
    2, 0, -3, -1, -6, -5, -9, -4, -6,
    -- layer=1 filter=194 channel=14
    12, -4, 1, -1, -1, -5, 7, 4, 0,
    -- layer=1 filter=194 channel=15
    -10, -7, -9, 8, -7, 0, -6, 1, 0,
    -- layer=1 filter=194 channel=16
    -27, -3, -6, -26, -23, -32, -14, -5, -4,
    -- layer=1 filter=194 channel=17
    -14, 2, -11, 2, -12, -8, 4, -2, -10,
    -- layer=1 filter=194 channel=18
    -8, -8, 0, -7, -8, 4, -14, -18, -20,
    -- layer=1 filter=194 channel=19
    -3, 0, -4, -9, 0, -12, -9, -9, 7,
    -- layer=1 filter=194 channel=20
    0, -14, -2, -17, -21, -22, -22, -6, -23,
    -- layer=1 filter=194 channel=21
    -1, 9, -9, -2, 12, 7, 0, -7, -6,
    -- layer=1 filter=194 channel=22
    -15, -1, -16, -19, -19, -19, -14, -18, -23,
    -- layer=1 filter=194 channel=23
    0, -4, -9, 1, -6, -4, -4, -8, 0,
    -- layer=1 filter=194 channel=24
    7, 10, -1, 9, -7, 5, 12, 10, 11,
    -- layer=1 filter=194 channel=25
    -20, -7, 4, -9, -16, -11, -6, -9, -5,
    -- layer=1 filter=194 channel=26
    -7, -14, -18, -2, -5, -4, 2, -9, -26,
    -- layer=1 filter=194 channel=27
    -15, -7, 0, -4, -6, 0, 3, 0, -3,
    -- layer=1 filter=194 channel=28
    -10, -9, 3, -1, -13, 0, -15, -11, -4,
    -- layer=1 filter=194 channel=29
    -1, -7, -1, -14, -7, -5, -14, -3, -4,
    -- layer=1 filter=194 channel=30
    -5, 3, 8, 11, 1, -7, -12, -15, -20,
    -- layer=1 filter=194 channel=31
    2, 12, -1, -1, 13, 9, 1, 3, -14,
    -- layer=1 filter=194 channel=32
    -5, 4, -10, -12, -1, 2, 2, -2, -13,
    -- layer=1 filter=194 channel=33
    5, 0, -7, -10, 3, -16, -6, -8, 0,
    -- layer=1 filter=194 channel=34
    -4, 7, -5, -1, -1, -8, -11, 8, 7,
    -- layer=1 filter=194 channel=35
    4, 0, -11, -11, 0, -9, -3, -3, -8,
    -- layer=1 filter=194 channel=36
    -3, -1, -11, 4, -1, 6, 2, -13, -6,
    -- layer=1 filter=194 channel=37
    -11, -8, 0, -21, -20, -8, 10, 8, -15,
    -- layer=1 filter=194 channel=38
    0, 4, 5, -3, 0, -3, -9, -7, -7,
    -- layer=1 filter=194 channel=39
    -1, 2, 1, 4, -10, 7, 6, 6, -11,
    -- layer=1 filter=194 channel=40
    4, -1, 11, 0, 5, -7, -7, 6, 7,
    -- layer=1 filter=194 channel=41
    0, 7, -8, -4, 2, 5, -4, -7, 1,
    -- layer=1 filter=194 channel=42
    -7, -6, -16, -1, 6, 12, -1, 6, 3,
    -- layer=1 filter=194 channel=43
    -13, 9, 3, -6, 3, -3, -7, 2, -17,
    -- layer=1 filter=194 channel=44
    -2, 1, -18, -6, -14, -1, -7, -13, -17,
    -- layer=1 filter=194 channel=45
    1, -6, -8, -9, 4, -1, 0, -13, -13,
    -- layer=1 filter=194 channel=46
    -3, -4, 3, -5, 3, 1, 0, -3, -10,
    -- layer=1 filter=194 channel=47
    -11, 4, 2, 5, -9, 0, 0, -2, -9,
    -- layer=1 filter=194 channel=48
    0, 0, 5, 1, -6, -11, -7, -9, -6,
    -- layer=1 filter=194 channel=49
    0, 2, 2, 4, 8, -4, -4, 6, 0,
    -- layer=1 filter=194 channel=50
    4, -2, -9, 7, -9, -5, -5, -7, 2,
    -- layer=1 filter=194 channel=51
    0, -3, -7, -5, 0, -6, -12, -3, -4,
    -- layer=1 filter=194 channel=52
    7, 6, -4, 6, -9, 6, 0, 1, -9,
    -- layer=1 filter=194 channel=53
    -5, -4, 0, 6, 0, -4, 0, 3, -2,
    -- layer=1 filter=194 channel=54
    -19, -14, -16, -9, -8, -10, -1, -15, 0,
    -- layer=1 filter=194 channel=55
    -10, -4, -2, -16, -9, -9, 3, 0, 5,
    -- layer=1 filter=194 channel=56
    -3, -1, -9, -1, 2, 1, 5, -1, 0,
    -- layer=1 filter=194 channel=57
    -18, -1, -4, -15, -4, -14, -9, -5, 8,
    -- layer=1 filter=194 channel=58
    0, -16, 6, -15, -20, -1, 6, -15, 3,
    -- layer=1 filter=194 channel=59
    -9, 0, 0, -3, 7, -6, 8, 0, 2,
    -- layer=1 filter=194 channel=60
    -4, 6, -9, -4, 1, 10, -9, 5, 11,
    -- layer=1 filter=194 channel=61
    0, -2, -5, 9, 5, -1, 1, 1, -6,
    -- layer=1 filter=194 channel=62
    -12, -8, -3, -20, -8, -14, -7, -8, -13,
    -- layer=1 filter=194 channel=63
    -8, -9, -12, -13, -9, -4, -2, -15, -8,
    -- layer=1 filter=194 channel=64
    3, 6, -2, 7, -9, -12, -10, 6, 3,
    -- layer=1 filter=194 channel=65
    -2, 6, -4, 1, -1, -4, -10, -11, -2,
    -- layer=1 filter=194 channel=66
    3, -16, -7, -4, -10, -8, -10, -5, -1,
    -- layer=1 filter=194 channel=67
    12, 6, 10, 16, 9, 8, 0, 0, 7,
    -- layer=1 filter=194 channel=68
    -12, -3, -4, 8, -4, -15, 3, -18, -5,
    -- layer=1 filter=194 channel=69
    -27, -8, -19, -9, -21, -21, -7, 3, -18,
    -- layer=1 filter=194 channel=70
    -7, -1, 9, -4, -10, -9, -2, 0, 2,
    -- layer=1 filter=194 channel=71
    10, -10, 1, 2, -3, 6, 4, 1, 3,
    -- layer=1 filter=194 channel=72
    -9, -5, 0, -12, 8, -9, -3, -11, 0,
    -- layer=1 filter=194 channel=73
    1, -11, -3, -2, -6, -10, -4, 6, -10,
    -- layer=1 filter=194 channel=74
    5, 7, 5, -6, 7, -5, 8, -1, 5,
    -- layer=1 filter=194 channel=75
    -6, 8, 14, 19, 17, 1, -11, -16, 3,
    -- layer=1 filter=194 channel=76
    -2, 3, -1, 6, -3, -6, -4, 2, -3,
    -- layer=1 filter=194 channel=77
    7, 7, -8, 2, -8, 2, 1, -11, 6,
    -- layer=1 filter=194 channel=78
    3, -2, 1, -11, 1, 5, -8, -6, 0,
    -- layer=1 filter=194 channel=79
    -7, -12, -20, -11, -7, -14, -20, -10, -23,
    -- layer=1 filter=194 channel=80
    -6, 3, 10, 0, 1, 12, -8, -2, 10,
    -- layer=1 filter=194 channel=81
    7, -6, -1, 1, -7, 2, -1, 1, -2,
    -- layer=1 filter=194 channel=82
    11, 7, -2, 3, -6, -6, 7, 9, 2,
    -- layer=1 filter=194 channel=83
    4, -9, 1, -6, -4, 7, -2, -5, -9,
    -- layer=1 filter=194 channel=84
    -6, -5, 3, -4, 5, -2, -10, -16, -27,
    -- layer=1 filter=194 channel=85
    -5, 4, 6, -13, -9, 3, -2, 9, -6,
    -- layer=1 filter=194 channel=86
    -5, 0, 3, -15, -10, -18, -9, -16, -4,
    -- layer=1 filter=194 channel=87
    6, 7, -9, 8, 6, -6, -5, -5, 6,
    -- layer=1 filter=194 channel=88
    9, -6, -5, 14, 6, 0, 12, 10, -4,
    -- layer=1 filter=194 channel=89
    0, 0, 3, 3, -2, -2, -6, -3, -2,
    -- layer=1 filter=194 channel=90
    3, -15, 2, -11, 2, -6, -3, -4, 2,
    -- layer=1 filter=194 channel=91
    2, -5, 3, -8, -16, 0, -11, -13, -16,
    -- layer=1 filter=194 channel=92
    5, 3, 2, -4, 1, -3, -5, -1, 5,
    -- layer=1 filter=194 channel=93
    -11, 1, -3, -10, 6, 7, 5, -6, 0,
    -- layer=1 filter=194 channel=94
    1, -2, -7, 1, -1, 0, 5, -8, 0,
    -- layer=1 filter=194 channel=95
    4, 8, -3, 6, -10, -13, -18, -8, -17,
    -- layer=1 filter=194 channel=96
    4, -5, 0, -1, 8, 3, 5, -2, -2,
    -- layer=1 filter=194 channel=97
    -2, -2, -14, -9, -8, -3, -6, -7, -12,
    -- layer=1 filter=194 channel=98
    -13, -6, -7, -16, -22, -19, -12, -11, -3,
    -- layer=1 filter=194 channel=99
    -2, -6, -2, -4, 4, -7, -9, -8, -3,
    -- layer=1 filter=194 channel=100
    -6, 4, -2, 0, 1, 3, 7, 6, 6,
    -- layer=1 filter=194 channel=101
    -14, 0, -9, -5, -6, -6, -7, -9, -2,
    -- layer=1 filter=194 channel=102
    3, 0, -7, 1, -9, -6, 2, -9, -3,
    -- layer=1 filter=194 channel=103
    -10, -13, -9, 0, -2, 4, -8, -9, 0,
    -- layer=1 filter=194 channel=104
    4, 1, 0, -4, -2, 5, -6, -8, -5,
    -- layer=1 filter=194 channel=105
    -3, -7, -13, 0, -10, 3, 2, 0, -10,
    -- layer=1 filter=194 channel=106
    -4, 5, -11, 7, 0, -19, -4, -20, -14,
    -- layer=1 filter=194 channel=107
    0, 9, 4, -10, 4, -7, -10, 6, 0,
    -- layer=1 filter=194 channel=108
    -2, 3, -8, -4, 2, 1, 2, -1, -7,
    -- layer=1 filter=194 channel=109
    3, -8, -11, 4, -2, 5, 8, 7, -3,
    -- layer=1 filter=194 channel=110
    0, 8, 4, -10, -3, 1, -1, 1, 0,
    -- layer=1 filter=194 channel=111
    -4, 3, 2, -6, -9, -1, -4, -16, -24,
    -- layer=1 filter=194 channel=112
    -8, -6, -2, 0, 6, -3, -4, 3, -2,
    -- layer=1 filter=194 channel=113
    -16, -15, -16, -6, 1, 3, -16, 1, -13,
    -- layer=1 filter=194 channel=114
    -17, -14, 0, -9, -8, -23, -2, -4, 0,
    -- layer=1 filter=194 channel=115
    -1, -2, -12, -6, -13, 1, -14, 0, -1,
    -- layer=1 filter=194 channel=116
    8, 1, 6, -10, 8, -2, 8, 7, -6,
    -- layer=1 filter=194 channel=117
    -8, -5, 11, -12, -18, -13, -21, -10, -18,
    -- layer=1 filter=194 channel=118
    -9, 4, -3, 0, -14, -1, -2, -9, -9,
    -- layer=1 filter=194 channel=119
    -4, -3, -3, -7, -11, -5, 6, -13, -18,
    -- layer=1 filter=194 channel=120
    -4, -1, -6, 3, 6, -8, -11, -9, -7,
    -- layer=1 filter=194 channel=121
    -6, -9, -6, 4, 10, 14, 4, 6, 0,
    -- layer=1 filter=194 channel=122
    -8, -2, 1, -4, 5, 8, -6, 8, 0,
    -- layer=1 filter=194 channel=123
    0, -14, -18, -2, -8, -1, -8, 4, -9,
    -- layer=1 filter=194 channel=124
    1, 9, 6, 4, 5, -4, 3, -2, -12,
    -- layer=1 filter=194 channel=125
    0, -3, 8, 8, -15, -7, -16, 0, -3,
    -- layer=1 filter=194 channel=126
    -6, -8, -5, 4, 8, -11, -7, -9, -2,
    -- layer=1 filter=194 channel=127
    1, 9, -1, 13, -3, -5, -12, -7, -8,
    -- layer=1 filter=195 channel=0
    -5, 3, -2, 13, 0, 1, 0, -4, -9,
    -- layer=1 filter=195 channel=1
    12, 15, -15, -28, -11, 19, -41, -2, 27,
    -- layer=1 filter=195 channel=2
    4, 5, 0, -12, 5, -12, -29, -16, -7,
    -- layer=1 filter=195 channel=3
    6, -11, 7, -5, 2, 2, 2, -2, 8,
    -- layer=1 filter=195 channel=4
    0, 3, 1, 13, 0, 7, 4, -2, 4,
    -- layer=1 filter=195 channel=5
    44, 16, -6, -9, 10, 16, -29, 10, 10,
    -- layer=1 filter=195 channel=6
    0, 51, 82, -94, -20, 21, -73, -34, 18,
    -- layer=1 filter=195 channel=7
    -36, 13, 12, -11, -20, 40, -1, 25, 45,
    -- layer=1 filter=195 channel=8
    41, 20, -18, 1, 18, 27, -19, 5, 19,
    -- layer=1 filter=195 channel=9
    -68, -31, 13, 33, -11, 23, -42, 0, -29,
    -- layer=1 filter=195 channel=10
    -13, 32, 35, -5, 1, 53, 9, 34, 42,
    -- layer=1 filter=195 channel=11
    28, 7, -5, 48, 32, -16, 42, 14, -3,
    -- layer=1 filter=195 channel=12
    0, 54, 0, -33, -38, -3, -39, -13, 7,
    -- layer=1 filter=195 channel=13
    -24, -26, 26, -78, -23, 9, -70, 2, 22,
    -- layer=1 filter=195 channel=14
    -72, 38, 4, 0, -36, 10, -20, -14, 12,
    -- layer=1 filter=195 channel=15
    4, -40, -44, -33, 1, -27, -79, -43, 22,
    -- layer=1 filter=195 channel=16
    30, -16, -34, -4, 8, 8, -16, 15, 10,
    -- layer=1 filter=195 channel=17
    -5, 0, 0, -19, -4, -7, -32, -11, -11,
    -- layer=1 filter=195 channel=18
    -11, -3, 8, 10, 18, 18, 16, -10, 10,
    -- layer=1 filter=195 channel=19
    -5, -30, 44, 23, 27, 28, -19, 27, -2,
    -- layer=1 filter=195 channel=20
    -43, -17, 14, -80, -34, 8, -89, -33, -6,
    -- layer=1 filter=195 channel=21
    -34, 8, 3, -51, -8, 35, -55, -25, 3,
    -- layer=1 filter=195 channel=22
    -30, -13, 8, -63, -25, 11, -34, -16, 14,
    -- layer=1 filter=195 channel=23
    -57, 17, 27, -46, 11, 33, 6, 17, 54,
    -- layer=1 filter=195 channel=24
    -6, -45, 4, -13, -2, 28, -3, 18, 13,
    -- layer=1 filter=195 channel=25
    -26, -22, -10, -15, -33, 33, -15, 15, 22,
    -- layer=1 filter=195 channel=26
    -30, -52, 2, -59, 28, -5, -8, 21, 29,
    -- layer=1 filter=195 channel=27
    7, -27, -42, 6, -21, -57, 29, -28, -35,
    -- layer=1 filter=195 channel=28
    -44, 3, 4, -13, -43, 26, -20, 25, 23,
    -- layer=1 filter=195 channel=29
    -62, -54, -66, -29, -48, -47, -14, -37, -41,
    -- layer=1 filter=195 channel=30
    -10, 7, 47, 3, 11, 34, -27, -15, 8,
    -- layer=1 filter=195 channel=31
    -31, 27, 35, -27, -16, 16, -60, -45, 5,
    -- layer=1 filter=195 channel=32
    -39, -46, 9, -49, 11, -10, -24, 4, 33,
    -- layer=1 filter=195 channel=33
    -11, -11, 2, -15, -15, 6, -4, -13, 6,
    -- layer=1 filter=195 channel=34
    -11, -4, 21, -7, 0, 17, -11, 27, -1,
    -- layer=1 filter=195 channel=35
    -8, -9, -1, -6, 1, -6, -7, -6, -2,
    -- layer=1 filter=195 channel=36
    33, 17, -8, 59, 16, -2, 47, 22, -13,
    -- layer=1 filter=195 channel=37
    32, 14, -29, -3, 14, 24, -8, 22, 24,
    -- layer=1 filter=195 channel=38
    -30, -10, 70, -64, -27, 52, -80, -27, 10,
    -- layer=1 filter=195 channel=39
    19, 10, -11, 12, 12, 2, -8, -7, -9,
    -- layer=1 filter=195 channel=40
    -74, 12, 44, -25, -16, 16, -35, -38, 17,
    -- layer=1 filter=195 channel=41
    -30, -25, 8, -8, 14, 0, 3, 27, -22,
    -- layer=1 filter=195 channel=42
    -26, 11, -2, -17, -2, -2, -40, -38, -21,
    -- layer=1 filter=195 channel=43
    16, -3, -28, -20, 4, 16, -26, 21, 17,
    -- layer=1 filter=195 channel=44
    -33, -42, 1, -37, 25, 23, -6, 33, 34,
    -- layer=1 filter=195 channel=45
    6, -30, -13, -46, -5, -13, -48, -23, 20,
    -- layer=1 filter=195 channel=46
    -23, 0, 57, -2, 19, 11, -68, -13, 10,
    -- layer=1 filter=195 channel=47
    -58, -6, 12, -58, -8, 8, -19, -8, 22,
    -- layer=1 filter=195 channel=48
    -13, -14, 31, -22, -6, 28, -22, -11, 28,
    -- layer=1 filter=195 channel=49
    -5, 6, -6, -16, -17, 2, -45, -41, -6,
    -- layer=1 filter=195 channel=50
    -22, -34, 10, 2, -7, 3, -16, -36, -13,
    -- layer=1 filter=195 channel=51
    -39, -7, 36, -41, -37, 24, -40, -7, 17,
    -- layer=1 filter=195 channel=52
    0, 5, -17, 8, -7, 15, 2, -11, 7,
    -- layer=1 filter=195 channel=53
    -2, -7, -5, 4, -9, 1, 5, -8, -14,
    -- layer=1 filter=195 channel=54
    -7, -23, -18, 10, 12, 37, -23, 58, 32,
    -- layer=1 filter=195 channel=55
    44, 3, -29, 36, 11, -13, 42, 13, -14,
    -- layer=1 filter=195 channel=56
    4, 7, -4, 7, -6, 1, -6, 9, 5,
    -- layer=1 filter=195 channel=57
    -57, -22, 29, -19, -53, 30, -22, -14, 18,
    -- layer=1 filter=195 channel=58
    -80, 25, 54, -24, 29, 59, 21, 13, 51,
    -- layer=1 filter=195 channel=59
    8, 18, 2, 8, -1, 4, -12, -7, -16,
    -- layer=1 filter=195 channel=60
    3, -8, 1, 12, -9, 11, 3, 5, 8,
    -- layer=1 filter=195 channel=61
    2, -6, 8, 11, 5, -6, -2, 5, -7,
    -- layer=1 filter=195 channel=62
    43, -1, -25, -15, 35, 23, -15, 17, 19,
    -- layer=1 filter=195 channel=63
    18, -2, -11, 42, 22, 3, 21, 11, -9,
    -- layer=1 filter=195 channel=64
    3, -2, 8, -18, -7, 5, -16, -6, -10,
    -- layer=1 filter=195 channel=65
    -26, 22, 34, -42, 4, 34, -32, -2, 5,
    -- layer=1 filter=195 channel=66
    11, 0, 0, 28, 0, -4, 0, 0, -17,
    -- layer=1 filter=195 channel=67
    4, -17, 46, -34, 8, 94, -66, -19, 25,
    -- layer=1 filter=195 channel=68
    -18, -35, 1, -37, 20, 7, 7, 17, 36,
    -- layer=1 filter=195 channel=69
    31, -27, -34, -17, -5, -11, -32, 1, 10,
    -- layer=1 filter=195 channel=70
    44, 106, 50, -53, -36, 46, -60, -37, 10,
    -- layer=1 filter=195 channel=71
    -6, 20, 15, -2, 3, 23, -13, 8, 12,
    -- layer=1 filter=195 channel=72
    -27, -3, 51, 11, 12, 5, -33, -6, 0,
    -- layer=1 filter=195 channel=73
    -6, 3, -5, -7, -5, 9, -7, 0, 7,
    -- layer=1 filter=195 channel=74
    -15, 9, 7, -16, 16, 20, -16, -25, 14,
    -- layer=1 filter=195 channel=75
    -12, 40, 53, -9, -2, 1, -24, 0, 8,
    -- layer=1 filter=195 channel=76
    -10, -13, 5, 0, 17, 0, 16, 6, 8,
    -- layer=1 filter=195 channel=77
    -35, -8, 18, -49, -19, 22, -16, 0, 4,
    -- layer=1 filter=195 channel=78
    1, -8, -14, 11, -12, -4, -3, 14, -14,
    -- layer=1 filter=195 channel=79
    24, -11, -20, -19, 4, 0, -36, -4, 4,
    -- layer=1 filter=195 channel=80
    4, -4, 7, 2, 1, -2, -5, -8, -4,
    -- layer=1 filter=195 channel=81
    0, -15, -13, -15, -14, 6, -7, 7, -9,
    -- layer=1 filter=195 channel=82
    -21, 3, 40, -66, -24, 53, -55, -28, 15,
    -- layer=1 filter=195 channel=83
    16, -8, -8, -48, 6, -16, -43, -29, 19,
    -- layer=1 filter=195 channel=84
    -16, -9, 16, -9, 27, 17, 21, 20, 37,
    -- layer=1 filter=195 channel=85
    -39, 20, 42, -46, 17, 48, 6, 31, 26,
    -- layer=1 filter=195 channel=86
    7, 6, -9, 26, -2, -14, 10, -8, -14,
    -- layer=1 filter=195 channel=87
    -70, 9, 71, 20, 4, 22, -60, 20, -15,
    -- layer=1 filter=195 channel=88
    -9, -14, 28, -17, -13, 21, -19, -28, 4,
    -- layer=1 filter=195 channel=89
    -48, -4, 33, -58, -4, 23, -31, -3, 33,
    -- layer=1 filter=195 channel=90
    -39, -68, -35, -41, -9, -14, -24, 0, 26,
    -- layer=1 filter=195 channel=91
    -38, -13, 22, -66, -50, 17, -75, -66, 0,
    -- layer=1 filter=195 channel=92
    26, -43, -51, -22, -18, -27, -13, -7, -5,
    -- layer=1 filter=195 channel=93
    -12, 6, 7, -13, 1, 18, -19, -6, 5,
    -- layer=1 filter=195 channel=94
    1, 21, 8, 22, 0, 0, -2, -6, -10,
    -- layer=1 filter=195 channel=95
    -21, -2, 20, 2, 31, 20, -4, 26, 28,
    -- layer=1 filter=195 channel=96
    -7, 0, 9, -7, 1, -2, 2, 12, -1,
    -- layer=1 filter=195 channel=97
    -2, 5, 1, 3, -9, -15, -5, -2, -11,
    -- layer=1 filter=195 channel=98
    31, -1, -13, -16, 13, 1, -37, 7, 8,
    -- layer=1 filter=195 channel=99
    -49, -32, -10, -18, -37, 35, 17, 48, 27,
    -- layer=1 filter=195 channel=100
    36, 5, -15, 26, 30, -12, 36, -6, -12,
    -- layer=1 filter=195 channel=101
    -56, 0, 31, -71, -16, 33, -64, -31, 8,
    -- layer=1 filter=195 channel=102
    -19, 11, 30, -7, -18, -2, -37, -22, -5,
    -- layer=1 filter=195 channel=103
    22, -11, -6, 38, 18, -9, 30, -8, -17,
    -- layer=1 filter=195 channel=104
    -53, 4, 24, -30, 1, 13, 0, 4, -2,
    -- layer=1 filter=195 channel=105
    -8, 12, -3, 23, -3, -8, 11, 5, -17,
    -- layer=1 filter=195 channel=106
    -45, -14, 34, -78, 5, 13, -71, 7, 15,
    -- layer=1 filter=195 channel=107
    -7, -9, -7, 0, 13, 0, 2, 4, 5,
    -- layer=1 filter=195 channel=108
    -24, -67, -12, -43, 12, 23, -18, 7, 30,
    -- layer=1 filter=195 channel=109
    0, -4, -3, 5, -1, -8, -9, 3, -7,
    -- layer=1 filter=195 channel=110
    -11, 2, 12, -3, 5, -13, -15, -11, 0,
    -- layer=1 filter=195 channel=111
    -5, -4, 11, -15, 19, 4, 6, 6, 22,
    -- layer=1 filter=195 channel=112
    1, -21, -7, -11, 17, 18, 1, 8, 29,
    -- layer=1 filter=195 channel=113
    -49, -2, 17, -42, -29, 15, -68, -49, -8,
    -- layer=1 filter=195 channel=114
    21, -5, -54, 11, 12, -22, -17, 0, -11,
    -- layer=1 filter=195 channel=115
    17, 19, 2, 13, 0, 11, 0, -1, -12,
    -- layer=1 filter=195 channel=116
    -7, -5, 7, 0, 0, 5, 5, 3, 5,
    -- layer=1 filter=195 channel=117
    14, -11, 7, -14, -4, 8, 30, 23, 23,
    -- layer=1 filter=195 channel=118
    -15, 0, 27, -1, 22, 25, -18, 11, 15,
    -- layer=1 filter=195 channel=119
    -25, -53, -1, -52, 0, 10, 0, 10, 41,
    -- layer=1 filter=195 channel=120
    -32, -2, 9, -26, -11, 18, -18, -13, -4,
    -- layer=1 filter=195 channel=121
    -3, 14, -9, 11, -8, -15, -5, -3, -12,
    -- layer=1 filter=195 channel=122
    2, 10, -4, 2, -7, -2, 0, -6, -4,
    -- layer=1 filter=195 channel=123
    15, 5, -27, 43, 25, -15, 37, 0, -12,
    -- layer=1 filter=195 channel=124
    -7, 9, 2, 0, 2, 0, 7, -8, 5,
    -- layer=1 filter=195 channel=125
    43, 70, 89, -71, -21, 15, -70, -48, -7,
    -- layer=1 filter=195 channel=126
    42, 30, 0, -15, 14, 32, -6, 13, 2,
    -- layer=1 filter=195 channel=127
    -13, 11, 35, 1, 15, 6, -9, -3, 8,
    -- layer=1 filter=196 channel=0
    -4, -5, -7, -1, -1, -8, 5, -11, -12,
    -- layer=1 filter=196 channel=1
    2, 2, -7, 6, -5, -5, 0, 0, 6,
    -- layer=1 filter=196 channel=2
    -11, 3, -9, -10, -9, 7, -3, 8, -11,
    -- layer=1 filter=196 channel=3
    10, 0, -2, 7, -10, 4, 7, 3, 1,
    -- layer=1 filter=196 channel=4
    2, 0, -5, -3, 2, -12, 2, -5, -2,
    -- layer=1 filter=196 channel=5
    8, -4, -6, -5, 5, 5, -2, -7, -3,
    -- layer=1 filter=196 channel=6
    -11, 1, -7, 5, 3, -7, 5, -10, -7,
    -- layer=1 filter=196 channel=7
    -1, -4, 2, -3, 7, 3, 7, -1, 0,
    -- layer=1 filter=196 channel=8
    -4, 5, -8, -1, 8, 0, -7, -3, -11,
    -- layer=1 filter=196 channel=9
    1, -9, 3, 0, -4, -1, -10, -1, 5,
    -- layer=1 filter=196 channel=10
    9, 0, 2, 5, -8, 0, -7, 4, -9,
    -- layer=1 filter=196 channel=11
    -6, -7, 0, 1, 3, -4, 2, 5, -9,
    -- layer=1 filter=196 channel=12
    0, -6, 1, -9, 3, -6, 1, 3, 7,
    -- layer=1 filter=196 channel=13
    -2, -10, 0, -7, -8, 1, -5, -7, 9,
    -- layer=1 filter=196 channel=14
    -4, -12, 2, -2, -9, 2, -6, 4, 0,
    -- layer=1 filter=196 channel=15
    -12, 3, -10, 6, -9, 3, -9, 0, 2,
    -- layer=1 filter=196 channel=16
    0, -10, -9, -11, -4, -5, -4, -12, 0,
    -- layer=1 filter=196 channel=17
    3, 0, -3, -4, 7, -5, -4, 3, 6,
    -- layer=1 filter=196 channel=18
    1, -2, 7, -3, -13, 0, 0, -2, -7,
    -- layer=1 filter=196 channel=19
    2, 2, -3, 5, 2, 5, -1, -8, 0,
    -- layer=1 filter=196 channel=20
    3, 0, -1, 6, 7, -9, -10, 0, -12,
    -- layer=1 filter=196 channel=21
    8, -2, 3, -4, 7, 3, 8, 2, 6,
    -- layer=1 filter=196 channel=22
    4, 4, 8, 6, 7, 9, 3, 8, 8,
    -- layer=1 filter=196 channel=23
    0, 2, 7, 4, -5, -8, 4, 2, -4,
    -- layer=1 filter=196 channel=24
    8, -3, 0, -3, -10, -10, 4, 7, -8,
    -- layer=1 filter=196 channel=25
    8, 0, 0, -3, 0, -11, -4, 1, 3,
    -- layer=1 filter=196 channel=26
    -3, -2, -3, 0, 6, 6, -7, 7, 10,
    -- layer=1 filter=196 channel=27
    -2, 6, -7, -6, -9, -8, -3, -8, 9,
    -- layer=1 filter=196 channel=28
    0, -5, -9, -5, -1, -12, -8, 7, 1,
    -- layer=1 filter=196 channel=29
    -1, 7, -1, -1, -1, 7, -4, -8, -8,
    -- layer=1 filter=196 channel=30
    -6, -2, -6, 1, -4, 0, 4, -1, 4,
    -- layer=1 filter=196 channel=31
    -8, -3, -4, 4, -1, -7, 8, 7, 9,
    -- layer=1 filter=196 channel=32
    3, 0, 6, 7, -7, 2, -2, -5, -4,
    -- layer=1 filter=196 channel=33
    1, -9, 6, 3, -8, 0, 6, -9, 6,
    -- layer=1 filter=196 channel=34
    -9, 8, 1, 0, -7, 2, 4, 2, 1,
    -- layer=1 filter=196 channel=35
    -1, -10, -6, -9, 7, -2, 3, 5, 7,
    -- layer=1 filter=196 channel=36
    5, -6, -3, -3, -3, -13, -5, -2, 6,
    -- layer=1 filter=196 channel=37
    3, 3, 0, 5, -6, -5, -2, -11, -6,
    -- layer=1 filter=196 channel=38
    -4, -7, -9, 8, 2, 5, 9, 5, -8,
    -- layer=1 filter=196 channel=39
    -8, 7, 8, -8, -3, 8, -1, 1, 0,
    -- layer=1 filter=196 channel=40
    5, 5, -13, 4, 3, -2, 9, 1, -7,
    -- layer=1 filter=196 channel=41
    8, -1, 6, -6, -6, 1, 0, 0, 4,
    -- layer=1 filter=196 channel=42
    -11, -12, -10, 4, -14, -7, 5, 0, -2,
    -- layer=1 filter=196 channel=43
    1, -3, -6, 7, 8, 0, 4, 0, 8,
    -- layer=1 filter=196 channel=44
    -5, 3, -11, -1, 6, -7, 8, -7, 3,
    -- layer=1 filter=196 channel=45
    0, 7, -3, 0, 6, -1, -9, -5, 6,
    -- layer=1 filter=196 channel=46
    -5, -7, -2, -1, -8, -7, -4, -3, 6,
    -- layer=1 filter=196 channel=47
    -11, 3, 8, -8, 6, -9, 7, -3, 6,
    -- layer=1 filter=196 channel=48
    6, 7, 7, 3, 6, 2, -10, -5, 3,
    -- layer=1 filter=196 channel=49
    1, 0, -8, 5, 3, -12, -11, -2, -7,
    -- layer=1 filter=196 channel=50
    2, -7, 3, -9, 7, 3, 2, 3, -5,
    -- layer=1 filter=196 channel=51
    -3, -10, 2, -4, 0, 2, 5, -6, 1,
    -- layer=1 filter=196 channel=52
    7, 0, 0, 2, -4, 4, -4, -1, -7,
    -- layer=1 filter=196 channel=53
    4, -4, 4, -5, 3, 2, -5, -2, -1,
    -- layer=1 filter=196 channel=54
    -3, 0, -12, -4, -11, 0, -13, -11, -9,
    -- layer=1 filter=196 channel=55
    -2, -9, 4, 8, 0, -11, 3, -7, 0,
    -- layer=1 filter=196 channel=56
    -6, 2, 4, -8, -7, 6, 2, 8, 6,
    -- layer=1 filter=196 channel=57
    -10, 1, -8, -9, 6, -5, 4, 1, -3,
    -- layer=1 filter=196 channel=58
    0, 9, -10, 1, -12, 0, -7, -10, 0,
    -- layer=1 filter=196 channel=59
    5, -4, -11, 0, 0, 0, 2, -4, 1,
    -- layer=1 filter=196 channel=60
    -10, 8, 6, -7, -5, 7, -1, -7, 6,
    -- layer=1 filter=196 channel=61
    3, -6, 7, 8, 0, 5, 7, 9, -3,
    -- layer=1 filter=196 channel=62
    -7, 2, -8, -7, 3, 6, 2, -5, 1,
    -- layer=1 filter=196 channel=63
    0, -4, -2, 0, 5, 4, 6, 0, 1,
    -- layer=1 filter=196 channel=64
    -9, 5, 3, 0, -1, -5, 1, -12, -5,
    -- layer=1 filter=196 channel=65
    -3, -8, 6, 0, -11, 2, -11, -2, -7,
    -- layer=1 filter=196 channel=66
    -9, 4, -7, -1, 2, 7, -4, -7, 5,
    -- layer=1 filter=196 channel=67
    -1, -7, 6, -7, 1, -10, 7, 0, 4,
    -- layer=1 filter=196 channel=68
    7, 0, 0, 6, -1, 9, 1, 0, 0,
    -- layer=1 filter=196 channel=69
    -8, 5, -2, -2, -5, -1, 7, 0, -9,
    -- layer=1 filter=196 channel=70
    8, 2, -11, -9, 2, 0, 0, -10, 9,
    -- layer=1 filter=196 channel=71
    1, 5, -3, -12, 0, 6, -12, -10, -12,
    -- layer=1 filter=196 channel=72
    -11, -10, -1, -12, -11, 3, 0, -1, -5,
    -- layer=1 filter=196 channel=73
    -7, -12, 0, -9, 3, -9, -12, -8, 6,
    -- layer=1 filter=196 channel=74
    3, -4, -1, 6, 2, 3, 0, 5, 4,
    -- layer=1 filter=196 channel=75
    -9, -8, -11, 3, -4, -7, -9, 7, 6,
    -- layer=1 filter=196 channel=76
    1, 0, 1, -2, 7, 0, -8, 1, -7,
    -- layer=1 filter=196 channel=77
    2, 5, -9, 2, -11, 6, 6, 6, -7,
    -- layer=1 filter=196 channel=78
    -4, -9, 5, 7, -3, -1, -2, 1, -8,
    -- layer=1 filter=196 channel=79
    0, -9, 6, -8, -2, 8, -12, 1, -6,
    -- layer=1 filter=196 channel=80
    2, 6, -5, 2, 4, -4, 0, 7, 0,
    -- layer=1 filter=196 channel=81
    4, -6, -11, -7, -8, -12, 4, -7, -1,
    -- layer=1 filter=196 channel=82
    -4, 8, -7, 2, 5, 7, 7, 2, 6,
    -- layer=1 filter=196 channel=83
    4, -9, 0, 5, -5, 2, -10, -11, -1,
    -- layer=1 filter=196 channel=84
    -1, 0, 0, -8, -2, 5, 0, -1, 2,
    -- layer=1 filter=196 channel=85
    -3, -4, -6, 2, 4, 5, 2, 6, 7,
    -- layer=1 filter=196 channel=86
    1, -9, 6, -8, 3, -13, -10, -10, -2,
    -- layer=1 filter=196 channel=87
    2, 4, -10, -11, -10, -2, 8, -5, -11,
    -- layer=1 filter=196 channel=88
    -4, -7, -3, 8, -9, 4, 9, -3, 0,
    -- layer=1 filter=196 channel=89
    -5, -11, 8, 5, -7, 8, -1, 3, -12,
    -- layer=1 filter=196 channel=90
    4, 6, 0, -2, 3, -10, 2, -10, -8,
    -- layer=1 filter=196 channel=91
    -2, 4, 0, -3, -10, 0, -5, 8, -9,
    -- layer=1 filter=196 channel=92
    1, -10, 5, -2, 2, -6, -5, -1, -1,
    -- layer=1 filter=196 channel=93
    7, 7, 0, 2, 0, 0, -3, -6, -9,
    -- layer=1 filter=196 channel=94
    -2, 0, -8, 1, -11, 0, -2, 4, -10,
    -- layer=1 filter=196 channel=95
    -8, 0, 0, 5, -3, -8, -3, 0, -5,
    -- layer=1 filter=196 channel=96
    -3, 0, -5, 5, 0, -11, -8, 7, -12,
    -- layer=1 filter=196 channel=97
    0, -5, 2, 6, -10, -11, 6, 1, -9,
    -- layer=1 filter=196 channel=98
    -11, -5, 2, 2, -1, -11, -4, -10, -4,
    -- layer=1 filter=196 channel=99
    -8, -12, 8, 7, -4, 2, 5, 6, 2,
    -- layer=1 filter=196 channel=100
    -2, -3, 5, -4, -2, 5, 4, -4, 5,
    -- layer=1 filter=196 channel=101
    -11, -10, 0, 8, 6, -9, -10, -4, -6,
    -- layer=1 filter=196 channel=102
    4, 7, -12, 5, -6, 0, -8, -8, 8,
    -- layer=1 filter=196 channel=103
    -3, -4, -9, -7, 7, -8, -10, -5, 4,
    -- layer=1 filter=196 channel=104
    -9, 8, -9, -11, -8, 7, 6, -4, -5,
    -- layer=1 filter=196 channel=105
    -11, 8, 8, 6, -1, -8, -3, 0, 3,
    -- layer=1 filter=196 channel=106
    -3, 3, 6, -11, -6, 1, -9, 5, -7,
    -- layer=1 filter=196 channel=107
    0, 7, -8, 7, 0, -6, 6, -11, 0,
    -- layer=1 filter=196 channel=108
    6, 0, -1, -8, -8, 0, 0, -10, -5,
    -- layer=1 filter=196 channel=109
    9, -4, -3, -3, -8, -8, 8, 0, 3,
    -- layer=1 filter=196 channel=110
    1, 0, -12, 6, 0, -2, 4, -4, 4,
    -- layer=1 filter=196 channel=111
    0, 6, -5, 0, -6, -9, 3, -7, 6,
    -- layer=1 filter=196 channel=112
    -4, 0, -5, 5, 0, -11, -7, 3, 1,
    -- layer=1 filter=196 channel=113
    6, -1, 5, 6, 1, 3, -9, -6, 9,
    -- layer=1 filter=196 channel=114
    -6, 5, -9, -2, 3, 7, 0, -9, 4,
    -- layer=1 filter=196 channel=115
    -12, -4, -5, -9, 4, -2, -10, 3, -6,
    -- layer=1 filter=196 channel=116
    6, 4, 9, 9, 0, 0, -1, -9, 5,
    -- layer=1 filter=196 channel=117
    -8, 3, -12, 6, 1, -3, 0, -12, 4,
    -- layer=1 filter=196 channel=118
    -1, -3, -7, -5, 3, -8, 1, -11, 4,
    -- layer=1 filter=196 channel=119
    -1, -11, 3, 1, 5, -3, -1, -5, -5,
    -- layer=1 filter=196 channel=120
    -5, -9, -10, -9, 0, 3, -1, -2, 7,
    -- layer=1 filter=196 channel=121
    4, -7, -5, -1, -8, -7, -7, 4, -8,
    -- layer=1 filter=196 channel=122
    0, 7, 1, 8, 0, -5, -10, -10, -8,
    -- layer=1 filter=196 channel=123
    4, -8, 4, -6, -3, 6, 0, -10, 2,
    -- layer=1 filter=196 channel=124
    -11, -10, -4, 8, 2, -10, -7, -5, -3,
    -- layer=1 filter=196 channel=125
    4, 0, -4, 8, -9, -5, 4, 0, -10,
    -- layer=1 filter=196 channel=126
    7, -1, 9, -5, 8, 0, -6, 9, 8,
    -- layer=1 filter=196 channel=127
    -7, 0, 0, -8, -8, -4, -12, -9, 0,
    -- layer=1 filter=197 channel=0
    4, -3, -6, 4, -5, -11, 5, -2, -5,
    -- layer=1 filter=197 channel=1
    13, -4, -24, 24, 9, -8, 6, 15, -5,
    -- layer=1 filter=197 channel=2
    -1, 4, 12, -5, 17, 11, 17, 12, 18,
    -- layer=1 filter=197 channel=3
    7, -11, 9, 3, -7, -8, 6, 0, -11,
    -- layer=1 filter=197 channel=4
    18, 7, 15, -3, -8, -10, -7, -8, -9,
    -- layer=1 filter=197 channel=5
    39, 19, 17, 20, 8, -5, -20, 6, -27,
    -- layer=1 filter=197 channel=6
    -19, -44, -29, -78, -59, -56, -28, -6, -5,
    -- layer=1 filter=197 channel=7
    35, 13, 24, -28, -38, -41, -53, -47, -96,
    -- layer=1 filter=197 channel=8
    19, -1, 9, 46, 26, 26, 31, 38, 17,
    -- layer=1 filter=197 channel=9
    9, 7, 50, 6, 11, 6, -12, 17, -1,
    -- layer=1 filter=197 channel=10
    34, 31, 9, -31, -23, -44, -20, -71, -100,
    -- layer=1 filter=197 channel=11
    9, 29, 18, -6, -1, 1, -27, -28, -3,
    -- layer=1 filter=197 channel=12
    -12, -50, 10, -40, -16, -37, -39, -12, -54,
    -- layer=1 filter=197 channel=13
    -31, -17, -23, -23, -33, -10, 27, 26, 50,
    -- layer=1 filter=197 channel=14
    66, 28, 29, -15, 0, -4, -60, -51, -59,
    -- layer=1 filter=197 channel=15
    38, 22, 3, 38, -16, 7, -46, 3, -12,
    -- layer=1 filter=197 channel=16
    35, 37, 32, 27, 24, 22, 34, 51, 8,
    -- layer=1 filter=197 channel=17
    -34, -22, -13, -7, -11, -2, 27, 1, 5,
    -- layer=1 filter=197 channel=18
    13, -6, 13, -3, 0, 7, -49, -44, -33,
    -- layer=1 filter=197 channel=19
    41, 65, 65, 85, 83, 85, 76, 37, 37,
    -- layer=1 filter=197 channel=20
    -33, -22, -35, -19, -17, -5, 36, 51, 42,
    -- layer=1 filter=197 channel=21
    -8, -30, -19, 7, -1, 2, 37, 44, 41,
    -- layer=1 filter=197 channel=22
    -50, -42, -35, 5, -14, 11, 47, 59, 38,
    -- layer=1 filter=197 channel=23
    50, 27, 29, 16, -20, -33, -58, -71, -64,
    -- layer=1 filter=197 channel=24
    2, -12, -3, -6, -4, 18, 30, 18, 27,
    -- layer=1 filter=197 channel=25
    25, 35, 31, 4, 15, 3, 3, 23, -20,
    -- layer=1 filter=197 channel=26
    -4, 36, 9, 0, -9, -25, -26, -11, 10,
    -- layer=1 filter=197 channel=27
    13, -4, -1, -20, -23, -31, -15, 6, -4,
    -- layer=1 filter=197 channel=28
    41, 23, 22, -6, -8, -26, 0, 1, -30,
    -- layer=1 filter=197 channel=29
    7, 6, 5, -7, -6, -16, 17, 34, 13,
    -- layer=1 filter=197 channel=30
    7, 0, 1, 20, 30, 16, -4, -15, -31,
    -- layer=1 filter=197 channel=31
    -21, -46, -21, -49, -41, -40, -64, -55, -62,
    -- layer=1 filter=197 channel=32
    19, 41, 46, -25, -32, -36, -87, -114, -39,
    -- layer=1 filter=197 channel=33
    -36, -17, -19, -23, -9, -9, -15, -10, -7,
    -- layer=1 filter=197 channel=34
    -4, -13, 0, -1, -27, -26, -28, -24, -3,
    -- layer=1 filter=197 channel=35
    16, 14, 9, 24, 3, 5, 31, 19, 29,
    -- layer=1 filter=197 channel=36
    -8, 9, 7, -19, 8, -5, -39, -25, -17,
    -- layer=1 filter=197 channel=37
    38, 12, 29, 24, 13, 16, -4, 1, -22,
    -- layer=1 filter=197 channel=38
    -30, -35, -34, -20, -28, -19, 33, 42, 34,
    -- layer=1 filter=197 channel=39
    5, 3, 2, 0, 0, 4, -17, 8, -1,
    -- layer=1 filter=197 channel=40
    -11, -28, -18, -46, -29, -47, -12, -36, -19,
    -- layer=1 filter=197 channel=41
    19, 28, 35, -25, 14, -14, -49, -68, 6,
    -- layer=1 filter=197 channel=42
    -6, -7, 0, 4, 24, 7, 6, 23, 5,
    -- layer=1 filter=197 channel=43
    14, 31, 0, 37, 18, 17, 18, 52, -5,
    -- layer=1 filter=197 channel=44
    -7, 38, 0, -20, -66, -47, -68, -64, -15,
    -- layer=1 filter=197 channel=45
    -5, -21, -10, 4, -19, -2, 3, 28, 27,
    -- layer=1 filter=197 channel=46
    35, 49, 23, 39, 49, 34, 74, 35, 16,
    -- layer=1 filter=197 channel=47
    60, -12, 16, -18, -25, -64, -101, -107, -58,
    -- layer=1 filter=197 channel=48
    -20, -27, -31, -14, -12, 0, 38, 28, 44,
    -- layer=1 filter=197 channel=49
    9, -23, -12, -23, -14, -11, 0, 0, 15,
    -- layer=1 filter=197 channel=50
    -9, -29, -2, 2, -13, -8, 11, -2, 4,
    -- layer=1 filter=197 channel=51
    2, 0, -13, -16, -19, -15, 18, 21, 9,
    -- layer=1 filter=197 channel=52
    12, 7, 14, 12, 12, 21, 0, 10, -9,
    -- layer=1 filter=197 channel=53
    4, 31, 0, 5, 22, 19, 10, 8, 10,
    -- layer=1 filter=197 channel=54
    31, 33, 41, 2, 11, 9, 31, 0, -24,
    -- layer=1 filter=197 channel=55
    26, 34, 16, 9, 10, -2, -32, -9, -22,
    -- layer=1 filter=197 channel=56
    -1, -14, 6, 0, -2, -4, 2, -10, -4,
    -- layer=1 filter=197 channel=57
    -6, 0, -3, -49, -33, -38, -25, -46, -47,
    -- layer=1 filter=197 channel=58
    44, -3, 33, -30, -51, -56, -40, -117, -95,
    -- layer=1 filter=197 channel=59
    1, -8, -20, 2, 3, 2, 9, 2, -8,
    -- layer=1 filter=197 channel=60
    15, 9, 0, 20, 0, 15, 4, 9, -6,
    -- layer=1 filter=197 channel=61
    -7, -9, -10, 7, 1, 0, 0, 3, -2,
    -- layer=1 filter=197 channel=62
    23, 33, 27, 35, 38, 39, 35, 50, 4,
    -- layer=1 filter=197 channel=63
    16, 5, 5, 4, -2, 4, -32, -22, -23,
    -- layer=1 filter=197 channel=64
    -7, 0, -15, 0, 5, -10, 11, 31, 21,
    -- layer=1 filter=197 channel=65
    -32, -27, -37, -1, -1, 0, 37, 29, 39,
    -- layer=1 filter=197 channel=66
    4, -2, -4, -1, -16, 0, -13, -24, -10,
    -- layer=1 filter=197 channel=67
    -39, -20, -36, -63, -39, -31, -37, 4, 13,
    -- layer=1 filter=197 channel=68
    -8, 31, 35, -27, -68, -29, -98, -69, -15,
    -- layer=1 filter=197 channel=69
    39, 26, 11, 27, 12, 0, -2, 29, -3,
    -- layer=1 filter=197 channel=70
    46, 11, 0, -23, -36, -28, -37, -66, -34,
    -- layer=1 filter=197 channel=71
    -8, -14, -19, 12, 11, 10, 7, 16, 2,
    -- layer=1 filter=197 channel=72
    -16, -9, 12, 3, 29, 17, 36, -21, -2,
    -- layer=1 filter=197 channel=73
    -10, -6, -4, 5, 9, -5, -11, 0, -8,
    -- layer=1 filter=197 channel=74
    -4, -3, 25, -43, -29, -10, -74, -70, -36,
    -- layer=1 filter=197 channel=75
    13, -60, -15, 1, 9, 38, -44, -10, -36,
    -- layer=1 filter=197 channel=76
    -6, 9, 6, -9, 0, -2, -35, -12, -3,
    -- layer=1 filter=197 channel=77
    -19, -30, -35, -9, -15, 3, 15, 29, 27,
    -- layer=1 filter=197 channel=78
    -3, -12, -3, -11, -23, -8, -11, -16, -17,
    -- layer=1 filter=197 channel=79
    15, 17, 17, 31, 16, 31, 31, 48, 24,
    -- layer=1 filter=197 channel=80
    15, 6, 7, -2, 4, 6, 21, 2, 10,
    -- layer=1 filter=197 channel=81
    -25, -15, -22, -2, -8, 8, 25, 19, 18,
    -- layer=1 filter=197 channel=82
    -21, -37, -30, -10, -13, -2, 34, 41, 40,
    -- layer=1 filter=197 channel=83
    1, -11, -7, 23, -23, -8, -23, 9, 8,
    -- layer=1 filter=197 channel=84
    10, 21, 33, 12, 28, 24, -48, -33, -12,
    -- layer=1 filter=197 channel=85
    30, 3, 21, 19, 4, -27, -61, -123, -65,
    -- layer=1 filter=197 channel=86
    1, -5, 18, -21, -11, 7, -9, -15, 3,
    -- layer=1 filter=197 channel=87
    12, 23, 22, 18, 36, 24, 70, 17, 10,
    -- layer=1 filter=197 channel=88
    -20, -10, -20, -3, 8, 0, 33, 37, 29,
    -- layer=1 filter=197 channel=89
    -21, -11, -25, -5, -14, -3, 33, 23, 47,
    -- layer=1 filter=197 channel=90
    10, 31, 15, -2, -49, -35, -64, -51, -15,
    -- layer=1 filter=197 channel=91
    -10, -32, -13, -13, -16, -19, 24, 22, 30,
    -- layer=1 filter=197 channel=92
    -26, 33, 21, -23, -51, 1, -23, -15, 5,
    -- layer=1 filter=197 channel=93
    -26, -22, -24, -1, -3, -6, 22, 24, 28,
    -- layer=1 filter=197 channel=94
    -10, 4, 4, -21, -17, -7, -15, -4, -5,
    -- layer=1 filter=197 channel=95
    11, 5, 14, 4, 39, 25, -61, -33, -3,
    -- layer=1 filter=197 channel=96
    6, 5, 10, -10, -6, -16, -17, -24, -8,
    -- layer=1 filter=197 channel=97
    -19, -12, -7, -10, 0, -2, 8, 20, 1,
    -- layer=1 filter=197 channel=98
    -17, 1, -2, 31, 16, 23, 40, 39, 19,
    -- layer=1 filter=197 channel=99
    54, 32, 3, -47, -49, -55, -56, -78, -103,
    -- layer=1 filter=197 channel=100
    -3, 10, 23, -31, -8, -10, -30, -27, 0,
    -- layer=1 filter=197 channel=101
    -35, -23, -17, -17, -13, -16, 30, 17, 28,
    -- layer=1 filter=197 channel=102
    -33, -13, 8, -28, -25, -12, -3, 12, 17,
    -- layer=1 filter=197 channel=103
    7, 5, 17, 10, -7, -10, -24, -12, -18,
    -- layer=1 filter=197 channel=104
    39, -12, 26, 4, -13, -27, -84, -47, -36,
    -- layer=1 filter=197 channel=105
    -12, 4, -6, -19, -3, -4, -14, 1, -10,
    -- layer=1 filter=197 channel=106
    -14, 1, -7, -30, -32, -40, 6, 2, 38,
    -- layer=1 filter=197 channel=107
    -38, -19, -21, -11, -10, -9, -9, -17, -12,
    -- layer=1 filter=197 channel=108
    7, 15, 8, -27, -27, -30, -44, -53, -9,
    -- layer=1 filter=197 channel=109
    6, -13, 7, -8, -3, 3, -1, 6, -2,
    -- layer=1 filter=197 channel=110
    8, -1, 6, -3, -11, 6, 7, 0, -1,
    -- layer=1 filter=197 channel=111
    12, 8, 10, 9, 34, 27, -22, -50, -10,
    -- layer=1 filter=197 channel=112
    6, 42, 17, 28, 17, 44, -63, -3, -3,
    -- layer=1 filter=197 channel=113
    -23, -14, -13, -13, -20, -3, 14, -8, 16,
    -- layer=1 filter=197 channel=114
    58, 42, 26, 53, 30, 12, -15, 9, 6,
    -- layer=1 filter=197 channel=115
    -4, 4, 3, -17, -19, -11, -10, -8, -10,
    -- layer=1 filter=197 channel=116
    7, 9, -11, 6, 8, 7, -9, -3, 7,
    -- layer=1 filter=197 channel=117
    54, 49, 36, 56, 39, 57, -7, -16, 18,
    -- layer=1 filter=197 channel=118
    3, 3, 20, 10, 23, 5, -44, -45, -8,
    -- layer=1 filter=197 channel=119
    13, 37, 32, -8, -25, -46, -73, -82, -51,
    -- layer=1 filter=197 channel=120
    1, -15, -22, -13, -2, -12, 41, 46, 31,
    -- layer=1 filter=197 channel=121
    35, 13, 5, 22, 32, 8, 21, 5, -30,
    -- layer=1 filter=197 channel=122
    3, -6, -8, -2, -8, 9, 2, 5, 10,
    -- layer=1 filter=197 channel=123
    10, 1, 7, 9, 15, 10, -8, -20, -27,
    -- layer=1 filter=197 channel=124
    6, 6, -8, 8, 5, 2, 11, 12, -1,
    -- layer=1 filter=197 channel=125
    35, 41, 13, -12, -32, -45, -19, -58, -39,
    -- layer=1 filter=197 channel=126
    -14, -12, -12, 52, 21, 24, 29, 47, 7,
    -- layer=1 filter=197 channel=127
    0, 9, 18, 11, 37, 19, -50, -38, -20,
    -- layer=1 filter=198 channel=0
    -9, -2, 1, 6, -3, 4, 0, 4, -6,
    -- layer=1 filter=198 channel=1
    -10, -3, -14, 0, 2, 5, -4, -3, -11,
    -- layer=1 filter=198 channel=2
    0, 3, -6, -9, 0, -11, 9, -5, 10,
    -- layer=1 filter=198 channel=3
    6, 0, -1, -8, 0, 0, -4, 2, 2,
    -- layer=1 filter=198 channel=4
    -9, -4, 2, -3, 0, 8, 0, 0, -9,
    -- layer=1 filter=198 channel=5
    8, 11, -14, -8, 1, -5, -8, -1, -8,
    -- layer=1 filter=198 channel=6
    -8, 9, 0, -5, 0, 5, -8, 5, -1,
    -- layer=1 filter=198 channel=7
    -9, -13, -8, 12, -6, -11, -14, -2, 8,
    -- layer=1 filter=198 channel=8
    4, -5, -3, -6, 1, -11, -5, 0, 6,
    -- layer=1 filter=198 channel=9
    0, -2, -3, 0, -3, -8, 0, 12, -11,
    -- layer=1 filter=198 channel=10
    -6, -5, -7, 10, -13, 3, -5, -7, -1,
    -- layer=1 filter=198 channel=11
    -3, -16, -17, -16, -7, -4, -16, 3, -18,
    -- layer=1 filter=198 channel=12
    1, 9, -14, 0, -14, 5, 5, 3, 1,
    -- layer=1 filter=198 channel=13
    -4, -13, -3, -12, -12, -5, -6, 2, -11,
    -- layer=1 filter=198 channel=14
    -2, -6, -9, 0, -12, -2, -1, 4, -10,
    -- layer=1 filter=198 channel=15
    -10, 14, -1, 0, 3, -2, 0, -12, 5,
    -- layer=1 filter=198 channel=16
    4, 8, -12, -14, 0, -14, -11, -1, 5,
    -- layer=1 filter=198 channel=17
    -15, -15, 6, -2, 5, -14, 5, -14, -10,
    -- layer=1 filter=198 channel=18
    -12, -15, -11, -8, -14, -6, -1, 4, 8,
    -- layer=1 filter=198 channel=19
    6, -8, 2, -9, -4, 3, 4, 7, -10,
    -- layer=1 filter=198 channel=20
    -9, -8, -11, 4, -17, -8, -12, 1, -2,
    -- layer=1 filter=198 channel=21
    4, 5, -9, -9, -9, -4, -7, -18, -6,
    -- layer=1 filter=198 channel=22
    -1, -2, -11, -4, -7, 0, -8, -12, -1,
    -- layer=1 filter=198 channel=23
    -1, -9, 6, 8, -8, -14, 0, -5, 0,
    -- layer=1 filter=198 channel=24
    -4, -4, -12, -1, -2, 1, -17, -14, -12,
    -- layer=1 filter=198 channel=25
    9, -4, -7, 12, 5, -4, -16, -5, 3,
    -- layer=1 filter=198 channel=26
    -2, 2, 0, -15, 4, -3, 0, -6, -21,
    -- layer=1 filter=198 channel=27
    0, -10, -7, 7, 2, 7, 2, 4, -9,
    -- layer=1 filter=198 channel=28
    -11, 13, -9, -2, 2, 0, -6, -2, 3,
    -- layer=1 filter=198 channel=29
    -1, 9, -8, 2, -1, -9, 4, -8, 4,
    -- layer=1 filter=198 channel=30
    -10, -13, -4, -8, -3, 0, 5, -3, -15,
    -- layer=1 filter=198 channel=31
    -5, -10, 2, -12, -6, 11, -7, 1, 4,
    -- layer=1 filter=198 channel=32
    0, -11, -2, -5, 0, -6, 0, -13, -17,
    -- layer=1 filter=198 channel=33
    -7, 6, -5, 0, 5, 0, -7, 9, 3,
    -- layer=1 filter=198 channel=34
    4, -9, -9, 3, -9, -11, -3, 1, -10,
    -- layer=1 filter=198 channel=35
    2, -5, 4, -3, 2, -4, -7, 0, -10,
    -- layer=1 filter=198 channel=36
    -8, -5, -3, -3, 3, -10, -8, -4, -10,
    -- layer=1 filter=198 channel=37
    9, 2, -8, 1, -7, 3, -1, -4, 0,
    -- layer=1 filter=198 channel=38
    0, 0, -6, -10, -16, -1, -14, 0, -3,
    -- layer=1 filter=198 channel=39
    -8, 4, 8, -6, -3, -5, -1, 7, -7,
    -- layer=1 filter=198 channel=40
    -10, 1, 1, -4, -1, -12, -1, -2, 2,
    -- layer=1 filter=198 channel=41
    2, -3, 7, 1, 0, -12, -4, 10, -11,
    -- layer=1 filter=198 channel=42
    12, 6, -10, 5, -13, -2, 2, -12, -15,
    -- layer=1 filter=198 channel=43
    11, 5, -1, 13, -9, -10, -7, 8, -11,
    -- layer=1 filter=198 channel=44
    -2, 4, -1, -8, 6, -9, 1, -4, -7,
    -- layer=1 filter=198 channel=45
    -7, 0, 5, 2, -7, -10, -2, -11, -15,
    -- layer=1 filter=198 channel=46
    6, 1, -8, -14, 6, -7, 16, 8, -1,
    -- layer=1 filter=198 channel=47
    -10, -6, 0, 1, -8, 0, -10, -8, -6,
    -- layer=1 filter=198 channel=48
    -5, -6, 5, 7, 2, -5, -9, -13, -15,
    -- layer=1 filter=198 channel=49
    4, -4, -5, -12, 0, -13, -12, 3, -8,
    -- layer=1 filter=198 channel=50
    -4, 5, -10, 0, 9, -8, 6, 4, -2,
    -- layer=1 filter=198 channel=51
    0, 0, -3, -3, -2, 2, -6, -2, -2,
    -- layer=1 filter=198 channel=52
    -6, 7, 3, -7, 8, 6, -5, 2, -10,
    -- layer=1 filter=198 channel=53
    -10, 8, -10, 7, -7, -8, 2, 7, 5,
    -- layer=1 filter=198 channel=54
    0, -4, -7, 4, 6, -1, 4, -5, 5,
    -- layer=1 filter=198 channel=55
    -13, -18, 0, -6, -2, -12, -10, -11, 5,
    -- layer=1 filter=198 channel=56
    -1, 3, -10, -7, 4, 2, -10, -1, -1,
    -- layer=1 filter=198 channel=57
    -4, -5, 2, 2, -2, -4, -3, -10, 1,
    -- layer=1 filter=198 channel=58
    -1, 1, -3, 10, -8, -1, -13, -11, -4,
    -- layer=1 filter=198 channel=59
    -11, -3, -8, -10, 1, -8, 0, -2, -4,
    -- layer=1 filter=198 channel=60
    6, 9, -8, 0, -4, -3, 3, 8, 4,
    -- layer=1 filter=198 channel=61
    -2, 2, 3, 0, -9, 8, -1, 6, 9,
    -- layer=1 filter=198 channel=62
    12, 2, -17, -17, -5, -5, 7, -5, -4,
    -- layer=1 filter=198 channel=63
    -13, -17, -15, -7, 1, -6, -13, -3, -7,
    -- layer=1 filter=198 channel=64
    -13, 7, -3, -4, -4, -1, -7, -7, 0,
    -- layer=1 filter=198 channel=65
    -10, 8, -6, -3, 3, -13, 2, 1, -5,
    -- layer=1 filter=198 channel=66
    -17, -16, -2, 4, -13, 0, -11, 4, -5,
    -- layer=1 filter=198 channel=67
    2, 2, -6, 2, -3, 8, -6, 0, -7,
    -- layer=1 filter=198 channel=68
    -6, -14, -10, 0, 6, 3, -16, 1, -5,
    -- layer=1 filter=198 channel=69
    -1, 2, -4, -6, 0, -17, -12, 1, -13,
    -- layer=1 filter=198 channel=70
    -1, -10, -10, 12, -3, -7, 0, -14, -8,
    -- layer=1 filter=198 channel=71
    -9, 9, -15, -5, -10, -5, -2, -3, -10,
    -- layer=1 filter=198 channel=72
    0, -9, 0, -7, -2, 9, 8, 0, 4,
    -- layer=1 filter=198 channel=73
    -10, 5, 3, 9, 1, 3, 3, -4, -10,
    -- layer=1 filter=198 channel=74
    -1, -11, -2, -5, 11, 0, 0, 7, -4,
    -- layer=1 filter=198 channel=75
    8, -3, -7, 2, 1, -3, -1, -2, -7,
    -- layer=1 filter=198 channel=76
    -8, -6, 1, -5, 4, 4, -11, -3, -9,
    -- layer=1 filter=198 channel=77
    -2, 0, -12, -6, 7, -10, 5, 0, 2,
    -- layer=1 filter=198 channel=78
    -1, 4, 2, -5, 2, -8, -1, 8, -8,
    -- layer=1 filter=198 channel=79
    4, -10, -7, 4, 3, 0, 0, -11, -15,
    -- layer=1 filter=198 channel=80
    8, -11, 2, 6, 5, -7, 2, -4, -2,
    -- layer=1 filter=198 channel=81
    6, -9, -6, 0, -4, 4, -6, -7, -9,
    -- layer=1 filter=198 channel=82
    -4, -6, 0, -1, -11, -4, -12, -17, 2,
    -- layer=1 filter=198 channel=83
    2, -4, -1, -3, 2, 0, -6, 0, 5,
    -- layer=1 filter=198 channel=84
    -6, -4, -7, -18, -5, 5, -6, 3, -5,
    -- layer=1 filter=198 channel=85
    6, -6, 2, 0, -6, -13, -3, 6, -7,
    -- layer=1 filter=198 channel=86
    1, -7, -21, -9, -7, -6, -12, -14, -3,
    -- layer=1 filter=198 channel=87
    1, -1, 1, 3, -7, 0, 9, 12, -9,
    -- layer=1 filter=198 channel=88
    12, 8, 3, 4, -5, 4, 0, -9, -9,
    -- layer=1 filter=198 channel=89
    -14, 2, -4, -6, 6, -9, -14, -17, 0,
    -- layer=1 filter=198 channel=90
    1, -13, -15, 3, 9, -4, -13, -7, -8,
    -- layer=1 filter=198 channel=91
    -13, -5, -11, 2, -5, 1, 1, -14, 0,
    -- layer=1 filter=198 channel=92
    -13, -5, 2, 0, -6, -7, 5, -11, 2,
    -- layer=1 filter=198 channel=93
    -1, -1, -10, -14, -8, -10, -5, -13, -6,
    -- layer=1 filter=198 channel=94
    0, 1, 4, -14, 2, 2, -9, -10, -8,
    -- layer=1 filter=198 channel=95
    0, -13, -1, -11, 7, -2, -13, 7, -11,
    -- layer=1 filter=198 channel=96
    0, 0, 8, -8, -3, 9, -7, 0, -6,
    -- layer=1 filter=198 channel=97
    -17, 1, -5, -9, -13, 0, -16, -12, -14,
    -- layer=1 filter=198 channel=98
    -3, 4, -1, -2, 3, 1, -16, -13, -1,
    -- layer=1 filter=198 channel=99
    -8, -9, 9, -20, 9, -3, -3, -16, 0,
    -- layer=1 filter=198 channel=100
    -6, 2, -10, -2, 2, 1, 5, 9, 5,
    -- layer=1 filter=198 channel=101
    -4, -12, -15, -15, -1, -6, -11, -5, -10,
    -- layer=1 filter=198 channel=102
    3, 1, -9, -12, 0, -7, -13, -4, -5,
    -- layer=1 filter=198 channel=103
    4, -4, -6, -9, -5, 13, -8, -10, 3,
    -- layer=1 filter=198 channel=104
    -7, 6, 0, -11, -4, -7, 5, 7, -3,
    -- layer=1 filter=198 channel=105
    -14, -10, -12, -3, -8, -1, -16, 0, 0,
    -- layer=1 filter=198 channel=106
    -9, -12, -12, -19, -12, 0, -3, -12, -20,
    -- layer=1 filter=198 channel=107
    8, 0, 5, -6, -11, -9, 0, 0, 0,
    -- layer=1 filter=198 channel=108
    -4, -2, 4, 4, -9, -4, -7, 4, -1,
    -- layer=1 filter=198 channel=109
    0, -9, 10, -1, 9, 3, 10, 5, -10,
    -- layer=1 filter=198 channel=110
    3, -5, -6, 1, -9, 1, -3, 5, 4,
    -- layer=1 filter=198 channel=111
    -4, -13, -3, -5, -12, 2, -2, -1, -11,
    -- layer=1 filter=198 channel=112
    6, -10, -16, -9, 9, 0, -7, -10, -11,
    -- layer=1 filter=198 channel=113
    18, -2, -1, 3, 5, -16, 3, -13, 0,
    -- layer=1 filter=198 channel=114
    0, -4, -13, 4, 5, -10, 7, -9, 3,
    -- layer=1 filter=198 channel=115
    -14, 0, -10, 4, -11, -12, -13, -13, -5,
    -- layer=1 filter=198 channel=116
    7, 9, 5, -7, -10, 2, -4, 8, -3,
    -- layer=1 filter=198 channel=117
    -3, -8, -14, -6, 6, 1, -5, -10, -5,
    -- layer=1 filter=198 channel=118
    -17, -17, 4, -10, 2, -1, -2, 8, 1,
    -- layer=1 filter=198 channel=119
    3, -11, 4, -6, -10, -12, -11, -13, -5,
    -- layer=1 filter=198 channel=120
    -4, 0, -5, -4, 5, -13, 0, -20, 4,
    -- layer=1 filter=198 channel=121
    -15, -9, -6, -6, -7, -3, -6, 1, 5,
    -- layer=1 filter=198 channel=122
    -1, 8, 3, 10, 9, 6, -6, -7, 4,
    -- layer=1 filter=198 channel=123
    -9, 4, 0, -6, -2, -14, 0, -3, -6,
    -- layer=1 filter=198 channel=124
    6, -7, -3, 6, 0, -3, -6, -7, -8,
    -- layer=1 filter=198 channel=125
    12, 6, 6, 12, -3, 4, -15, -4, 1,
    -- layer=1 filter=198 channel=126
    -10, -8, 1, 6, -10, 1, 5, 6, -4,
    -- layer=1 filter=198 channel=127
    -16, -15, 2, -18, 0, -10, -12, -5, -5,
    -- layer=1 filter=199 channel=0
    -8, -12, -15, -9, -8, 2, -32, -16, 4,
    -- layer=1 filter=199 channel=1
    -22, 4, -20, 1, -35, -16, -1, -7, -7,
    -- layer=1 filter=199 channel=2
    15, 10, -16, 7, -2, 3, 1, 2, -9,
    -- layer=1 filter=199 channel=3
    1, -5, 7, 7, 6, -10, 0, -9, -5,
    -- layer=1 filter=199 channel=4
    -10, -4, 0, -5, 3, 3, 10, -6, 4,
    -- layer=1 filter=199 channel=5
    -28, 12, -14, 22, -2, -7, 10, 17, 0,
    -- layer=1 filter=199 channel=6
    -5, 16, 23, 8, 8, -4, 76, 34, -14,
    -- layer=1 filter=199 channel=7
    -18, -5, 26, 12, -26, -21, 0, -11, 27,
    -- layer=1 filter=199 channel=8
    -39, -1, -19, -3, -26, -26, 8, 9, 28,
    -- layer=1 filter=199 channel=9
    -21, -20, -4, -37, -9, -41, 2, -5, -11,
    -- layer=1 filter=199 channel=10
    -10, 7, 23, 13, -37, -6, -16, -15, 35,
    -- layer=1 filter=199 channel=11
    17, 25, 28, 3, 35, 36, -8, 13, 20,
    -- layer=1 filter=199 channel=12
    5, 42, 22, -9, -6, -20, 12, 60, -31,
    -- layer=1 filter=199 channel=13
    -12, -26, -7, 1, -8, 0, 7, 29, -6,
    -- layer=1 filter=199 channel=14
    -48, 8, 44, 24, -34, -17, 0, 42, 21,
    -- layer=1 filter=199 channel=15
    -41, -25, -19, -18, -10, -15, -38, -24, -19,
    -- layer=1 filter=199 channel=16
    -27, -11, -41, 30, 18, -19, 30, 22, 23,
    -- layer=1 filter=199 channel=17
    -6, 2, -6, -4, -2, -5, -14, -7, 2,
    -- layer=1 filter=199 channel=18
    -21, -15, 15, 33, 30, 9, 0, 40, 8,
    -- layer=1 filter=199 channel=19
    20, -55, -33, -12, 3, 13, -15, 19, 0,
    -- layer=1 filter=199 channel=20
    -7, -20, -8, 4, -31, -21, 19, 16, 24,
    -- layer=1 filter=199 channel=21
    -37, -30, -24, -1, -24, -25, 17, -47, -7,
    -- layer=1 filter=199 channel=22
    -9, 11, -1, 40, 7, 1, 34, 24, 33,
    -- layer=1 filter=199 channel=23
    4, -38, 31, -25, 13, 9, 7, 23, 25,
    -- layer=1 filter=199 channel=24
    -6, -30, -47, -16, -39, -19, -22, -8, 11,
    -- layer=1 filter=199 channel=25
    -13, 0, -1, 12, -24, -12, -14, 2, 46,
    -- layer=1 filter=199 channel=26
    -25, -15, -8, -4, -4, -8, -1, 17, 34,
    -- layer=1 filter=199 channel=27
    -13, 13, -9, 7, 24, 17, -19, -3, -3,
    -- layer=1 filter=199 channel=28
    -36, -7, 3, 48, -29, -8, 7, 1, 26,
    -- layer=1 filter=199 channel=29
    -33, -14, -7, -30, -10, -9, -53, -30, -12,
    -- layer=1 filter=199 channel=30
    -17, -73, -32, -26, -41, -49, -37, -12, -31,
    -- layer=1 filter=199 channel=31
    17, 21, 37, 22, 11, 15, 26, 45, -22,
    -- layer=1 filter=199 channel=32
    -34, -50, -24, -48, -48, -30, -21, -50, -16,
    -- layer=1 filter=199 channel=33
    -13, 0, 0, -14, -6, -18, 5, -12, -8,
    -- layer=1 filter=199 channel=34
    -8, -2, -5, -5, -12, -19, -8, 4, -24,
    -- layer=1 filter=199 channel=35
    2, 0, -6, -12, -6, -12, -6, -8, -2,
    -- layer=1 filter=199 channel=36
    6, 30, 28, 23, 43, 46, 12, 32, 38,
    -- layer=1 filter=199 channel=37
    2, 20, -23, 27, 6, -2, 12, 26, 4,
    -- layer=1 filter=199 channel=38
    -14, -34, -26, -7, -34, -18, 36, 5, -6,
    -- layer=1 filter=199 channel=39
    8, 21, 8, -17, 12, 17, 2, 17, 23,
    -- layer=1 filter=199 channel=40
    1, 24, -10, 54, -4, -50, 87, 95, 16,
    -- layer=1 filter=199 channel=41
    -19, -17, -9, -54, 9, -18, -38, -31, 17,
    -- layer=1 filter=199 channel=42
    19, -6, -4, 0, -13, -11, 21, 7, -21,
    -- layer=1 filter=199 channel=43
    -11, 8, -16, 29, -13, -19, 6, 26, 27,
    -- layer=1 filter=199 channel=44
    -66, -46, -30, -45, -64, -21, -21, -42, 0,
    -- layer=1 filter=199 channel=45
    -57, -42, -28, -2, -32, -17, -16, -9, 0,
    -- layer=1 filter=199 channel=46
    -4, -26, 16, -27, -5, 37, 15, 37, -14,
    -- layer=1 filter=199 channel=47
    19, -19, 9, -36, 16, 3, 9, 4, 10,
    -- layer=1 filter=199 channel=48
    -1, -41, -32, -9, -34, -27, -5, -5, -1,
    -- layer=1 filter=199 channel=49
    -16, 3, 10, -23, -24, -29, -19, -13, -2,
    -- layer=1 filter=199 channel=50
    0, -8, -1, -1, 0, -12, -17, -3, -15,
    -- layer=1 filter=199 channel=51
    -20, -6, -9, 0, -43, -55, 14, -8, 16,
    -- layer=1 filter=199 channel=52
    5, -8, -28, 2, -5, -2, 19, 17, -11,
    -- layer=1 filter=199 channel=53
    0, -5, -1, -7, -3, -2, 5, 0, -6,
    -- layer=1 filter=199 channel=54
    19, -10, -21, 16, 11, 0, -5, 19, 43,
    -- layer=1 filter=199 channel=55
    26, 37, 23, 28, 53, 54, -2, 30, 26,
    -- layer=1 filter=199 channel=56
    2, -9, -4, -10, 1, 1, -6, 2, -2,
    -- layer=1 filter=199 channel=57
    -13, 8, 22, 33, -11, -7, 11, 6, 32,
    -- layer=1 filter=199 channel=58
    7, -33, 13, -18, -5, -1, -22, 35, 40,
    -- layer=1 filter=199 channel=59
    -11, -13, -6, 12, 12, -10, -13, -5, 1,
    -- layer=1 filter=199 channel=60
    15, 0, -3, 13, -8, 14, 16, 11, 15,
    -- layer=1 filter=199 channel=61
    3, -10, 8, -2, -1, 2, 11, 0, -2,
    -- layer=1 filter=199 channel=62
    -37, -34, -45, -3, -18, -17, -5, 14, 28,
    -- layer=1 filter=199 channel=63
    -3, 17, 12, 6, 37, 35, 4, 0, 5,
    -- layer=1 filter=199 channel=64
    3, -7, -1, 4, 0, 0, 1, -17, -8,
    -- layer=1 filter=199 channel=65
    -24, -37, -20, -7, -15, -21, 7, -16, -8,
    -- layer=1 filter=199 channel=66
    -11, 10, 2, -3, 7, 11, -28, -1, -10,
    -- layer=1 filter=199 channel=67
    3, 18, 27, 4, -22, 34, 77, 9, 42,
    -- layer=1 filter=199 channel=68
    -51, -36, -33, -44, -85, -24, -27, -36, -10,
    -- layer=1 filter=199 channel=69
    -40, 0, -42, 14, 2, -25, -5, 28, 23,
    -- layer=1 filter=199 channel=70
    47, 94, 73, -18, -2, -14, 63, 29, 10,
    -- layer=1 filter=199 channel=71
    -17, -1, 3, 8, -9, 13, -21, 4, 0,
    -- layer=1 filter=199 channel=72
    7, -59, -28, -7, -9, 0, 4, 19, 0,
    -- layer=1 filter=199 channel=73
    0, 15, 11, 14, -3, -4, 15, 13, 5,
    -- layer=1 filter=199 channel=74
    -23, -22, -26, -33, -25, -22, 3, 14, -17,
    -- layer=1 filter=199 channel=75
    -48, -46, 3, -15, -69, -57, 20, 42, -19,
    -- layer=1 filter=199 channel=76
    -20, -29, -3, -13, -9, -23, -9, -28, -3,
    -- layer=1 filter=199 channel=77
    -3, -24, -16, 17, -32, -11, 17, -26, -1,
    -- layer=1 filter=199 channel=78
    16, 14, 15, 7, 17, 1, 2, 21, 25,
    -- layer=1 filter=199 channel=79
    -17, -13, -37, 17, -10, -30, 8, 18, 31,
    -- layer=1 filter=199 channel=80
    9, -7, -10, -10, 4, 8, 3, -6, -6,
    -- layer=1 filter=199 channel=81
    3, -18, -43, 1, -15, -26, -6, 0, 7,
    -- layer=1 filter=199 channel=82
    -31, -56, -27, -7, -39, -20, 17, -24, -16,
    -- layer=1 filter=199 channel=83
    -26, -15, -28, -13, -34, -42, -16, -17, -16,
    -- layer=1 filter=199 channel=84
    -40, -50, -55, -21, -22, -46, -2, 14, 14,
    -- layer=1 filter=199 channel=85
    -6, -17, 3, -33, 13, 6, -38, 27, -17,
    -- layer=1 filter=199 channel=86
    4, 37, 28, 6, 41, 23, 3, 24, 21,
    -- layer=1 filter=199 channel=87
    28, -12, -8, -6, 16, -17, -13, 26, -15,
    -- layer=1 filter=199 channel=88
    14, 2, 17, 9, -10, -1, 3, 11, 23,
    -- layer=1 filter=199 channel=89
    -51, -34, -24, -26, -47, -30, 14, -29, -27,
    -- layer=1 filter=199 channel=90
    -54, -56, -54, -32, -61, -49, -26, -43, -4,
    -- layer=1 filter=199 channel=91
    9, -25, -24, 5, -35, -41, 41, 0, -4,
    -- layer=1 filter=199 channel=92
    -53, -4, -44, -43, 7, 2, -14, -8, -11,
    -- layer=1 filter=199 channel=93
    -26, -36, -34, -24, -47, -25, -18, -26, -2,
    -- layer=1 filter=199 channel=94
    -18, 0, 0, -9, -4, -2, -28, -15, 1,
    -- layer=1 filter=199 channel=95
    -73, -52, -38, -16, -45, -46, -24, 2, -29,
    -- layer=1 filter=199 channel=96
    24, 11, 12, 21, 17, 5, 9, 4, 1,
    -- layer=1 filter=199 channel=97
    -19, 3, 0, 1, -4, -3, -9, -9, 15,
    -- layer=1 filter=199 channel=98
    -21, -37, -35, 14, -33, -21, 6, -3, 11,
    -- layer=1 filter=199 channel=99
    -54, -30, -4, 4, -52, -20, 2, -21, 32,
    -- layer=1 filter=199 channel=100
    -9, 23, 28, -3, 42, 43, -29, -4, -8,
    -- layer=1 filter=199 channel=101
    -27, -28, -19, -31, -39, -40, 29, -20, -17,
    -- layer=1 filter=199 channel=102
    -28, -20, -6, -5, -10, -23, -21, -22, -24,
    -- layer=1 filter=199 channel=103
    0, 15, 22, -13, 34, 29, -10, 6, -3,
    -- layer=1 filter=199 channel=104
    -9, -29, 10, -36, -8, 22, -4, 7, 45,
    -- layer=1 filter=199 channel=105
    -14, 9, 3, -11, 2, 13, -3, -14, 12,
    -- layer=1 filter=199 channel=106
    -17, -21, -16, -37, -64, -32, 18, -21, -47,
    -- layer=1 filter=199 channel=107
    -8, 0, 2, 9, 6, -2, -15, 2, 3,
    -- layer=1 filter=199 channel=108
    -49, -69, -44, -43, -61, -45, -40, -29, 9,
    -- layer=1 filter=199 channel=109
    7, -7, -8, -10, -9, 6, 5, 6, 4,
    -- layer=1 filter=199 channel=110
    6, 7, -8, 0, 3, 5, -7, -8, 7,
    -- layer=1 filter=199 channel=111
    -40, -56, -23, -15, -28, -57, -13, 18, 1,
    -- layer=1 filter=199 channel=112
    -21, -7, 5, -13, -16, -23, 0, -4, -1,
    -- layer=1 filter=199 channel=113
    -4, 1, 9, 2, 6, 3, 24, 14, 0,
    -- layer=1 filter=199 channel=114
    -3, 17, -5, 20, 34, 18, 34, 39, 26,
    -- layer=1 filter=199 channel=115
    -10, 30, 30, 13, 33, 22, -12, 13, 37,
    -- layer=1 filter=199 channel=116
    -6, 5, 4, -7, -8, 8, 1, 8, -4,
    -- layer=1 filter=199 channel=117
    -44, -30, 60, -7, -22, -90, 18, 48, 36,
    -- layer=1 filter=199 channel=118
    -39, -55, -38, -37, -29, -65, 5, 1, -34,
    -- layer=1 filter=199 channel=119
    -26, -40, -41, -56, -63, -50, -53, -62, -29,
    -- layer=1 filter=199 channel=120
    -13, -26, -20, 5, -23, -57, 6, -9, 6,
    -- layer=1 filter=199 channel=121
    -2, 6, 20, 1, 25, 27, -14, 10, -10,
    -- layer=1 filter=199 channel=122
    10, -7, -2, -10, 0, 4, -4, -2, -5,
    -- layer=1 filter=199 channel=123
    -11, 4, 22, 6, 44, 41, -19, 7, 16,
    -- layer=1 filter=199 channel=124
    10, -10, 3, 13, 12, 4, -3, 9, -1,
    -- layer=1 filter=199 channel=125
    13, 62, 62, 10, -11, -25, 45, 44, 14,
    -- layer=1 filter=199 channel=126
    -8, -19, -20, -5, -68, -70, -2, -46, -21,
    -- layer=1 filter=199 channel=127
    -41, -54, -5, -32, -24, -39, -4, -5, -32,
    -- layer=1 filter=200 channel=0
    6, -1, 0, 1, -3, 3, -3, -7, -11,
    -- layer=1 filter=200 channel=1
    -2, -5, -8, -7, 1, 5, 1, 1, -9,
    -- layer=1 filter=200 channel=2
    0, -8, -3, 2, -7, -5, 0, -4, 5,
    -- layer=1 filter=200 channel=3
    -9, 3, 0, 7, -4, 5, 0, 3, 6,
    -- layer=1 filter=200 channel=4
    -2, -5, -4, 0, 0, -3, 3, -7, -9,
    -- layer=1 filter=200 channel=5
    3, -1, -7, -7, -4, 5, 0, -9, -9,
    -- layer=1 filter=200 channel=6
    -6, -7, -1, -2, -7, 0, 6, -9, 0,
    -- layer=1 filter=200 channel=7
    4, 2, -3, 1, -10, 3, -3, -3, -10,
    -- layer=1 filter=200 channel=8
    4, 0, -4, -2, 3, -9, -7, -13, 2,
    -- layer=1 filter=200 channel=9
    -2, -4, -5, -14, 0, 1, -11, 4, 0,
    -- layer=1 filter=200 channel=10
    -4, -5, -3, -2, 0, 2, 5, 0, 6,
    -- layer=1 filter=200 channel=11
    2, 0, -1, 0, -5, -1, -13, 2, -5,
    -- layer=1 filter=200 channel=12
    10, -10, 7, 3, -4, 4, -14, -1, 6,
    -- layer=1 filter=200 channel=13
    -4, -15, -13, -3, -3, -6, -10, -1, -16,
    -- layer=1 filter=200 channel=14
    12, 3, -1, -3, -10, -12, -10, -14, -3,
    -- layer=1 filter=200 channel=15
    0, -3, 2, -12, 7, -9, -5, -5, 4,
    -- layer=1 filter=200 channel=16
    -6, -12, -7, 5, 0, -3, 0, -7, -15,
    -- layer=1 filter=200 channel=17
    -3, -11, 0, -5, 3, -12, 3, 4, 1,
    -- layer=1 filter=200 channel=18
    -7, -1, -3, 9, 4, 4, 5, 5, 2,
    -- layer=1 filter=200 channel=19
    0, 1, -3, -5, 0, 8, 7, -9, -2,
    -- layer=1 filter=200 channel=20
    -2, -6, -11, -10, -14, 7, -12, 5, -13,
    -- layer=1 filter=200 channel=21
    -8, 13, -3, -8, -12, -2, -11, 0, 4,
    -- layer=1 filter=200 channel=22
    6, 0, -4, -9, -11, -9, -5, 3, 4,
    -- layer=1 filter=200 channel=23
    5, -6, -9, -10, -10, 7, -12, -6, -8,
    -- layer=1 filter=200 channel=24
    6, -10, 6, -3, 3, 7, 0, -2, -20,
    -- layer=1 filter=200 channel=25
    5, -1, -8, 1, 0, 0, -11, -6, 4,
    -- layer=1 filter=200 channel=26
    -3, 0, -4, -9, -4, -7, -9, 0, 0,
    -- layer=1 filter=200 channel=27
    3, 11, -10, -10, -12, -14, -8, -5, 3,
    -- layer=1 filter=200 channel=28
    0, -14, -6, 7, 6, -8, -3, -10, -5,
    -- layer=1 filter=200 channel=29
    -4, 3, -2, 10, -7, 5, -11, -5, -2,
    -- layer=1 filter=200 channel=30
    -1, -6, 12, -9, 1, -4, 0, -1, -10,
    -- layer=1 filter=200 channel=31
    0, -5, -6, -7, -9, -5, -1, -5, -1,
    -- layer=1 filter=200 channel=32
    -2, 3, 3, -8, 3, -12, 0, -8, 0,
    -- layer=1 filter=200 channel=33
    3, -9, -4, 10, -10, 8, 3, -4, 3,
    -- layer=1 filter=200 channel=34
    6, 3, -1, 1, 3, 3, -2, 0, -2,
    -- layer=1 filter=200 channel=35
    1, 2, -11, -8, -1, -9, -10, 4, 0,
    -- layer=1 filter=200 channel=36
    4, 4, 0, 3, -2, -9, -3, -7, 5,
    -- layer=1 filter=200 channel=37
    -3, -8, -8, 8, -10, -7, -14, -14, -16,
    -- layer=1 filter=200 channel=38
    5, -1, 1, -10, -7, -2, -15, -5, -11,
    -- layer=1 filter=200 channel=39
    6, -1, -7, -9, 7, -9, 1, -9, -8,
    -- layer=1 filter=200 channel=40
    9, -4, -7, 4, 4, -19, 10, -1, -2,
    -- layer=1 filter=200 channel=41
    -4, -12, -14, -3, -5, -10, 5, 1, 6,
    -- layer=1 filter=200 channel=42
    -4, 8, -6, 1, 6, -6, 14, -8, 3,
    -- layer=1 filter=200 channel=43
    -1, -1, 0, 2, -7, -3, 1, -7, 0,
    -- layer=1 filter=200 channel=44
    5, 5, 0, -10, -3, -4, -10, -6, 4,
    -- layer=1 filter=200 channel=45
    0, -6, 0, -15, 5, 0, -12, -8, -14,
    -- layer=1 filter=200 channel=46
    -7, -3, -7, 8, -12, -11, -8, 5, -13,
    -- layer=1 filter=200 channel=47
    3, 15, -2, -18, 4, -7, 5, 10, -1,
    -- layer=1 filter=200 channel=48
    -12, 0, -7, -9, 3, -8, 1, -7, -1,
    -- layer=1 filter=200 channel=49
    -13, -3, -1, -12, 8, -10, -3, 4, -17,
    -- layer=1 filter=200 channel=50
    -11, -7, 3, -6, -10, 2, 2, -11, -4,
    -- layer=1 filter=200 channel=51
    -6, -10, -7, 3, -5, -2, 2, -3, -12,
    -- layer=1 filter=200 channel=52
    -2, -7, 8, 10, 7, 1, 2, 6, -1,
    -- layer=1 filter=200 channel=53
    5, -9, 0, 0, -10, -11, -3, -8, -3,
    -- layer=1 filter=200 channel=54
    -2, -10, -9, -1, 10, -3, -12, 2, -5,
    -- layer=1 filter=200 channel=55
    6, 0, -1, 8, -2, -3, 3, -16, -13,
    -- layer=1 filter=200 channel=56
    7, -5, -11, -10, 5, -1, 0, -2, 2,
    -- layer=1 filter=200 channel=57
    1, 1, 0, -10, -1, -6, -5, -12, 4,
    -- layer=1 filter=200 channel=58
    1, -7, -2, 5, 2, -6, -1, -4, -3,
    -- layer=1 filter=200 channel=59
    1, 0, -4, 0, -1, 2, -1, 0, 2,
    -- layer=1 filter=200 channel=60
    0, 0, -10, -6, 9, 11, 7, -5, 0,
    -- layer=1 filter=200 channel=61
    0, -8, -5, -9, 3, -1, 2, -6, -3,
    -- layer=1 filter=200 channel=62
    6, -11, 4, 5, 5, -5, 1, -13, -6,
    -- layer=1 filter=200 channel=63
    -15, -4, 0, -4, 3, 2, 3, -3, 4,
    -- layer=1 filter=200 channel=64
    -4, -12, -3, -10, -12, -5, -2, 0, -9,
    -- layer=1 filter=200 channel=65
    -11, -11, -4, -10, -10, 7, 4, -1, 0,
    -- layer=1 filter=200 channel=66
    -1, -2, -1, -6, 0, -9, -5, -10, 3,
    -- layer=1 filter=200 channel=67
    4, 11, 0, -5, -5, -2, 4, -7, 3,
    -- layer=1 filter=200 channel=68
    -13, -4, 6, -8, 13, -15, -9, 0, -16,
    -- layer=1 filter=200 channel=69
    8, -13, 8, 3, -2, 4, 3, -7, -7,
    -- layer=1 filter=200 channel=70
    -11, -3, 10, -13, 0, -8, 4, -7, -8,
    -- layer=1 filter=200 channel=71
    -4, -8, -9, -2, -6, -1, -6, -4, 1,
    -- layer=1 filter=200 channel=72
    7, 3, -5, -15, 4, -5, 7, 0, 6,
    -- layer=1 filter=200 channel=73
    0, 4, 2, -1, -1, -6, 6, -1, -7,
    -- layer=1 filter=200 channel=74
    -4, 6, -4, -10, -5, 5, 8, -7, -5,
    -- layer=1 filter=200 channel=75
    -7, -2, 0, -2, -12, -17, 3, 5, 2,
    -- layer=1 filter=200 channel=76
    -1, -5, -11, 1, -3, 4, -5, 5, 7,
    -- layer=1 filter=200 channel=77
    -11, -3, -10, -2, -8, -1, 1, 5, 0,
    -- layer=1 filter=200 channel=78
    2, -2, 6, -1, -7, 0, 6, 5, -6,
    -- layer=1 filter=200 channel=79
    9, -15, 0, 0, 6, 8, -13, -5, -1,
    -- layer=1 filter=200 channel=80
    9, 10, 6, 9, -9, 7, 1, 6, 0,
    -- layer=1 filter=200 channel=81
    2, -2, 4, -3, 4, 9, 1, -1, -5,
    -- layer=1 filter=200 channel=82
    2, -3, -3, -4, 4, -2, 1, 1, -8,
    -- layer=1 filter=200 channel=83
    3, -1, -10, 5, 0, -2, 1, -3, 0,
    -- layer=1 filter=200 channel=84
    0, 4, -9, -13, 6, 3, 10, -9, -8,
    -- layer=1 filter=200 channel=85
    0, 3, -4, 2, 6, 7, -5, 2, -4,
    -- layer=1 filter=200 channel=86
    -6, -6, 3, 0, -15, -10, -1, -6, 1,
    -- layer=1 filter=200 channel=87
    -3, -11, 0, 2, -6, 5, -9, -7, 2,
    -- layer=1 filter=200 channel=88
    -9, -17, -3, -2, 5, 5, -12, -11, -1,
    -- layer=1 filter=200 channel=89
    -17, 3, -10, 1, -3, -15, 1, -3, -3,
    -- layer=1 filter=200 channel=90
    0, -8, -12, 3, 1, -4, -7, -13, 0,
    -- layer=1 filter=200 channel=91
    -3, -9, -15, -13, -7, -5, -7, 1, -1,
    -- layer=1 filter=200 channel=92
    3, -6, 0, -12, -10, 7, 0, -2, 1,
    -- layer=1 filter=200 channel=93
    1, 3, 5, 2, -2, 8, -4, 2, -8,
    -- layer=1 filter=200 channel=94
    2, -1, 4, 0, -3, 6, 6, -7, -4,
    -- layer=1 filter=200 channel=95
    -12, -12, -4, 0, 5, -1, 10, -5, 3,
    -- layer=1 filter=200 channel=96
    2, -12, -4, -10, 7, -6, -11, -12, -5,
    -- layer=1 filter=200 channel=97
    -4, 5, -11, 7, -5, -12, 5, 0, 0,
    -- layer=1 filter=200 channel=98
    7, -13, -12, -5, 4, 3, 0, -15, -12,
    -- layer=1 filter=200 channel=99
    -7, -9, 2, 8, -10, -6, -7, 3, -11,
    -- layer=1 filter=200 channel=100
    0, -5, -5, -4, 5, 4, -8, -1, -10,
    -- layer=1 filter=200 channel=101
    -3, -3, -6, -9, 2, -9, 5, -4, -9,
    -- layer=1 filter=200 channel=102
    -5, 4, -7, -4, -13, 6, 0, 4, -8,
    -- layer=1 filter=200 channel=103
    5, -10, -7, -9, 7, -1, -13, -1, 2,
    -- layer=1 filter=200 channel=104
    6, -11, -9, -4, -9, -12, 7, -3, 8,
    -- layer=1 filter=200 channel=105
    -10, -15, -11, -1, -13, 0, -11, -3, 0,
    -- layer=1 filter=200 channel=106
    -3, 4, -11, -13, 0, 0, 0, 0, -3,
    -- layer=1 filter=200 channel=107
    4, -7, -7, 0, -1, 0, 4, -2, 1,
    -- layer=1 filter=200 channel=108
    0, 2, 11, -1, 5, -8, 7, -4, -15,
    -- layer=1 filter=200 channel=109
    1, 6, 7, 8, 1, -1, 6, 5, 1,
    -- layer=1 filter=200 channel=110
    -8, -13, -1, 7, -7, -3, 4, -5, 2,
    -- layer=1 filter=200 channel=111
    10, -11, 7, -10, 0, 5, -7, -6, 0,
    -- layer=1 filter=200 channel=112
    -6, -4, 5, 2, 4, 4, 5, 0, -1,
    -- layer=1 filter=200 channel=113
    0, 7, 10, -6, -10, -11, -4, -13, -5,
    -- layer=1 filter=200 channel=114
    3, -1, -1, 5, 2, -14, -13, -13, -12,
    -- layer=1 filter=200 channel=115
    -3, -5, -10, 0, -3, -10, 0, -4, -5,
    -- layer=1 filter=200 channel=116
    -1, -1, 1, 1, 8, -1, 9, 10, 8,
    -- layer=1 filter=200 channel=117
    4, 2, 3, -7, 7, 6, 0, -5, 2,
    -- layer=1 filter=200 channel=118
    -4, 1, 2, 5, -4, 0, 2, -7, -4,
    -- layer=1 filter=200 channel=119
    -9, -2, 8, -12, 12, -10, 3, -12, -6,
    -- layer=1 filter=200 channel=120
    -11, -2, -15, -1, 4, -4, -3, -3, 2,
    -- layer=1 filter=200 channel=121
    11, -2, -2, -5, -13, -11, 4, -7, 8,
    -- layer=1 filter=200 channel=122
    1, 6, 5, -4, -6, -1, 4, 2, 6,
    -- layer=1 filter=200 channel=123
    -6, 2, 5, 0, -8, -7, 8, -6, -13,
    -- layer=1 filter=200 channel=124
    8, 1, -4, 0, 0, 0, 3, 1, 4,
    -- layer=1 filter=200 channel=125
    0, -6, -6, 9, 2, -6, -1, 0, -7,
    -- layer=1 filter=200 channel=126
    -3, 8, 0, 0, 4, 5, -8, -11, -7,
    -- layer=1 filter=200 channel=127
    -4, 5, 6, -5, 4, -3, 9, -10, 6,
    -- layer=1 filter=201 channel=0
    7, 5, 4, 2, 4, -2, 8, -7, -2,
    -- layer=1 filter=201 channel=1
    -5, -7, -2, 4, -2, -12, -3, 7, 6,
    -- layer=1 filter=201 channel=2
    0, 0, 8, -10, -6, -2, -2, 5, 2,
    -- layer=1 filter=201 channel=3
    3, -6, -8, 3, -4, 11, 7, 5, 4,
    -- layer=1 filter=201 channel=4
    5, 0, -5, 6, 2, 5, -12, -5, -2,
    -- layer=1 filter=201 channel=5
    1, 0, 3, -2, -7, 5, -8, -8, 0,
    -- layer=1 filter=201 channel=6
    -8, 1, -9, -8, 4, -11, -10, 0, -6,
    -- layer=1 filter=201 channel=7
    1, -6, -2, -8, 5, -1, -10, 4, -1,
    -- layer=1 filter=201 channel=8
    6, 0, 5, 6, 7, -9, -4, -7, 3,
    -- layer=1 filter=201 channel=9
    4, -8, 7, -3, -7, 4, -11, -2, -10,
    -- layer=1 filter=201 channel=10
    5, 1, -7, -6, -4, -3, 8, 7, 0,
    -- layer=1 filter=201 channel=11
    -1, -1, -7, -1, -10, -13, -1, 0, -8,
    -- layer=1 filter=201 channel=12
    9, -4, 0, 8, 6, 0, -2, -1, 7,
    -- layer=1 filter=201 channel=13
    2, 7, 5, -11, 8, -2, -2, 8, -5,
    -- layer=1 filter=201 channel=14
    10, 8, 5, -5, -10, 7, 4, 5, 2,
    -- layer=1 filter=201 channel=15
    1, 0, 0, -9, 5, 2, 5, -5, -12,
    -- layer=1 filter=201 channel=16
    -8, -2, -3, -2, 8, -4, 3, 7, 0,
    -- layer=1 filter=201 channel=17
    -7, -3, -1, -5, -8, -1, 0, -2, -10,
    -- layer=1 filter=201 channel=18
    -3, -11, 0, -10, -9, -8, -10, -2, 6,
    -- layer=1 filter=201 channel=19
    -2, -4, 5, -9, 0, -12, -2, 5, 0,
    -- layer=1 filter=201 channel=20
    6, -9, 5, -11, -8, -10, -7, -6, 5,
    -- layer=1 filter=201 channel=21
    0, 5, 6, 5, -1, -5, 2, 4, 5,
    -- layer=1 filter=201 channel=22
    2, 8, -2, 3, 10, -4, -4, -10, 1,
    -- layer=1 filter=201 channel=23
    -8, -12, -2, -8, -8, 0, 2, -12, -7,
    -- layer=1 filter=201 channel=24
    0, 7, -2, -1, 8, 7, 7, 6, 1,
    -- layer=1 filter=201 channel=25
    -7, 2, 10, 6, -1, -5, 2, -6, -6,
    -- layer=1 filter=201 channel=26
    -9, -2, -4, 0, -1, 8, -3, 12, 2,
    -- layer=1 filter=201 channel=27
    0, -5, -1, 9, -11, -7, 0, 0, 1,
    -- layer=1 filter=201 channel=28
    0, 1, -3, 8, 0, -6, 5, 0, -11,
    -- layer=1 filter=201 channel=29
    -2, 7, 0, -11, -1, 5, 0, -2, -12,
    -- layer=1 filter=201 channel=30
    -10, -11, 2, 0, -8, 1, -5, -3, -5,
    -- layer=1 filter=201 channel=31
    5, -1, -8, -4, -10, 8, -6, -9, 0,
    -- layer=1 filter=201 channel=32
    8, 9, 1, -7, -12, 4, -7, -1, -1,
    -- layer=1 filter=201 channel=33
    -1, -9, -6, -8, 3, 0, -8, 2, 0,
    -- layer=1 filter=201 channel=34
    -7, 0, 6, 7, 4, 8, 0, 0, -5,
    -- layer=1 filter=201 channel=35
    -12, 3, -12, 5, 0, 2, 5, 8, 5,
    -- layer=1 filter=201 channel=36
    2, -8, -12, -10, -10, -12, -10, 1, 0,
    -- layer=1 filter=201 channel=37
    9, -1, 0, -8, -6, -1, -4, -2, 5,
    -- layer=1 filter=201 channel=38
    3, 0, 0, -5, 3, 3, -5, 0, 7,
    -- layer=1 filter=201 channel=39
    -2, 4, 1, 4, 6, 6, 1, 0, 3,
    -- layer=1 filter=201 channel=40
    2, 2, 10, 3, -7, -4, -6, 9, -11,
    -- layer=1 filter=201 channel=41
    -4, 7, -2, 2, 4, 2, -12, -5, 4,
    -- layer=1 filter=201 channel=42
    -1, -5, -8, 4, 0, -6, 4, -6, 5,
    -- layer=1 filter=201 channel=43
    7, 3, -5, -10, -8, 3, -6, -2, -4,
    -- layer=1 filter=201 channel=44
    -12, -7, 7, -3, -1, -13, -7, -3, -13,
    -- layer=1 filter=201 channel=45
    3, -11, -9, -9, -9, 4, -8, -5, -7,
    -- layer=1 filter=201 channel=46
    -8, 5, 6, 0, 1, 3, 5, 5, -1,
    -- layer=1 filter=201 channel=47
    8, -7, -1, 3, 3, 1, 9, 1, -8,
    -- layer=1 filter=201 channel=48
    -10, 3, -8, 5, -6, -10, 0, -5, -5,
    -- layer=1 filter=201 channel=49
    8, -13, -12, 5, 2, 4, 0, 6, 7,
    -- layer=1 filter=201 channel=50
    -4, 0, -7, -9, 0, 7, -3, 6, 0,
    -- layer=1 filter=201 channel=51
    8, 0, -3, -6, 1, 3, -9, -8, 4,
    -- layer=1 filter=201 channel=52
    3, -10, 3, 7, 0, -8, -5, -6, -7,
    -- layer=1 filter=201 channel=53
    1, -2, -3, -9, -7, -3, -8, -12, 2,
    -- layer=1 filter=201 channel=54
    -4, -9, 7, -2, 3, -2, -4, -12, 3,
    -- layer=1 filter=201 channel=55
    2, 0, 2, 1, -4, -3, -9, -2, -11,
    -- layer=1 filter=201 channel=56
    -3, 7, 2, 0, 0, 8, -5, -10, 4,
    -- layer=1 filter=201 channel=57
    6, -7, -10, -1, 6, -2, -6, 2, 7,
    -- layer=1 filter=201 channel=58
    1, -8, 2, 6, -9, 7, 4, -7, -7,
    -- layer=1 filter=201 channel=59
    7, -9, -1, -10, 0, 3, 5, -8, -2,
    -- layer=1 filter=201 channel=60
    3, -6, 5, 6, 9, 3, -8, 1, 4,
    -- layer=1 filter=201 channel=61
    3, -5, -10, 3, 9, -7, 1, 1, -3,
    -- layer=1 filter=201 channel=62
    7, 6, 3, -9, 3, -7, -9, 6, -9,
    -- layer=1 filter=201 channel=63
    1, -8, -3, 6, -5, 0, 6, 0, -5,
    -- layer=1 filter=201 channel=64
    -1, -10, -12, 7, -5, -3, -4, -2, -6,
    -- layer=1 filter=201 channel=65
    -8, -1, -1, -5, 0, -7, -6, 4, -7,
    -- layer=1 filter=201 channel=66
    -8, -11, 2, -10, -7, -5, 7, -8, -5,
    -- layer=1 filter=201 channel=67
    0, -8, -5, 4, -4, 6, -2, -3, 7,
    -- layer=1 filter=201 channel=68
    6, 3, -2, 0, -7, 4, -3, -3, -12,
    -- layer=1 filter=201 channel=69
    5, -5, -9, 1, -5, -1, -6, 2, 4,
    -- layer=1 filter=201 channel=70
    -5, -3, -1, 8, 3, 11, -4, -5, -9,
    -- layer=1 filter=201 channel=71
    -8, -7, -4, -8, 3, -1, -11, -1, 2,
    -- layer=1 filter=201 channel=72
    0, -2, 5, -7, 4, -10, 3, -2, -3,
    -- layer=1 filter=201 channel=73
    -1, 0, -12, -7, 1, 5, -3, 3, 4,
    -- layer=1 filter=201 channel=74
    -2, 6, 5, -1, 0, -1, 5, -10, 4,
    -- layer=1 filter=201 channel=75
    -5, 8, 7, 6, 6, 1, 0, 9, -9,
    -- layer=1 filter=201 channel=76
    -11, -1, 0, 7, -3, -12, 4, 7, -6,
    -- layer=1 filter=201 channel=77
    2, 7, -8, -10, -11, 0, -12, -8, -6,
    -- layer=1 filter=201 channel=78
    1, -11, 5, 0, 4, -3, -9, 3, 0,
    -- layer=1 filter=201 channel=79
    -2, -10, 2, -4, 1, 6, -3, 3, 4,
    -- layer=1 filter=201 channel=80
    1, 6, -7, 2, 1, -5, 9, 0, -1,
    -- layer=1 filter=201 channel=81
    2, 0, 3, -9, -11, 1, 3, 6, -12,
    -- layer=1 filter=201 channel=82
    0, 0, 1, -12, -7, -7, -11, -8, -5,
    -- layer=1 filter=201 channel=83
    -2, 8, 7, 0, 7, -6, 7, -8, 5,
    -- layer=1 filter=201 channel=84
    4, 0, -1, -10, 4, -3, 1, 10, 7,
    -- layer=1 filter=201 channel=85
    -9, -7, -4, 8, 8, -7, 4, -1, -2,
    -- layer=1 filter=201 channel=86
    0, 1, -4, 1, -10, -7, 3, -3, 5,
    -- layer=1 filter=201 channel=87
    -6, -2, -12, -4, -5, 7, 1, 2, -11,
    -- layer=1 filter=201 channel=88
    1, -9, 6, 5, 6, 2, 5, -1, -1,
    -- layer=1 filter=201 channel=89
    -1, 8, -4, 6, -9, -6, 2, -10, -2,
    -- layer=1 filter=201 channel=90
    4, 0, 1, 4, 0, -9, 5, 2, -6,
    -- layer=1 filter=201 channel=91
    1, 5, 6, -8, 0, -8, 5, 7, -10,
    -- layer=1 filter=201 channel=92
    -2, -8, -12, -5, 0, -4, -5, -7, 4,
    -- layer=1 filter=201 channel=93
    -1, 8, -7, -6, -6, 8, 2, 4, -3,
    -- layer=1 filter=201 channel=94
    5, -7, 6, 6, 7, -9, 0, 0, 4,
    -- layer=1 filter=201 channel=95
    -2, 8, -11, 0, 0, 6, -4, -1, 5,
    -- layer=1 filter=201 channel=96
    -8, -3, 0, 3, -11, 4, 5, 1, 3,
    -- layer=1 filter=201 channel=97
    -3, -8, -2, 3, -4, 7, 4, 4, 2,
    -- layer=1 filter=201 channel=98
    -9, -2, 10, 6, -4, -6, 4, -8, -10,
    -- layer=1 filter=201 channel=99
    6, -5, -9, 4, -10, 5, -4, -4, -11,
    -- layer=1 filter=201 channel=100
    -12, -11, 0, 5, 5, -12, 0, 6, -6,
    -- layer=1 filter=201 channel=101
    -5, 7, 0, -11, -10, -3, 3, -11, 0,
    -- layer=1 filter=201 channel=102
    -8, -4, 1, 3, -2, 8, 4, 1, -1,
    -- layer=1 filter=201 channel=103
    4, -8, -3, 4, -5, 0, -7, -5, -2,
    -- layer=1 filter=201 channel=104
    0, -9, -10, -3, 0, 6, -2, -9, -7,
    -- layer=1 filter=201 channel=105
    -5, 2, 5, 0, -5, 7, 4, 7, -12,
    -- layer=1 filter=201 channel=106
    0, 6, 6, 4, -6, -6, 9, -2, -10,
    -- layer=1 filter=201 channel=107
    -4, 7, 3, 5, -4, 2, -7, 5, -3,
    -- layer=1 filter=201 channel=108
    -11, -5, 7, 0, -1, -7, -2, 8, 7,
    -- layer=1 filter=201 channel=109
    4, 6, -5, 9, -4, 8, 0, -5, -6,
    -- layer=1 filter=201 channel=110
    -4, -4, -11, 1, -9, -7, -8, 0, -1,
    -- layer=1 filter=201 channel=111
    -8, 0, 1, -6, -7, -5, -8, 3, 0,
    -- layer=1 filter=201 channel=112
    -4, -10, -6, 5, -2, 0, 5, 1, 5,
    -- layer=1 filter=201 channel=113
    4, -5, -6, 3, 3, 1, 5, -2, 4,
    -- layer=1 filter=201 channel=114
    -4, 5, 5, -10, 0, -4, -8, 1, -6,
    -- layer=1 filter=201 channel=115
    -9, 0, 1, -11, -2, -6, 3, 4, 4,
    -- layer=1 filter=201 channel=116
    -2, -6, -2, 3, 5, -6, 8, 9, -1,
    -- layer=1 filter=201 channel=117
    4, 8, -7, -11, 0, 0, 9, 11, 4,
    -- layer=1 filter=201 channel=118
    -11, -2, 6, -3, -5, 1, -3, -2, -1,
    -- layer=1 filter=201 channel=119
    -11, 1, -2, -5, 5, -10, 8, 6, 10,
    -- layer=1 filter=201 channel=120
    -8, 4, -2, -11, -7, -5, 5, 6, 1,
    -- layer=1 filter=201 channel=121
    0, -2, -3, 6, 7, 3, -10, 4, -6,
    -- layer=1 filter=201 channel=122
    4, 8, 1, -4, -4, 2, -9, 8, 8,
    -- layer=1 filter=201 channel=123
    -12, -12, -4, -12, -4, -12, 1, -9, -10,
    -- layer=1 filter=201 channel=124
    -10, 3, -4, -4, -7, 3, 7, -6, -9,
    -- layer=1 filter=201 channel=125
    -6, 4, 1, 0, 9, -7, -1, 5, 4,
    -- layer=1 filter=201 channel=126
    -9, -8, -5, -6, 8, -6, -3, 6, -9,
    -- layer=1 filter=201 channel=127
    -8, 0, 2, 1, 4, 6, 6, 0, 1,
    -- layer=1 filter=202 channel=0
    -1, -17, 3, 3, 0, -8, -10, 2, -13,
    -- layer=1 filter=202 channel=1
    0, -7, -8, 4, 5, 7, -10, -12, -2,
    -- layer=1 filter=202 channel=2
    3, -12, 7, 2, -2, -11, -5, -10, -13,
    -- layer=1 filter=202 channel=3
    1, 2, -2, 4, -9, -7, -7, -7, 1,
    -- layer=1 filter=202 channel=4
    0, -10, -12, 6, 5, 0, -8, 2, -9,
    -- layer=1 filter=202 channel=5
    -8, 0, 1, 17, 16, 1, -8, -8, -25,
    -- layer=1 filter=202 channel=6
    -2, -4, -9, 15, -7, 9, 12, 8, 2,
    -- layer=1 filter=202 channel=7
    -20, 0, -11, -2, -9, 0, -5, 2, -23,
    -- layer=1 filter=202 channel=8
    0, -2, 1, 2, -4, 5, -19, -12, 1,
    -- layer=1 filter=202 channel=9
    0, -18, -10, -10, 3, 0, -2, 9, -5,
    -- layer=1 filter=202 channel=10
    -12, -4, -18, 5, -3, -20, -11, -10, -23,
    -- layer=1 filter=202 channel=11
    -7, -6, -17, -21, -13, -4, -6, -7, 0,
    -- layer=1 filter=202 channel=12
    -16, -2, -2, -3, 2, -5, -13, 0, -20,
    -- layer=1 filter=202 channel=13
    -5, -5, -14, -5, -3, -1, -3, -3, 6,
    -- layer=1 filter=202 channel=14
    -5, -4, -4, -4, -6, -17, 6, 2, -17,
    -- layer=1 filter=202 channel=15
    5, 7, -3, 3, 0, -7, 1, -2, 1,
    -- layer=1 filter=202 channel=16
    5, 4, -2, 9, 12, 6, -14, -20, -24,
    -- layer=1 filter=202 channel=17
    -17, -13, -16, -2, 1, -3, -10, -3, 0,
    -- layer=1 filter=202 channel=18
    -6, 1, -4, -3, -20, -17, -6, 0, -14,
    -- layer=1 filter=202 channel=19
    -7, 0, -11, -11, -1, 1, 1, 2, -12,
    -- layer=1 filter=202 channel=20
    -17, -1, -4, -7, -8, 6, -2, 7, -2,
    -- layer=1 filter=202 channel=21
    0, -4, -19, -4, -15, -14, -14, -21, -12,
    -- layer=1 filter=202 channel=22
    4, -1, -19, 5, 10, 0, 8, 0, -10,
    -- layer=1 filter=202 channel=23
    -19, 6, -9, -7, -9, -8, -12, -6, 2,
    -- layer=1 filter=202 channel=24
    -9, -1, -9, -17, -6, -24, -13, -21, -7,
    -- layer=1 filter=202 channel=25
    -10, -10, -13, -5, 0, 1, -20, -4, -6,
    -- layer=1 filter=202 channel=26
    -3, -19, -13, -2, -23, 8, 3, -10, 5,
    -- layer=1 filter=202 channel=27
    2, 6, 7, 1, 5, -1, 4, -13, -5,
    -- layer=1 filter=202 channel=28
    -8, -21, 0, 0, 0, -16, -8, -11, -6,
    -- layer=1 filter=202 channel=29
    -10, -10, -13, -12, -7, 1, -19, -17, -10,
    -- layer=1 filter=202 channel=30
    -7, 0, -15, -4, -25, -31, -19, -19, -8,
    -- layer=1 filter=202 channel=31
    -8, -10, -2, 5, -17, -9, 3, 2, -3,
    -- layer=1 filter=202 channel=32
    -12, -16, -14, -7, -11, -10, -5, -3, 0,
    -- layer=1 filter=202 channel=33
    -11, -12, -1, 2, -4, -5, -3, -6, 1,
    -- layer=1 filter=202 channel=34
    -1, 7, 1, -4, 4, -4, 0, 3, 7,
    -- layer=1 filter=202 channel=35
    -8, -2, -4, -6, -2, 5, 5, -2, -4,
    -- layer=1 filter=202 channel=36
    -1, -16, -15, -14, 1, 2, -12, -2, -14,
    -- layer=1 filter=202 channel=37
    8, -7, -3, -3, -2, -6, -28, -7, -31,
    -- layer=1 filter=202 channel=38
    -7, -8, -22, 2, -1, -14, -3, -2, 1,
    -- layer=1 filter=202 channel=39
    2, -10, -12, -6, -4, -4, -13, -8, -3,
    -- layer=1 filter=202 channel=40
    2, 0, 2, -11, 4, 5, 0, 14, -1,
    -- layer=1 filter=202 channel=41
    7, -11, 6, -12, -11, -7, 6, 0, 3,
    -- layer=1 filter=202 channel=42
    0, -8, 3, -2, 0, 4, -3, -18, -15,
    -- layer=1 filter=202 channel=43
    -1, 0, -14, 0, 0, 0, -19, -9, -12,
    -- layer=1 filter=202 channel=44
    -1, -7, 2, 0, -3, -15, -9, -14, -3,
    -- layer=1 filter=202 channel=45
    -13, -14, -11, -7, -7, -12, -12, -23, -6,
    -- layer=1 filter=202 channel=46
    7, 2, 2, 0, -10, 3, 10, 4, -12,
    -- layer=1 filter=202 channel=47
    -11, -14, 0, -10, -13, -5, -5, -4, 9,
    -- layer=1 filter=202 channel=48
    -5, -1, -2, -16, -14, -17, -13, -8, -8,
    -- layer=1 filter=202 channel=49
    -15, -12, -21, -12, 0, -19, -5, -14, -3,
    -- layer=1 filter=202 channel=50
    -11, 4, -7, -6, -4, 3, -4, -10, -7,
    -- layer=1 filter=202 channel=51
    -10, -19, 0, -17, -9, -18, -3, -14, -17,
    -- layer=1 filter=202 channel=52
    -5, 4, 9, -7, -3, 4, -4, 7, 10,
    -- layer=1 filter=202 channel=53
    -5, 4, 6, 7, 3, -3, 1, -9, -3,
    -- layer=1 filter=202 channel=54
    4, -3, -17, 0, -3, -13, -2, -16, -19,
    -- layer=1 filter=202 channel=55
    -7, -4, -6, 2, 6, 8, 5, 7, 9,
    -- layer=1 filter=202 channel=56
    -7, 6, 6, 3, 6, -10, 5, 4, -11,
    -- layer=1 filter=202 channel=57
    -4, -9, 0, -1, -15, -1, -9, -5, -10,
    -- layer=1 filter=202 channel=58
    -4, -6, -7, 2, -14, -4, 3, 2, 0,
    -- layer=1 filter=202 channel=59
    2, 0, 7, 1, -1, 7, -10, -10, -3,
    -- layer=1 filter=202 channel=60
    -10, -8, 3, 6, 2, 4, -5, 1, -8,
    -- layer=1 filter=202 channel=61
    6, 3, -5, 0, 4, -7, 3, 0, -8,
    -- layer=1 filter=202 channel=62
    -3, -7, 0, 15, 0, -4, -24, -29, -17,
    -- layer=1 filter=202 channel=63
    -1, -8, -8, -21, -19, -6, -10, 0, -4,
    -- layer=1 filter=202 channel=64
    -10, -17, -4, -11, -12, -2, -3, 0, -10,
    -- layer=1 filter=202 channel=65
    -5, -12, -3, -3, -5, 0, -1, -14, -12,
    -- layer=1 filter=202 channel=66
    1, -2, -5, 0, 3, -13, 5, 1, -4,
    -- layer=1 filter=202 channel=67
    12, 7, -11, 18, 12, 1, -7, 3, 11,
    -- layer=1 filter=202 channel=68
    -4, -17, 0, -17, -11, -21, -16, -7, -6,
    -- layer=1 filter=202 channel=69
    -12, 1, -2, -2, 11, 13, -17, -21, -10,
    -- layer=1 filter=202 channel=70
    1, -8, 3, 4, 4, -5, 23, 15, 10,
    -- layer=1 filter=202 channel=71
    -15, -2, -12, -15, -16, -19, -14, -11, -11,
    -- layer=1 filter=202 channel=72
    -15, 0, -1, -3, -12, -5, -2, -3, -5,
    -- layer=1 filter=202 channel=73
    5, 8, 4, -2, -6, -1, 0, -7, 3,
    -- layer=1 filter=202 channel=74
    -11, 4, -9, -9, -4, -12, -5, 7, 2,
    -- layer=1 filter=202 channel=75
    -10, -7, -4, -12, -22, -19, 0, -18, -27,
    -- layer=1 filter=202 channel=76
    -14, -7, -5, -8, -4, 0, -14, -3, -16,
    -- layer=1 filter=202 channel=77
    -10, -17, 0, -18, -15, -18, -9, 0, -15,
    -- layer=1 filter=202 channel=78
    -5, 0, 4, -6, 2, -10, -3, -2, -9,
    -- layer=1 filter=202 channel=79
    -4, 0, 1, 10, 9, 3, -23, -8, -10,
    -- layer=1 filter=202 channel=80
    2, -3, -4, 0, -4, -2, -8, -9, -4,
    -- layer=1 filter=202 channel=81
    0, -12, -6, -8, -14, -14, -4, -2, -18,
    -- layer=1 filter=202 channel=82
    -21, -8, -8, -19, -12, -8, -18, -10, -1,
    -- layer=1 filter=202 channel=83
    -3, -17, -8, -4, 3, -15, -13, -9, -15,
    -- layer=1 filter=202 channel=84
    -4, 0, 0, -12, -22, -2, -9, -11, 10,
    -- layer=1 filter=202 channel=85
    -2, 2, -1, -6, 0, 1, -2, -1, 0,
    -- layer=1 filter=202 channel=86
    -1, 2, 2, 2, 0, 0, -4, 0, -14,
    -- layer=1 filter=202 channel=87
    -8, 7, -9, 2, -2, -2, 3, -5, 3,
    -- layer=1 filter=202 channel=88
    -7, -16, -27, -7, -18, -10, -6, -5, -10,
    -- layer=1 filter=202 channel=89
    -3, -24, -26, -23, -20, -19, -22, -16, -17,
    -- layer=1 filter=202 channel=90
    -12, -10, -16, -11, -18, 1, 3, -18, 1,
    -- layer=1 filter=202 channel=91
    -11, -12, -8, 0, -15, -3, -11, 8, 5,
    -- layer=1 filter=202 channel=92
    -13, 4, -9, 7, 3, 0, -8, -9, 9,
    -- layer=1 filter=202 channel=93
    -11, -9, -17, -8, 1, 1, -7, -12, 0,
    -- layer=1 filter=202 channel=94
    -17, -13, -8, -1, -2, -6, 5, -4, -7,
    -- layer=1 filter=202 channel=95
    0, -13, -15, -11, -11, -17, -4, -20, -15,
    -- layer=1 filter=202 channel=96
    -4, -6, -7, -11, 3, -4, -8, -2, 0,
    -- layer=1 filter=202 channel=97
    -18, -15, -1, 3, 0, -11, -6, -5, -6,
    -- layer=1 filter=202 channel=98
    2, -8, -8, 12, 8, 5, -28, -10, -19,
    -- layer=1 filter=202 channel=99
    -5, -5, -11, -14, -18, -1, -10, -11, -7,
    -- layer=1 filter=202 channel=100
    -9, -3, -13, 1, -12, 3, -11, 1, -4,
    -- layer=1 filter=202 channel=101
    -6, -8, -20, 2, -4, -10, -7, -9, -4,
    -- layer=1 filter=202 channel=102
    2, -14, -9, -1, -15, -12, 4, -4, -14,
    -- layer=1 filter=202 channel=103
    0, -16, -11, -23, -10, -21, -10, 4, -5,
    -- layer=1 filter=202 channel=104
    -7, -1, -12, -12, -10, -9, -17, -12, -11,
    -- layer=1 filter=202 channel=105
    -7, -5, -9, -16, -7, -10, 0, -9, -10,
    -- layer=1 filter=202 channel=106
    -16, -22, -20, -7, -16, -11, 3, 3, -1,
    -- layer=1 filter=202 channel=107
    6, -5, 7, -4, 8, -10, 0, 6, -8,
    -- layer=1 filter=202 channel=108
    -10, -2, -16, -8, -21, 0, -5, -23, -10,
    -- layer=1 filter=202 channel=109
    2, -1, 8, -6, 6, 2, 9, 9, -6,
    -- layer=1 filter=202 channel=110
    -16, -7, -14, 0, -1, -10, -1, 2, -1,
    -- layer=1 filter=202 channel=111
    2, -6, -16, -15, -13, -15, -16, -9, -9,
    -- layer=1 filter=202 channel=112
    -3, -4, 3, -9, -2, 6, -2, -5, 3,
    -- layer=1 filter=202 channel=113
    -2, 1, -6, 2, -3, 4, 12, 4, 0,
    -- layer=1 filter=202 channel=114
    7, 3, 7, 5, 13, -2, -14, -5, -24,
    -- layer=1 filter=202 channel=115
    -9, -4, -16, -2, -11, -12, 4, -11, 4,
    -- layer=1 filter=202 channel=116
    -9, 3, -9, 5, 5, 4, -2, 10, -7,
    -- layer=1 filter=202 channel=117
    -4, -3, 5, -7, -11, -14, 8, 1, -11,
    -- layer=1 filter=202 channel=118
    4, -3, -8, -16, -23, -23, -20, -5, -9,
    -- layer=1 filter=202 channel=119
    -4, -15, -4, -5, -29, -17, -16, -13, -6,
    -- layer=1 filter=202 channel=120
    -3, -7, -15, 2, 3, -8, -4, -17, -8,
    -- layer=1 filter=202 channel=121
    -4, -8, -9, 0, -10, -13, -15, -14, -17,
    -- layer=1 filter=202 channel=122
    -4, -4, 9, 1, -6, 5, -5, 2, -8,
    -- layer=1 filter=202 channel=123
    -5, -16, -1, -2, -13, -12, -16, -11, -20,
    -- layer=1 filter=202 channel=124
    8, -1, -7, 2, 7, -1, -8, -9, -3,
    -- layer=1 filter=202 channel=125
    -1, 2, -2, 6, 0, 9, 8, 14, 7,
    -- layer=1 filter=202 channel=126
    -12, -3, -7, 8, 9, -4, -18, 0, -11,
    -- layer=1 filter=202 channel=127
    5, 0, -7, -19, -16, -14, -2, -4, 0,
    -- layer=1 filter=203 channel=0
    -12, 4, 5, -11, 0, 5, 7, 4, -10,
    -- layer=1 filter=203 channel=1
    -5, -7, -12, -7, -5, -1, -1, -11, 9,
    -- layer=1 filter=203 channel=2
    5, 0, 1, -8, 0, 1, 6, 10, -8,
    -- layer=1 filter=203 channel=3
    2, -5, 0, 9, 3, -8, -4, -8, 6,
    -- layer=1 filter=203 channel=4
    -10, 2, 5, 5, 8, 4, -9, -3, -9,
    -- layer=1 filter=203 channel=5
    -1, -8, 0, 3, -10, 0, -4, -7, 6,
    -- layer=1 filter=203 channel=6
    -3, -7, -6, -9, -10, -6, 0, 4, 0,
    -- layer=1 filter=203 channel=7
    -6, -9, -1, -9, -14, 4, 4, -1, -14,
    -- layer=1 filter=203 channel=8
    -1, 8, -7, 0, 7, 4, -4, -4, -4,
    -- layer=1 filter=203 channel=9
    7, -7, -7, -3, -1, 6, 3, -6, -3,
    -- layer=1 filter=203 channel=10
    -4, 5, -6, -2, 3, -9, -11, -1, -11,
    -- layer=1 filter=203 channel=11
    2, 7, -12, -2, 6, 3, 1, 0, -9,
    -- layer=1 filter=203 channel=12
    -1, -7, 0, 2, 5, 9, 9, 1, 6,
    -- layer=1 filter=203 channel=13
    2, -9, 4, -11, -1, 0, -10, 3, -10,
    -- layer=1 filter=203 channel=14
    -3, -2, 4, 4, -1, 0, 1, -1, -6,
    -- layer=1 filter=203 channel=15
    -8, 3, -7, -8, 2, 3, 7, -2, -3,
    -- layer=1 filter=203 channel=16
    -13, -8, -11, -5, -12, -11, -10, 9, -6,
    -- layer=1 filter=203 channel=17
    2, 8, -5, 3, 0, -1, -9, 1, -6,
    -- layer=1 filter=203 channel=18
    4, -4, -5, -8, -5, 7, -7, 1, -12,
    -- layer=1 filter=203 channel=19
    0, 0, 4, 0, 5, 0, 6, -11, 3,
    -- layer=1 filter=203 channel=20
    -5, -8, -3, 8, -6, -7, 0, 6, 5,
    -- layer=1 filter=203 channel=21
    -10, -1, 1, -7, -13, 7, -10, 0, -6,
    -- layer=1 filter=203 channel=22
    7, 6, 6, 2, 5, -2, -1, 9, -7,
    -- layer=1 filter=203 channel=23
    -7, -4, -11, -12, -10, 6, -10, -12, 8,
    -- layer=1 filter=203 channel=24
    -1, -8, -10, -3, -10, -11, -8, -2, -2,
    -- layer=1 filter=203 channel=25
    7, -11, 4, -13, -5, -12, -9, -5, -4,
    -- layer=1 filter=203 channel=26
    6, 0, -10, -12, -12, -6, 0, -12, -11,
    -- layer=1 filter=203 channel=27
    -6, 5, -3, 5, 3, -4, 5, 5, 8,
    -- layer=1 filter=203 channel=28
    -11, -4, 7, -3, -6, -6, 7, 3, 8,
    -- layer=1 filter=203 channel=29
    5, -8, -4, 5, 4, -12, -7, -5, 2,
    -- layer=1 filter=203 channel=30
    -1, -3, 9, 1, 3, -5, -4, -8, 5,
    -- layer=1 filter=203 channel=31
    6, -9, 7, -9, -4, -3, 7, 8, 3,
    -- layer=1 filter=203 channel=32
    -3, 1, 5, 7, -1, -10, -11, 1, -7,
    -- layer=1 filter=203 channel=33
    3, 2, -4, -10, -1, -8, 9, -8, 9,
    -- layer=1 filter=203 channel=34
    1, 4, 3, -5, 4, -9, 7, -4, 3,
    -- layer=1 filter=203 channel=35
    7, 5, -9, -5, -2, 3, -3, 8, 5,
    -- layer=1 filter=203 channel=36
    0, -4, 2, -9, 8, -4, -3, 4, 4,
    -- layer=1 filter=203 channel=37
    4, 3, 3, 5, 2, 5, -6, -1, -6,
    -- layer=1 filter=203 channel=38
    4, -3, 4, -7, -3, 1, -3, 7, -5,
    -- layer=1 filter=203 channel=39
    1, -1, -8, -5, 3, 1, -4, -2, -7,
    -- layer=1 filter=203 channel=40
    -6, -2, 0, -11, -12, -11, -12, 3, -7,
    -- layer=1 filter=203 channel=41
    3, 8, -3, -8, -1, -10, 7, -8, 5,
    -- layer=1 filter=203 channel=42
    -5, 8, -6, 7, 7, 10, -8, -8, 4,
    -- layer=1 filter=203 channel=43
    5, 3, -6, 0, -12, 4, -8, -11, -6,
    -- layer=1 filter=203 channel=44
    6, 0, -6, -3, 4, -7, -1, 0, -2,
    -- layer=1 filter=203 channel=45
    4, -5, 2, -6, 4, 4, -11, -12, -3,
    -- layer=1 filter=203 channel=46
    9, 2, -2, 0, -7, 9, 12, 10, 6,
    -- layer=1 filter=203 channel=47
    5, -4, 10, 5, -8, 7, 0, -3, 5,
    -- layer=1 filter=203 channel=48
    0, -8, -3, 4, 0, -7, 6, -7, -6,
    -- layer=1 filter=203 channel=49
    -7, 0, 3, -7, 7, -9, 0, -8, -9,
    -- layer=1 filter=203 channel=50
    -11, -9, -10, -1, -9, 4, -4, -7, -4,
    -- layer=1 filter=203 channel=51
    8, -1, -8, 6, -6, -1, 3, 0, -9,
    -- layer=1 filter=203 channel=52
    9, 2, 2, 8, 1, -7, -9, 4, -4,
    -- layer=1 filter=203 channel=53
    -5, 1, 5, 0, 0, -5, -5, 6, 8,
    -- layer=1 filter=203 channel=54
    7, 0, 1, -10, 1, -3, -1, 1, -11,
    -- layer=1 filter=203 channel=55
    -9, -10, 0, -3, -10, 0, 5, -11, 4,
    -- layer=1 filter=203 channel=56
    1, 7, -3, 3, 1, 5, 4, 6, 9,
    -- layer=1 filter=203 channel=57
    0, -8, 0, 8, 7, 6, 0, -5, -8,
    -- layer=1 filter=203 channel=58
    0, 0, 6, 0, -4, -11, -5, 1, 1,
    -- layer=1 filter=203 channel=59
    3, 3, -10, -9, -6, -6, 5, -10, -4,
    -- layer=1 filter=203 channel=60
    -6, -8, 5, 8, 9, -10, -11, 6, 5,
    -- layer=1 filter=203 channel=61
    -4, 0, -2, 5, -9, 6, -1, 0, -1,
    -- layer=1 filter=203 channel=62
    -4, 0, 5, -2, -3, -1, 6, 4, -4,
    -- layer=1 filter=203 channel=63
    6, -4, -4, 0, -1, 5, 6, -1, 6,
    -- layer=1 filter=203 channel=64
    -9, -1, 6, -4, -4, 0, 7, 2, 6,
    -- layer=1 filter=203 channel=65
    2, 7, 3, -9, -8, -5, -6, -5, 5,
    -- layer=1 filter=203 channel=66
    -11, 1, -9, 6, -4, -4, -2, -5, -11,
    -- layer=1 filter=203 channel=67
    1, -9, -3, -10, -8, -1, 8, -4, -10,
    -- layer=1 filter=203 channel=68
    -3, 0, -11, -1, -5, 4, 7, -10, -6,
    -- layer=1 filter=203 channel=69
    6, -10, 3, -6, 4, 0, 0, -9, 7,
    -- layer=1 filter=203 channel=70
    0, 0, 5, -12, 8, 2, 8, 2, 2,
    -- layer=1 filter=203 channel=71
    7, -7, -4, -1, 3, 2, -6, -11, -10,
    -- layer=1 filter=203 channel=72
    -10, 2, 2, 2, -6, -2, -12, 4, 4,
    -- layer=1 filter=203 channel=73
    6, 3, -12, 5, 8, -7, 0, 5, 3,
    -- layer=1 filter=203 channel=74
    2, 7, 0, 2, 0, 2, -3, 4, -1,
    -- layer=1 filter=203 channel=75
    3, -7, -7, 9, -8, 0, 2, 3, -6,
    -- layer=1 filter=203 channel=76
    -2, 1, -4, -9, -11, 6, -8, -9, 4,
    -- layer=1 filter=203 channel=77
    0, -4, -9, 7, -4, 3, -4, -1, -4,
    -- layer=1 filter=203 channel=78
    6, -7, 2, -1, 6, 0, 7, 2, -10,
    -- layer=1 filter=203 channel=79
    -5, 6, 3, 4, -6, 2, 2, 5, 3,
    -- layer=1 filter=203 channel=80
    -7, 0, -2, -8, -1, 2, 5, -5, -1,
    -- layer=1 filter=203 channel=81
    -2, 3, 3, -5, 6, 8, 2, 0, -7,
    -- layer=1 filter=203 channel=82
    -7, -2, 1, -8, -4, -2, 1, -2, -5,
    -- layer=1 filter=203 channel=83
    1, 5, -6, -6, 8, 7, -10, -7, 2,
    -- layer=1 filter=203 channel=84
    6, 0, -11, -3, -5, 1, -8, -9, -6,
    -- layer=1 filter=203 channel=85
    3, -4, -3, 0, -9, -2, -1, -3, -4,
    -- layer=1 filter=203 channel=86
    6, 2, 4, 1, -11, 0, -5, 1, -9,
    -- layer=1 filter=203 channel=87
    4, -9, 7, -11, 4, -3, 5, -11, 0,
    -- layer=1 filter=203 channel=88
    -6, 2, -4, 0, -3, 1, 8, -3, 0,
    -- layer=1 filter=203 channel=89
    -9, 2, 0, -11, -7, 7, -5, 7, 5,
    -- layer=1 filter=203 channel=90
    0, 3, 0, -11, -11, -5, -7, 1, 7,
    -- layer=1 filter=203 channel=91
    5, -8, -4, 5, 1, 8, -10, 4, 0,
    -- layer=1 filter=203 channel=92
    7, 3, -6, -9, 0, -4, 3, -6, -9,
    -- layer=1 filter=203 channel=93
    6, -8, -6, -1, 6, 0, -9, 0, 7,
    -- layer=1 filter=203 channel=94
    -7, -12, 7, 2, -2, 0, -7, -3, -4,
    -- layer=1 filter=203 channel=95
    2, -7, 1, 1, 7, 0, -8, -5, -3,
    -- layer=1 filter=203 channel=96
    -9, -2, -1, 0, -10, -8, 0, 8, -6,
    -- layer=1 filter=203 channel=97
    0, -5, 0, -4, 4, 1, -11, -10, 6,
    -- layer=1 filter=203 channel=98
    -8, -7, 0, 0, 4, -9, 4, 7, -5,
    -- layer=1 filter=203 channel=99
    7, 3, 2, 4, -3, -6, 3, -11, -2,
    -- layer=1 filter=203 channel=100
    3, 5, 5, -3, -10, -9, -6, -2, -3,
    -- layer=1 filter=203 channel=101
    -4, -7, -2, 0, 0, -4, -1, -10, 8,
    -- layer=1 filter=203 channel=102
    -4, -9, -9, -8, 5, -6, 6, -3, -10,
    -- layer=1 filter=203 channel=103
    -6, -10, 5, -1, -3, -3, 7, -10, 5,
    -- layer=1 filter=203 channel=104
    -5, -4, -3, 8, -10, 8, 2, 5, 1,
    -- layer=1 filter=203 channel=105
    -4, -8, 7, 0, -3, 2, -3, 4, 0,
    -- layer=1 filter=203 channel=106
    -4, -1, -6, 1, 2, 5, -10, 4, -4,
    -- layer=1 filter=203 channel=107
    -2, -2, -8, -4, 0, -10, -11, 10, -7,
    -- layer=1 filter=203 channel=108
    -5, -5, 5, 3, 0, 2, -11, -7, -3,
    -- layer=1 filter=203 channel=109
    -2, -6, -1, 4, 3, 8, -9, -2, -9,
    -- layer=1 filter=203 channel=110
    -4, -4, -2, -2, -8, 0, 0, 2, 7,
    -- layer=1 filter=203 channel=111
    4, 6, 8, -1, 5, -2, 2, -1, 1,
    -- layer=1 filter=203 channel=112
    -3, 8, 6, -1, 4, -11, -1, -8, -8,
    -- layer=1 filter=203 channel=113
    -5, -1, 7, -6, -6, -3, 2, -9, 8,
    -- layer=1 filter=203 channel=114
    -1, -7, 6, -6, -11, 2, -4, -5, -2,
    -- layer=1 filter=203 channel=115
    0, -7, 2, -4, 0, -6, 0, -4, 9,
    -- layer=1 filter=203 channel=116
    8, -7, -8, 0, 4, 2, 9, -10, -1,
    -- layer=1 filter=203 channel=117
    -5, -2, 0, -11, -10, -1, 5, -12, 1,
    -- layer=1 filter=203 channel=118
    -4, -5, 0, 4, -3, -7, 1, -4, -10,
    -- layer=1 filter=203 channel=119
    -4, -16, -9, 1, 2, -7, -2, 6, 6,
    -- layer=1 filter=203 channel=120
    -10, 7, -9, -11, 0, -6, -11, 2, 3,
    -- layer=1 filter=203 channel=121
    1, -11, -10, -6, -13, 6, -5, -4, 0,
    -- layer=1 filter=203 channel=122
    -3, -2, 8, 0, 10, 4, 3, -9, 3,
    -- layer=1 filter=203 channel=123
    -6, -11, 0, 3, -9, 6, -5, -11, 7,
    -- layer=1 filter=203 channel=124
    2, 4, 0, 5, -2, -2, -10, 0, 6,
    -- layer=1 filter=203 channel=125
    -7, 10, 6, -9, 5, 0, 7, -3, -7,
    -- layer=1 filter=203 channel=126
    -4, 2, -2, 8, -1, 8, -4, -6, 6,
    -- layer=1 filter=203 channel=127
    6, -1, -5, 1, 10, 0, -3, 0, 8,
    -- layer=1 filter=204 channel=0
    0, 6, 6, -6, -2, 14, -4, -8, 0,
    -- layer=1 filter=204 channel=1
    -14, -27, -21, 9, -10, -16, 10, 12, 10,
    -- layer=1 filter=204 channel=2
    -16, -3, 0, -3, 16, 7, 22, 45, 42,
    -- layer=1 filter=204 channel=3
    -8, -8, 4, -4, 7, -8, 5, -4, 13,
    -- layer=1 filter=204 channel=4
    -7, -17, -4, -2, 1, -2, 6, 0, -5,
    -- layer=1 filter=204 channel=5
    -7, -15, -6, -5, -13, -19, 20, 4, 0,
    -- layer=1 filter=204 channel=6
    -59, -60, -68, -8, -16, -17, 36, 15, 38,
    -- layer=1 filter=204 channel=7
    -39, -108, -66, -103, -217, -89, -80, -155, -95,
    -- layer=1 filter=204 channel=8
    13, -1, 12, 24, 2, 2, 15, 32, 36,
    -- layer=1 filter=204 channel=9
    -53, -43, -11, -17, -20, -8, 27, 19, 11,
    -- layer=1 filter=204 channel=10
    -53, -104, -60, -72, -186, -96, -45, -133, -94,
    -- layer=1 filter=204 channel=11
    1, 4, 12, -13, 7, -1, -31, -39, -23,
    -- layer=1 filter=204 channel=12
    -37, -31, -7, -47, -11, 5, -4, 19, 32,
    -- layer=1 filter=204 channel=13
    -15, -7, -32, 8, -2, -12, 26, 21, 13,
    -- layer=1 filter=204 channel=14
    13, -40, -16, -52, -26, -17, 0, -16, -40,
    -- layer=1 filter=204 channel=15
    -31, -25, 1, -3, -27, -12, 0, -17, 7,
    -- layer=1 filter=204 channel=16
    26, 5, 26, 23, 19, 5, 22, 22, 22,
    -- layer=1 filter=204 channel=17
    3, -10, -11, 8, -4, -12, -1, -1, -24,
    -- layer=1 filter=204 channel=18
    -7, 11, -1, 7, -4, 14, 0, 17, 21,
    -- layer=1 filter=204 channel=19
    32, 23, 39, 63, 69, 44, 49, 25, 36,
    -- layer=1 filter=204 channel=20
    -14, -4, -11, 5, 1, -13, 28, 12, 11,
    -- layer=1 filter=204 channel=21
    -26, -12, -20, 3, -2, 1, 7, 23, 18,
    -- layer=1 filter=204 channel=22
    -36, -27, -27, 19, 7, -2, 35, 20, 31,
    -- layer=1 filter=204 channel=23
    25, -69, -6, -44, -101, -38, -38, -80, -26,
    -- layer=1 filter=204 channel=24
    0, 18, 11, -4, 8, 12, 10, 20, 9,
    -- layer=1 filter=204 channel=25
    -13, -58, -4, -25, -73, -63, -8, -42, -11,
    -- layer=1 filter=204 channel=26
    14, 16, 11, 21, -15, -31, 0, -3, -14,
    -- layer=1 filter=204 channel=27
    -8, 4, 3, -16, 10, -5, -31, -17, 5,
    -- layer=1 filter=204 channel=28
    -18, -55, -41, -22, -95, -65, -18, -81, -67,
    -- layer=1 filter=204 channel=29
    -5, 0, -19, -2, 9, 2, -17, 3, -10,
    -- layer=1 filter=204 channel=30
    46, 26, 34, 15, 11, 32, 45, 37, 41,
    -- layer=1 filter=204 channel=31
    -41, -47, -24, -9, -3, 9, 28, 63, 48,
    -- layer=1 filter=204 channel=32
    9, -5, -16, -24, -53, -71, -22, -51, -23,
    -- layer=1 filter=204 channel=33
    -10, -5, -3, 5, 1, 19, 19, 2, -7,
    -- layer=1 filter=204 channel=34
    -26, -40, -21, -16, 0, -16, -2, 23, -18,
    -- layer=1 filter=204 channel=35
    0, -8, -8, -2, 8, -3, 4, 4, 6,
    -- layer=1 filter=204 channel=36
    6, 20, 8, -13, 4, -3, -26, -14, -25,
    -- layer=1 filter=204 channel=37
    30, 14, 25, 0, 8, -4, 26, 17, 7,
    -- layer=1 filter=204 channel=38
    -17, -17, -29, 10, -3, -8, 28, 28, 14,
    -- layer=1 filter=204 channel=39
    9, 5, 10, -14, -18, -9, -9, -3, 11,
    -- layer=1 filter=204 channel=40
    -22, -54, -41, 8, 6, 10, 62, 46, 43,
    -- layer=1 filter=204 channel=41
    -21, -43, 6, -24, -85, -46, -36, -49, -14,
    -- layer=1 filter=204 channel=42
    -9, 1, 36, -3, -1, 20, 34, 23, 36,
    -- layer=1 filter=204 channel=43
    0, 3, 7, 26, -11, -8, 8, 11, 17,
    -- layer=1 filter=204 channel=44
    -45, -42, -49, -13, -62, -71, -45, -55, -38,
    -- layer=1 filter=204 channel=45
    -33, -26, -16, 8, -16, -1, 0, -6, -3,
    -- layer=1 filter=204 channel=46
    36, 12, 42, 61, 55, 23, 111, 71, 69,
    -- layer=1 filter=204 channel=47
    9, -66, 3, -49, -59, -59, -10, 1, -7,
    -- layer=1 filter=204 channel=48
    2, -3, -2, 7, -3, 2, 23, 7, 10,
    -- layer=1 filter=204 channel=49
    0, -21, 0, 5, 1, -2, 8, 14, 32,
    -- layer=1 filter=204 channel=50
    -23, -51, -36, -8, 7, 2, -3, 10, -2,
    -- layer=1 filter=204 channel=51
    2, -5, -13, 6, -17, -6, 36, 6, 21,
    -- layer=1 filter=204 channel=52
    16, 12, 21, 21, 2, 33, 7, 8, 21,
    -- layer=1 filter=204 channel=53
    13, 4, 9, 6, 1, 16, 16, 14, 20,
    -- layer=1 filter=204 channel=54
    6, -17, 16, -17, -39, -49, -11, -41, -5,
    -- layer=1 filter=204 channel=55
    8, 18, 29, 3, 19, 14, -14, 3, 8,
    -- layer=1 filter=204 channel=56
    -8, -4, 0, 6, 0, -2, -7, 7, -6,
    -- layer=1 filter=204 channel=57
    -47, -111, -42, -45, -106, -49, 12, -42, -27,
    -- layer=1 filter=204 channel=58
    -26, -153, -35, -116, -200, -71, -58, -124, -58,
    -- layer=1 filter=204 channel=59
    -10, -9, -17, -8, -10, -3, 5, -2, 5,
    -- layer=1 filter=204 channel=60
    14, 3, 8, 13, 4, 9, 20, 4, 11,
    -- layer=1 filter=204 channel=61
    -3, -8, -10, -1, 7, -1, -5, 0, -2,
    -- layer=1 filter=204 channel=62
    31, -1, 29, 25, 13, 4, 14, 34, 22,
    -- layer=1 filter=204 channel=63
    11, 23, 6, -6, 11, 19, -24, -21, -5,
    -- layer=1 filter=204 channel=64
    -9, -19, -32, -2, -4, -1, 5, 6, 1,
    -- layer=1 filter=204 channel=65
    7, 5, -2, 15, -1, -1, 11, 18, 9,
    -- layer=1 filter=204 channel=66
    12, 2, 14, -5, -3, 1, -29, -5, -13,
    -- layer=1 filter=204 channel=67
    -17, -12, -45, -6, -2, -16, -2, 8, -2,
    -- layer=1 filter=204 channel=68
    -57, -40, -44, -32, -82, -98, -62, -74, -50,
    -- layer=1 filter=204 channel=69
    8, 3, 13, 16, -1, 8, 14, 15, 14,
    -- layer=1 filter=204 channel=70
    -26, -33, -32, -13, -1, -10, 20, 25, 47,
    -- layer=1 filter=204 channel=71
    14, 12, -1, 20, 19, 27, 20, 24, 15,
    -- layer=1 filter=204 channel=72
    -2, -15, 15, 8, 4, 16, 55, 8, 39,
    -- layer=1 filter=204 channel=73
    -1, 3, -2, -11, -4, 1, 0, 4, -6,
    -- layer=1 filter=204 channel=74
    -9, -9, -34, -4, 1, -43, 24, -5, 9,
    -- layer=1 filter=204 channel=75
    -29, -36, -25, -37, 0, 15, 25, 32, 45,
    -- layer=1 filter=204 channel=76
    12, 0, 7, 13, -6, -27, 11, -4, 6,
    -- layer=1 filter=204 channel=77
    -14, 14, -3, 6, 13, 0, 4, 6, 0,
    -- layer=1 filter=204 channel=78
    -1, 3, -15, -15, -8, -2, 0, -15, -23,
    -- layer=1 filter=204 channel=79
    29, 2, 20, 22, 1, 3, 11, 19, 9,
    -- layer=1 filter=204 channel=80
    8, -12, 8, -1, 0, 2, -8, 0, 6,
    -- layer=1 filter=204 channel=81
    2, 1, 15, 14, 22, 10, 7, 21, 23,
    -- layer=1 filter=204 channel=82
    -12, -5, -9, 13, 14, 1, 22, 29, 17,
    -- layer=1 filter=204 channel=83
    8, -12, 24, 20, 1, -17, 24, 22, 25,
    -- layer=1 filter=204 channel=84
    19, 22, 26, 35, 26, 15, 25, 39, 59,
    -- layer=1 filter=204 channel=85
    11, -63, -15, -49, -93, -43, -32, -95, -45,
    -- layer=1 filter=204 channel=86
    5, 7, 16, -6, 10, 3, -26, -21, -14,
    -- layer=1 filter=204 channel=87
    20, -14, -6, 29, 25, 8, 55, 59, 24,
    -- layer=1 filter=204 channel=88
    -3, 1, 2, 0, 0, 3, 12, 3, 20,
    -- layer=1 filter=204 channel=89
    5, 10, -13, 19, 24, 5, 13, 15, 22,
    -- layer=1 filter=204 channel=90
    -45, -55, -65, -31, -74, -80, -45, -35, -55,
    -- layer=1 filter=204 channel=91
    0, -7, -20, 1, -3, -2, 37, 24, 23,
    -- layer=1 filter=204 channel=92
    -50, -5, -3, -30, -30, -40, 18, -12, -30,
    -- layer=1 filter=204 channel=93
    11, 8, 14, 17, 20, 20, 15, 11, 13,
    -- layer=1 filter=204 channel=94
    -10, 0, 6, -8, -5, -5, -22, -9, -21,
    -- layer=1 filter=204 channel=95
    22, 23, 13, 30, 16, 20, 25, 45, 56,
    -- layer=1 filter=204 channel=96
    0, -6, 4, -2, 4, 0, -12, 3, 11,
    -- layer=1 filter=204 channel=97
    10, 9, 13, 12, -6, 8, 0, 3, -12,
    -- layer=1 filter=204 channel=98
    -9, -13, 2, 25, -8, -17, 25, 14, 21,
    -- layer=1 filter=204 channel=99
    -49, -49, -48, -34, -82, -81, 11, -77, -84,
    -- layer=1 filter=204 channel=100
    3, 10, 9, -23, -18, 1, -30, -28, -25,
    -- layer=1 filter=204 channel=101
    -9, -12, -26, 20, 12, 1, 33, 14, 20,
    -- layer=1 filter=204 channel=102
    -9, -1, -24, 0, -25, -3, 13, -8, -15,
    -- layer=1 filter=204 channel=103
    -10, 1, 2, 6, 0, 22, -31, -20, -2,
    -- layer=1 filter=204 channel=104
    41, -26, 0, -26, -6, -28, -26, -10, -14,
    -- layer=1 filter=204 channel=105
    11, 3, 19, 6, 0, 12, -1, -16, -17,
    -- layer=1 filter=204 channel=106
    -12, -3, -23, 22, -1, -18, 25, 23, 31,
    -- layer=1 filter=204 channel=107
    -1, 3, 4, -2, 12, -11, -7, 0, 3,
    -- layer=1 filter=204 channel=108
    -25, -43, -32, -11, -80, -89, -24, -43, -53,
    -- layer=1 filter=204 channel=109
    0, 6, 9, -3, 3, 5, 7, 0, 2,
    -- layer=1 filter=204 channel=110
    10, 4, 2, -7, 0, -4, -4, 1, -14,
    -- layer=1 filter=204 channel=111
    18, 18, 21, 30, 12, 21, 47, 41, 28,
    -- layer=1 filter=204 channel=112
    9, 32, 15, 36, 27, 37, -3, 26, 55,
    -- layer=1 filter=204 channel=113
    -27, -32, -5, -12, -28, 5, 33, 28, 23,
    -- layer=1 filter=204 channel=114
    16, 18, 28, -2, 13, -11, 12, 7, 13,
    -- layer=1 filter=204 channel=115
    -3, 4, 15, -12, -17, 8, -14, -38, -14,
    -- layer=1 filter=204 channel=116
    -11, -3, 0, -4, -6, 5, -9, 4, -2,
    -- layer=1 filter=204 channel=117
    60, 25, 48, 85, 55, 63, 43, 53, 51,
    -- layer=1 filter=204 channel=118
    33, 22, 4, 34, 9, 8, 56, 36, 48,
    -- layer=1 filter=204 channel=119
    -22, -32, -11, -32, -84, -95, -41, -63, -54,
    -- layer=1 filter=204 channel=120
    -10, -8, -2, 12, -11, -9, 9, 21, 10,
    -- layer=1 filter=204 channel=121
    24, 15, 7, 18, 36, 35, 52, 50, 5,
    -- layer=1 filter=204 channel=122
    -9, 7, -4, 8, -3, -2, 7, 0, -9,
    -- layer=1 filter=204 channel=123
    12, 16, 19, 5, 17, 20, 7, 10, 21,
    -- layer=1 filter=204 channel=124
    -7, -4, -13, -11, -10, 10, -8, 3, -3,
    -- layer=1 filter=204 channel=125
    -46, -21, -51, -19, -5, -1, 42, 29, 38,
    -- layer=1 filter=204 channel=126
    -8, -11, -6, 71, 25, -3, 49, 62, 49,
    -- layer=1 filter=204 channel=127
    26, 23, 7, 29, 27, 29, 49, 35, 52,
    -- layer=1 filter=205 channel=0
    2, 4, 1, 1, -4, 3, -2, 3, -2,
    -- layer=1 filter=205 channel=1
    2, 6, -4, 2, 4, -10, 1, 0, 4,
    -- layer=1 filter=205 channel=2
    2, 5, -1, -1, 1, 2, -6, -4, 4,
    -- layer=1 filter=205 channel=3
    3, -2, 5, -1, -1, -3, -8, -6, 5,
    -- layer=1 filter=205 channel=4
    4, 0, -4, -11, -3, -5, -12, -7, 8,
    -- layer=1 filter=205 channel=5
    -10, 0, -4, 2, 7, -1, -12, 6, 2,
    -- layer=1 filter=205 channel=6
    8, -9, 3, -10, -4, 4, 3, -10, -4,
    -- layer=1 filter=205 channel=7
    -6, -9, 6, 1, -6, 9, 7, -4, -1,
    -- layer=1 filter=205 channel=8
    -3, -10, -1, 7, 3, -10, -2, 4, 5,
    -- layer=1 filter=205 channel=9
    -1, -4, -5, 7, -11, -4, -2, 7, 4,
    -- layer=1 filter=205 channel=10
    -4, 6, -12, -2, -5, 0, 0, -6, 3,
    -- layer=1 filter=205 channel=11
    -6, 6, -8, -7, -8, -7, 1, -4, -7,
    -- layer=1 filter=205 channel=12
    -6, 6, 4, -1, 7, 9, 3, -3, -6,
    -- layer=1 filter=205 channel=13
    -8, -9, 6, 1, -1, 0, 0, 8, 4,
    -- layer=1 filter=205 channel=14
    7, 3, 0, -4, 9, -8, 3, -10, 0,
    -- layer=1 filter=205 channel=15
    -4, -6, -1, 0, -9, -5, -10, -12, 8,
    -- layer=1 filter=205 channel=16
    -4, -1, 5, -2, -5, -5, 4, 0, 6,
    -- layer=1 filter=205 channel=17
    7, 3, 2, 3, -4, -12, -8, 8, 6,
    -- layer=1 filter=205 channel=18
    -7, 7, -5, 0, -7, -10, -4, 7, 9,
    -- layer=1 filter=205 channel=19
    6, -1, -13, 0, -3, -7, -6, 1, 7,
    -- layer=1 filter=205 channel=20
    -5, -11, 0, -9, 8, 1, 6, -2, -10,
    -- layer=1 filter=205 channel=21
    6, -9, 4, 5, -9, 2, -3, 0, -10,
    -- layer=1 filter=205 channel=22
    -10, 4, -4, -4, 0, -1, 7, 1, -1,
    -- layer=1 filter=205 channel=23
    -8, -2, -4, -12, -11, 2, 1, -9, -7,
    -- layer=1 filter=205 channel=24
    8, -7, 7, -11, -5, 0, -10, 3, 6,
    -- layer=1 filter=205 channel=25
    0, -6, -3, -5, 3, 7, 5, -6, -10,
    -- layer=1 filter=205 channel=26
    -11, 8, -5, 0, -2, 1, 0, -11, -6,
    -- layer=1 filter=205 channel=27
    0, -5, 7, 2, -8, -8, 2, -9, -8,
    -- layer=1 filter=205 channel=28
    -12, 2, 2, -2, 0, 1, 1, -10, 0,
    -- layer=1 filter=205 channel=29
    3, -2, -5, 5, 7, -5, 4, 0, 4,
    -- layer=1 filter=205 channel=30
    7, 2, -7, -4, -5, 2, 10, -2, -12,
    -- layer=1 filter=205 channel=31
    -2, -3, 0, -11, 0, -8, 7, 4, -8,
    -- layer=1 filter=205 channel=32
    2, -3, 0, 0, -1, 6, -2, 0, -2,
    -- layer=1 filter=205 channel=33
    -2, 4, -5, -8, 5, 3, 4, -3, 11,
    -- layer=1 filter=205 channel=34
    -10, -1, 5, 5, -10, 0, -1, -5, -3,
    -- layer=1 filter=205 channel=35
    -7, -10, -12, 6, 7, 3, -13, 2, -3,
    -- layer=1 filter=205 channel=36
    6, -11, -7, -5, -7, -1, 0, 8, 5,
    -- layer=1 filter=205 channel=37
    2, -3, 6, -1, -3, -1, 0, 9, -6,
    -- layer=1 filter=205 channel=38
    -4, -8, 9, 2, -4, 0, 2, 5, 2,
    -- layer=1 filter=205 channel=39
    -4, -10, 4, 7, -9, -8, 0, -7, 1,
    -- layer=1 filter=205 channel=40
    4, 2, 1, -8, 0, -1, -5, 4, 0,
    -- layer=1 filter=205 channel=41
    -2, -9, 3, -5, -13, 6, 2, 4, 3,
    -- layer=1 filter=205 channel=42
    -6, 6, 1, 5, 10, -6, -10, -7, -6,
    -- layer=1 filter=205 channel=43
    0, 0, -2, 4, 7, -1, -1, -8, -9,
    -- layer=1 filter=205 channel=44
    0, -5, 1, 5, -3, -5, 7, 0, 4,
    -- layer=1 filter=205 channel=45
    -4, 7, -8, 9, 0, -6, -9, 8, -7,
    -- layer=1 filter=205 channel=46
    -2, -1, 1, 1, -7, -9, 0, 3, 5,
    -- layer=1 filter=205 channel=47
    10, -11, 4, 4, 0, 1, 8, -1, 0,
    -- layer=1 filter=205 channel=48
    -1, -6, 2, -9, 4, -7, 5, -2, -5,
    -- layer=1 filter=205 channel=49
    -6, 8, 2, -5, 0, 5, -3, -4, 1,
    -- layer=1 filter=205 channel=50
    -3, -10, -11, -12, 0, -11, 8, 5, -6,
    -- layer=1 filter=205 channel=51
    -8, -7, 4, -1, 3, -9, 7, 2, -5,
    -- layer=1 filter=205 channel=52
    -1, -2, -6, 5, -2, -4, -5, -7, -6,
    -- layer=1 filter=205 channel=53
    -12, -5, 0, -11, -8, 7, 3, -4, 2,
    -- layer=1 filter=205 channel=54
    -2, 3, 3, 2, -7, -6, 5, -7, -6,
    -- layer=1 filter=205 channel=55
    -6, -8, -1, -3, -4, -2, 1, -9, 0,
    -- layer=1 filter=205 channel=56
    -7, 1, -5, 5, -12, 4, 2, 7, -8,
    -- layer=1 filter=205 channel=57
    1, 0, -9, 0, 5, -2, -11, 5, -3,
    -- layer=1 filter=205 channel=58
    -4, 3, 4, -9, -5, -1, -4, -10, -5,
    -- layer=1 filter=205 channel=59
    5, -2, -7, -3, 8, 4, -6, -4, -2,
    -- layer=1 filter=205 channel=60
    6, 8, -5, -3, 3, 4, 1, 2, 8,
    -- layer=1 filter=205 channel=61
    0, -8, 0, -1, -8, -2, 5, 4, 2,
    -- layer=1 filter=205 channel=62
    -2, 7, -4, 8, 5, 2, -1, -8, -9,
    -- layer=1 filter=205 channel=63
    -12, -11, 2, 5, 6, 7, -2, 0, -3,
    -- layer=1 filter=205 channel=64
    1, -5, -1, 8, 0, -6, -12, -9, -12,
    -- layer=1 filter=205 channel=65
    1, 0, -2, 5, 1, 0, -1, -1, 6,
    -- layer=1 filter=205 channel=66
    -4, -13, -2, 8, -7, -4, -11, -11, -4,
    -- layer=1 filter=205 channel=67
    3, -11, -3, -9, -9, 4, -10, 1, 4,
    -- layer=1 filter=205 channel=68
    -9, -4, 7, 7, 2, -11, 0, -11, -7,
    -- layer=1 filter=205 channel=69
    7, -4, 6, 5, -7, 1, 7, -4, -5,
    -- layer=1 filter=205 channel=70
    9, -4, -7, 1, -4, -3, 1, 8, 1,
    -- layer=1 filter=205 channel=71
    5, 8, -1, 4, 4, -12, 5, 1, -2,
    -- layer=1 filter=205 channel=72
    0, 4, -10, -7, -11, 4, -6, -6, -1,
    -- layer=1 filter=205 channel=73
    -11, -9, 4, -3, 8, -8, 4, 4, 5,
    -- layer=1 filter=205 channel=74
    0, -11, -6, -8, -8, 1, -4, 5, 7,
    -- layer=1 filter=205 channel=75
    7, 6, -4, -4, -1, 9, 0, 5, 0,
    -- layer=1 filter=205 channel=76
    -4, 3, 0, 7, 4, -12, 4, 1, -6,
    -- layer=1 filter=205 channel=77
    -3, -12, -6, 5, -5, -12, -12, -1, -7,
    -- layer=1 filter=205 channel=78
    -9, 2, -4, -8, -4, -7, 2, -9, -9,
    -- layer=1 filter=205 channel=79
    7, -9, 4, 4, 5, -8, 7, -3, -11,
    -- layer=1 filter=205 channel=80
    -9, 8, -7, -10, -6, 8, -10, -9, 6,
    -- layer=1 filter=205 channel=81
    0, 0, -1, 4, 7, -7, 7, 0, 0,
    -- layer=1 filter=205 channel=82
    6, -5, 2, 1, 6, -8, -11, -6, -5,
    -- layer=1 filter=205 channel=83
    7, 2, -7, -2, -3, 6, 1, 6, -7,
    -- layer=1 filter=205 channel=84
    -11, -1, 0, -7, 0, -4, -1, -9, -6,
    -- layer=1 filter=205 channel=85
    3, 5, 0, 0, -6, 7, -4, -2, -6,
    -- layer=1 filter=205 channel=86
    -8, -7, 4, -3, -9, -10, -5, -6, 6,
    -- layer=1 filter=205 channel=87
    -1, 0, -5, -10, -12, 5, 8, -1, 5,
    -- layer=1 filter=205 channel=88
    -4, 3, 1, 5, -7, -8, -3, 4, 2,
    -- layer=1 filter=205 channel=89
    4, 7, 4, -2, -4, 1, -2, -3, 0,
    -- layer=1 filter=205 channel=90
    -6, 0, -6, -9, -2, -1, 0, 0, -3,
    -- layer=1 filter=205 channel=91
    0, 8, -6, -7, -1, -3, 4, 3, 1,
    -- layer=1 filter=205 channel=92
    0, 1, 1, 7, -9, 1, -7, -4, 4,
    -- layer=1 filter=205 channel=93
    -7, 0, 7, -1, 5, 3, 8, -3, 6,
    -- layer=1 filter=205 channel=94
    -1, 2, -2, -11, -2, 0, -4, 3, -3,
    -- layer=1 filter=205 channel=95
    -3, -9, -10, 3, -10, 1, -6, 0, -8,
    -- layer=1 filter=205 channel=96
    1, 0, 6, -9, -10, 3, 5, 5, 3,
    -- layer=1 filter=205 channel=97
    6, -4, 4, -1, 4, 5, 5, 6, -4,
    -- layer=1 filter=205 channel=98
    -2, 4, -5, -13, 0, 0, 3, -8, 9,
    -- layer=1 filter=205 channel=99
    -4, 5, -6, 1, -6, -12, 4, -11, -5,
    -- layer=1 filter=205 channel=100
    -1, -12, 6, -12, -8, 5, 5, 0, -10,
    -- layer=1 filter=205 channel=101
    -9, -9, -4, -8, -2, 7, -11, -6, -12,
    -- layer=1 filter=205 channel=102
    -3, -1, 7, -11, -8, -12, -12, -8, 3,
    -- layer=1 filter=205 channel=103
    -9, -10, -12, -4, -12, -8, 3, -8, 2,
    -- layer=1 filter=205 channel=104
    -13, -5, 2, -3, -8, 1, 2, 1, -2,
    -- layer=1 filter=205 channel=105
    -12, -3, 0, 1, 0, -4, -2, -6, 6,
    -- layer=1 filter=205 channel=106
    -6, -9, -11, 2, 2, -9, -4, 1, 9,
    -- layer=1 filter=205 channel=107
    5, -10, -7, 2, -1, 1, -3, 8, -11,
    -- layer=1 filter=205 channel=108
    1, 4, 7, -1, 5, 1, -8, 8, 2,
    -- layer=1 filter=205 channel=109
    -3, -5, -9, -7, 4, 1, -4, -9, 7,
    -- layer=1 filter=205 channel=110
    -7, 3, 2, -1, 7, 1, 0, -7, 0,
    -- layer=1 filter=205 channel=111
    2, 9, 0, -12, -12, 1, 1, -2, -8,
    -- layer=1 filter=205 channel=112
    0, -5, 3, 7, 3, -3, 0, 3, 0,
    -- layer=1 filter=205 channel=113
    -7, 6, 6, -2, 12, 11, -6, 8, 0,
    -- layer=1 filter=205 channel=114
    10, 3, -8, -7, 8, -7, -8, -4, 7,
    -- layer=1 filter=205 channel=115
    0, -7, 2, 3, 2, 1, -6, 6, -2,
    -- layer=1 filter=205 channel=116
    8, 5, 0, -9, 9, -4, -1, -4, -2,
    -- layer=1 filter=205 channel=117
    -11, 3, -8, 3, -2, 5, -9, -9, 9,
    -- layer=1 filter=205 channel=118
    -7, 0, -7, 1, -1, -3, -2, 3, 8,
    -- layer=1 filter=205 channel=119
    5, -9, -9, -2, -1, 1, -7, 5, 3,
    -- layer=1 filter=205 channel=120
    6, -5, 2, -12, 0, 2, 0, 2, 5,
    -- layer=1 filter=205 channel=121
    -2, 6, 2, -2, 1, -6, 0, 0, 6,
    -- layer=1 filter=205 channel=122
    -3, -8, 3, 5, 0, 0, -4, -6, 7,
    -- layer=1 filter=205 channel=123
    5, 3, 8, -9, 8, -6, -5, -10, -5,
    -- layer=1 filter=205 channel=124
    4, -11, -10, 9, 0, 8, -6, -9, -7,
    -- layer=1 filter=205 channel=125
    5, 7, -11, -11, -2, -9, -5, -6, -7,
    -- layer=1 filter=205 channel=126
    2, 1, 4, -4, -9, 0, 7, -1, -7,
    -- layer=1 filter=205 channel=127
    4, -5, 3, 1, -6, -6, 4, 2, 8,
    -- layer=1 filter=206 channel=0
    -9, 3, -12, -4, -8, 0, 2, -2, -10,
    -- layer=1 filter=206 channel=1
    -2, 0, 2, 3, -9, -10, 2, 6, 6,
    -- layer=1 filter=206 channel=2
    1, 11, -4, -12, 10, -10, -2, 5, -4,
    -- layer=1 filter=206 channel=3
    -6, 5, 0, -9, -1, -1, 9, 1, 2,
    -- layer=1 filter=206 channel=4
    2, -7, -9, -9, 3, 5, -5, 2, -3,
    -- layer=1 filter=206 channel=5
    -11, 0, 3, 7, -2, 0, -18, 1, -14,
    -- layer=1 filter=206 channel=6
    3, 3, 8, -5, -3, -3, -12, -13, -8,
    -- layer=1 filter=206 channel=7
    -6, 3, 0, -9, 5, -4, -17, 6, 8,
    -- layer=1 filter=206 channel=8
    -12, 0, -4, -12, -8, 5, -5, -8, -9,
    -- layer=1 filter=206 channel=9
    8, -9, -9, -5, -9, 0, 1, -3, 0,
    -- layer=1 filter=206 channel=10
    4, 0, -11, 0, 7, 0, -5, 1, 1,
    -- layer=1 filter=206 channel=11
    -6, 1, -3, -7, -10, -7, -5, -2, -13,
    -- layer=1 filter=206 channel=12
    6, 1, -7, -9, 6, -7, -4, 9, -6,
    -- layer=1 filter=206 channel=13
    4, -12, 4, 0, -4, -7, -9, -12, -4,
    -- layer=1 filter=206 channel=14
    6, 5, -13, -1, 6, 3, 10, 8, -1,
    -- layer=1 filter=206 channel=15
    -1, 3, -7, 9, -4, -7, 10, 5, -5,
    -- layer=1 filter=206 channel=16
    -9, -2, 1, 5, 0, 1, 0, 1, -2,
    -- layer=1 filter=206 channel=17
    -7, -1, -4, 2, -12, -5, 2, -12, 1,
    -- layer=1 filter=206 channel=18
    5, 3, -9, 2, 3, -6, -9, -2, 6,
    -- layer=1 filter=206 channel=19
    -2, -9, -8, 7, 7, -10, -4, 5, 7,
    -- layer=1 filter=206 channel=20
    -4, 1, -8, -3, -1, -6, -4, 0, -6,
    -- layer=1 filter=206 channel=21
    -8, 1, -6, 5, -4, 1, 0, 1, -11,
    -- layer=1 filter=206 channel=22
    0, -8, 8, 3, 5, 6, -7, 4, 7,
    -- layer=1 filter=206 channel=23
    4, 3, 1, -7, -4, -2, -17, -5, 3,
    -- layer=1 filter=206 channel=24
    6, -1, -12, 2, 0, -3, 1, 3, 4,
    -- layer=1 filter=206 channel=25
    -9, -9, -13, -3, -3, -3, 1, -14, 1,
    -- layer=1 filter=206 channel=26
    -12, 2, -16, 2, -6, 2, -12, 2, 8,
    -- layer=1 filter=206 channel=27
    0, -7, 1, -9, -9, -5, -3, -6, -10,
    -- layer=1 filter=206 channel=28
    -9, 0, -13, -1, -12, -2, 5, -4, -7,
    -- layer=1 filter=206 channel=29
    -5, 0, 0, -13, -3, 4, -7, -2, 8,
    -- layer=1 filter=206 channel=30
    5, -9, 12, -6, 3, 3, -2, -2, 19,
    -- layer=1 filter=206 channel=31
    -1, 2, 4, 4, 2, 5, -9, 5, -2,
    -- layer=1 filter=206 channel=32
    6, 8, -10, -9, 0, 0, -1, -9, -3,
    -- layer=1 filter=206 channel=33
    6, 3, 0, 1, -8, 1, 4, 5, 8,
    -- layer=1 filter=206 channel=34
    -6, 8, 7, -11, -2, 5, 6, 2, 0,
    -- layer=1 filter=206 channel=35
    -9, -4, 8, -11, 1, -7, -2, -9, 6,
    -- layer=1 filter=206 channel=36
    -5, 0, 0, -5, 3, -9, -4, -9, -4,
    -- layer=1 filter=206 channel=37
    0, -10, -10, 8, 9, -5, -7, -11, 2,
    -- layer=1 filter=206 channel=38
    -8, -9, -3, -1, -5, 6, 5, -8, 10,
    -- layer=1 filter=206 channel=39
    -5, 4, -13, 3, -8, -6, 3, -1, -3,
    -- layer=1 filter=206 channel=40
    5, -7, -3, 5, -7, 6, -12, 0, 8,
    -- layer=1 filter=206 channel=41
    7, 0, 5, 1, -9, 4, 8, -8, 1,
    -- layer=1 filter=206 channel=42
    -2, 4, 4, -9, 3, 7, -6, 5, 7,
    -- layer=1 filter=206 channel=43
    8, -10, -11, 0, 4, -8, -7, -3, 4,
    -- layer=1 filter=206 channel=44
    -15, 1, 1, -13, 7, -8, 3, 3, 4,
    -- layer=1 filter=206 channel=45
    5, -7, 2, 0, -11, -3, -1, 0, 3,
    -- layer=1 filter=206 channel=46
    -3, 3, -12, -9, 6, 2, -10, 4, -12,
    -- layer=1 filter=206 channel=47
    -1, 1, -6, -4, -6, -10, -10, 5, 0,
    -- layer=1 filter=206 channel=48
    -11, 0, -3, 0, 3, 4, 7, -3, 7,
    -- layer=1 filter=206 channel=49
    0, -13, -7, 3, -7, 2, -10, 6, -7,
    -- layer=1 filter=206 channel=50
    -8, -2, -3, -5, -2, 2, 4, 3, -4,
    -- layer=1 filter=206 channel=51
    -6, -6, 3, -8, 6, -6, -12, -4, 3,
    -- layer=1 filter=206 channel=52
    7, 10, -9, 1, -10, 10, 0, -5, 1,
    -- layer=1 filter=206 channel=53
    0, 0, -6, -3, -9, -4, 2, -3, 4,
    -- layer=1 filter=206 channel=54
    -10, 4, -16, -2, -7, -10, 2, 5, -2,
    -- layer=1 filter=206 channel=55
    -5, -12, -13, -17, -8, -11, -14, -8, -13,
    -- layer=1 filter=206 channel=56
    -4, 5, 3, -1, -5, -7, -10, -3, 7,
    -- layer=1 filter=206 channel=57
    0, -1, 5, 2, -6, -3, 6, -14, 3,
    -- layer=1 filter=206 channel=58
    -16, 2, -14, -14, -5, -9, 0, -14, 7,
    -- layer=1 filter=206 channel=59
    0, -2, -5, -5, 1, 3, 6, -8, -5,
    -- layer=1 filter=206 channel=60
    -11, 7, 4, 9, -2, 5, 2, -8, 0,
    -- layer=1 filter=206 channel=61
    5, 2, 2, -1, 0, -8, 7, 0, -5,
    -- layer=1 filter=206 channel=62
    6, -12, -13, -9, -7, 0, -12, -9, -6,
    -- layer=1 filter=206 channel=63
    -4, 3, -11, -9, 0, 5, 0, 4, -5,
    -- layer=1 filter=206 channel=64
    -8, -10, -8, -9, 4, -2, 6, -11, 0,
    -- layer=1 filter=206 channel=65
    5, 4, 2, 6, -11, -5, 0, -3, 0,
    -- layer=1 filter=206 channel=66
    4, 3, 4, 1, 1, -4, -1, -16, -8,
    -- layer=1 filter=206 channel=67
    7, -5, 1, -2, 4, -3, -2, 1, 0,
    -- layer=1 filter=206 channel=68
    -14, -3, -5, -13, -3, -7, 0, 8, -8,
    -- layer=1 filter=206 channel=69
    -3, -15, -17, -2, -4, -6, -10, 0, -13,
    -- layer=1 filter=206 channel=70
    5, 6, -6, -4, -1, -2, -6, 5, 14,
    -- layer=1 filter=206 channel=71
    4, -13, -7, -1, -13, -13, -4, 1, -9,
    -- layer=1 filter=206 channel=72
    -8, 0, -5, 0, -2, 0, 1, -9, -3,
    -- layer=1 filter=206 channel=73
    -7, 6, -4, -9, -8, -9, -11, 5, 6,
    -- layer=1 filter=206 channel=74
    -3, 1, 4, -12, -9, 7, -7, 3, -4,
    -- layer=1 filter=206 channel=75
    -11, -1, 7, 4, 8, -10, -9, 0, 11,
    -- layer=1 filter=206 channel=76
    2, 2, 5, -13, -11, -5, 2, 2, 1,
    -- layer=1 filter=206 channel=77
    -5, 7, -10, -8, -11, -12, -7, 0, -8,
    -- layer=1 filter=206 channel=78
    -2, 4, -2, -1, 7, -8, 7, 5, -12,
    -- layer=1 filter=206 channel=79
    6, -4, 4, -8, 0, 0, -4, -4, -1,
    -- layer=1 filter=206 channel=80
    4, 6, 0, -7, 5, 1, 8, 2, 3,
    -- layer=1 filter=206 channel=81
    0, -7, -3, 1, -7, -12, -13, 2, -14,
    -- layer=1 filter=206 channel=82
    -9, -12, 5, -10, 0, -4, -4, -8, -12,
    -- layer=1 filter=206 channel=83
    7, 3, 0, 6, -7, -6, 2, -6, -2,
    -- layer=1 filter=206 channel=84
    -4, -2, 9, -2, -4, -10, 7, 7, -2,
    -- layer=1 filter=206 channel=85
    4, 2, 4, -5, 3, 2, -7, 0, -10,
    -- layer=1 filter=206 channel=86
    4, -10, 5, 6, 0, -3, 0, 0, -2,
    -- layer=1 filter=206 channel=87
    -3, 10, 5, -11, 0, -10, -2, -2, 3,
    -- layer=1 filter=206 channel=88
    9, -2, -2, 3, -3, -5, 1, -7, 1,
    -- layer=1 filter=206 channel=89
    1, -8, 8, 6, -8, 7, 5, -8, 4,
    -- layer=1 filter=206 channel=90
    -12, 6, -11, 5, 8, 5, -8, 0, -9,
    -- layer=1 filter=206 channel=91
    -7, -10, -4, 0, -5, 0, 3, -5, -7,
    -- layer=1 filter=206 channel=92
    1, -7, 1, 0, -2, 5, 6, -11, -8,
    -- layer=1 filter=206 channel=93
    -5, -12, 0, 0, 2, -1, 5, 3, -3,
    -- layer=1 filter=206 channel=94
    4, -8, -6, -4, 6, -3, -12, -1, -2,
    -- layer=1 filter=206 channel=95
    -13, 1, 0, -12, -4, -5, -6, 12, 11,
    -- layer=1 filter=206 channel=96
    -11, 2, -5, 7, -7, -1, 0, 1, -6,
    -- layer=1 filter=206 channel=97
    4, 6, -6, -10, -8, -5, 5, 1, 1,
    -- layer=1 filter=206 channel=98
    2, 8, 7, -2, -16, 6, -12, -16, -3,
    -- layer=1 filter=206 channel=99
    0, 4, 0, -12, -11, -6, 7, -1, 7,
    -- layer=1 filter=206 channel=100
    -3, -12, 5, -1, 7, 0, 4, -10, -8,
    -- layer=1 filter=206 channel=101
    -7, 1, 3, -8, -2, 5, -4, -11, 3,
    -- layer=1 filter=206 channel=102
    6, -7, -6, 0, 1, -9, -10, -1, -3,
    -- layer=1 filter=206 channel=103
    -11, -15, 6, 5, -15, -11, 8, -14, -11,
    -- layer=1 filter=206 channel=104
    -1, 3, -9, 8, 5, -4, 0, -9, -5,
    -- layer=1 filter=206 channel=105
    -14, 2, -6, -10, -5, -6, -6, -13, -9,
    -- layer=1 filter=206 channel=106
    -11, 3, -8, -11, -2, -5, -1, 13, 3,
    -- layer=1 filter=206 channel=107
    -6, -9, 1, -9, -4, 6, 4, 6, 2,
    -- layer=1 filter=206 channel=108
    -6, -8, -9, -10, 3, -11, 9, -5, 3,
    -- layer=1 filter=206 channel=109
    8, 3, 3, -3, 2, 6, -7, -4, 10,
    -- layer=1 filter=206 channel=110
    -5, 3, -4, 2, -1, 5, -2, -13, -1,
    -- layer=1 filter=206 channel=111
    -14, -1, 12, -12, -9, -7, -7, 8, 0,
    -- layer=1 filter=206 channel=112
    -10, 0, 8, -10, -4, -1, -3, 5, 2,
    -- layer=1 filter=206 channel=113
    -4, -13, -4, -7, 0, 0, 3, 6, 2,
    -- layer=1 filter=206 channel=114
    -14, 5, 5, 4, -2, 5, -14, 0, -15,
    -- layer=1 filter=206 channel=115
    2, 3, 0, 2, -6, -12, 3, -6, -7,
    -- layer=1 filter=206 channel=116
    4, 3, 8, 6, 0, -2, -1, 1, 0,
    -- layer=1 filter=206 channel=117
    -3, 0, 1, 3, 9, -9, -10, 5, -12,
    -- layer=1 filter=206 channel=118
    -2, -2, 11, -7, 6, -2, 2, 0, 8,
    -- layer=1 filter=206 channel=119
    -6, -15, -6, 3, -9, -4, 0, -2, 6,
    -- layer=1 filter=206 channel=120
    7, -14, -3, -1, -2, -2, -11, -14, -8,
    -- layer=1 filter=206 channel=121
    -1, -2, -12, 2, -16, -7, 4, 2, 0,
    -- layer=1 filter=206 channel=122
    2, 7, 4, -2, 4, 7, -7, -9, -7,
    -- layer=1 filter=206 channel=123
    -4, -6, -14, -16, -5, -12, 1, -8, -5,
    -- layer=1 filter=206 channel=124
    4, 1, 1, -8, -11, -5, -9, -4, -9,
    -- layer=1 filter=206 channel=125
    0, 6, -3, -8, 2, 8, 6, 4, 11,
    -- layer=1 filter=206 channel=126
    -8, 9, 6, -9, -15, 0, 7, 2, -6,
    -- layer=1 filter=206 channel=127
    0, 2, 1, -13, -8, -1, 10, 16, 14,
    -- layer=1 filter=207 channel=0
    -15, -7, 0, -2, -4, 1, -9, -13, 1,
    -- layer=1 filter=207 channel=1
    5, -18, -10, 0, 0, -5, -6, -10, 0,
    -- layer=1 filter=207 channel=2
    1, -2, -16, 0, 6, -2, 0, 0, -5,
    -- layer=1 filter=207 channel=3
    1, 0, 1, 2, 3, -2, 1, -5, 6,
    -- layer=1 filter=207 channel=4
    -9, 3, 6, -11, -12, 8, -7, -8, 8,
    -- layer=1 filter=207 channel=5
    1, -1, -8, -24, -23, -22, -19, -9, -23,
    -- layer=1 filter=207 channel=6
    -17, -25, -14, 9, -15, -3, -17, -21, -19,
    -- layer=1 filter=207 channel=7
    0, -12, -6, -16, -13, -23, -8, -19, -9,
    -- layer=1 filter=207 channel=8
    -6, -7, -6, -10, -22, -15, -15, -4, -12,
    -- layer=1 filter=207 channel=9
    -6, -1, -18, -15, -6, -5, -10, -15, -6,
    -- layer=1 filter=207 channel=10
    -17, -3, -1, -13, -18, -10, 0, -22, -15,
    -- layer=1 filter=207 channel=11
    6, 5, -7, 0, 7, -5, -3, 10, 8,
    -- layer=1 filter=207 channel=12
    3, -11, 0, -21, 18, 2, 9, 3, -13,
    -- layer=1 filter=207 channel=13
    -3, -13, -15, -8, 1, -11, -4, -8, -5,
    -- layer=1 filter=207 channel=14
    -14, 0, 2, -13, 10, -10, -10, -10, -3,
    -- layer=1 filter=207 channel=15
    -12, -6, -26, -15, -14, -17, 1, -16, -18,
    -- layer=1 filter=207 channel=16
    -7, -17, -22, -8, -11, -23, -6, -18, -8,
    -- layer=1 filter=207 channel=17
    -6, 7, -8, -8, -11, 2, 5, 2, -3,
    -- layer=1 filter=207 channel=18
    7, -1, -1, 1, -3, -4, -14, 1, 2,
    -- layer=1 filter=207 channel=19
    -12, -10, -12, -7, -6, -15, -11, 0, -8,
    -- layer=1 filter=207 channel=20
    -11, -14, -8, -6, 0, -8, 4, -4, -10,
    -- layer=1 filter=207 channel=21
    -16, -15, -15, -8, -23, -9, -20, -17, -16,
    -- layer=1 filter=207 channel=22
    -6, -11, -11, -2, 1, -7, 3, -6, 0,
    -- layer=1 filter=207 channel=23
    -16, -13, -16, -3, -22, -12, -24, -16, -9,
    -- layer=1 filter=207 channel=24
    -6, 1, -1, -2, -14, -17, -1, -2, -4,
    -- layer=1 filter=207 channel=25
    -11, -8, -17, -24, -19, -20, 3, -10, -5,
    -- layer=1 filter=207 channel=26
    -26, -1, -14, -11, -23, -7, -6, -12, 3,
    -- layer=1 filter=207 channel=27
    -14, -7, 8, -1, -6, 10, 6, 8, 8,
    -- layer=1 filter=207 channel=28
    -19, -5, -4, -25, -3, -15, -10, -7, -20,
    -- layer=1 filter=207 channel=29
    1, 9, 3, 2, 3, -6, 14, 11, -5,
    -- layer=1 filter=207 channel=30
    -3, -1, -23, -11, -5, -17, -25, -15, 0,
    -- layer=1 filter=207 channel=31
    1, -8, -9, -15, -9, -7, -6, -19, -2,
    -- layer=1 filter=207 channel=32
    -3, 0, -10, -13, -3, -6, -9, -5, -6,
    -- layer=1 filter=207 channel=33
    9, 6, -4, 1, -3, 4, 7, -9, -5,
    -- layer=1 filter=207 channel=34
    8, 3, -10, 5, 0, 6, -2, -10, -13,
    -- layer=1 filter=207 channel=35
    5, -11, 8, -12, 5, 5, -3, -1, -3,
    -- layer=1 filter=207 channel=36
    3, 2, -9, 5, -1, 6, -8, 0, 5,
    -- layer=1 filter=207 channel=37
    -5, -8, 0, -22, -8, -13, -9, -9, -6,
    -- layer=1 filter=207 channel=38
    -16, -16, -26, -10, -11, -22, -7, -8, -5,
    -- layer=1 filter=207 channel=39
    -4, -9, -7, 5, 4, -6, 0, 6, 8,
    -- layer=1 filter=207 channel=40
    -8, -26, -29, -4, -14, -23, -28, -33, -22,
    -- layer=1 filter=207 channel=41
    -1, 1, -7, -6, -9, -10, -10, 0, 1,
    -- layer=1 filter=207 channel=42
    4, 0, -7, 3, -2, 2, -10, -11, -6,
    -- layer=1 filter=207 channel=43
    -4, -6, -1, -23, -11, -15, -23, -18, -9,
    -- layer=1 filter=207 channel=44
    -9, -12, -7, 3, 1, 1, -14, -3, -17,
    -- layer=1 filter=207 channel=45
    -10, -14, -11, -6, 0, -4, -19, -2, 0,
    -- layer=1 filter=207 channel=46
    4, -7, -8, -28, -22, -17, -16, 5, 5,
    -- layer=1 filter=207 channel=47
    -1, -10, -8, -11, -8, -9, -18, -11, -1,
    -- layer=1 filter=207 channel=48
    -15, -23, -20, -4, -4, -17, -20, -14, -2,
    -- layer=1 filter=207 channel=49
    0, -11, -16, -10, -6, 0, -1, 12, -7,
    -- layer=1 filter=207 channel=50
    5, 0, 6, 0, 6, 0, -1, -4, -5,
    -- layer=1 filter=207 channel=51
    -6, -4, 0, -15, 0, -18, -12, -20, -4,
    -- layer=1 filter=207 channel=52
    -10, 3, 0, 0, 4, -8, -5, 6, 0,
    -- layer=1 filter=207 channel=53
    0, 1, -3, 7, -5, -6, -2, -8, 1,
    -- layer=1 filter=207 channel=54
    -8, -17, -5, -11, -3, -15, -2, -4, -7,
    -- layer=1 filter=207 channel=55
    -9, -5, -11, -5, 0, 13, -9, -5, -1,
    -- layer=1 filter=207 channel=56
    2, -2, 7, 6, -10, 3, -9, -11, -5,
    -- layer=1 filter=207 channel=57
    -25, -15, -19, -24, -24, -27, -15, -11, -20,
    -- layer=1 filter=207 channel=58
    -4, -20, -9, 1, -11, -6, -4, -31, -17,
    -- layer=1 filter=207 channel=59
    -4, -5, 0, -11, 2, -9, 0, 4, 2,
    -- layer=1 filter=207 channel=60
    10, 5, -9, 0, 9, -7, -5, 9, -2,
    -- layer=1 filter=207 channel=61
    0, 5, 5, 7, 5, 5, 0, 3, -7,
    -- layer=1 filter=207 channel=62
    -18, -12, -6, -19, -19, -10, -15, -18, -4,
    -- layer=1 filter=207 channel=63
    -14, -13, -4, -11, 4, 1, -6, -11, 6,
    -- layer=1 filter=207 channel=64
    -3, 1, 4, -7, -10, -5, -1, 8, 6,
    -- layer=1 filter=207 channel=65
    -5, -19, -22, -5, -16, -18, -1, -8, -17,
    -- layer=1 filter=207 channel=66
    -8, 5, -1, -2, 6, 6, -7, 2, 0,
    -- layer=1 filter=207 channel=67
    -21, -4, -7, -10, -6, 1, -6, 13, -7,
    -- layer=1 filter=207 channel=68
    -12, 1, -7, -13, -19, -12, -4, 6, -4,
    -- layer=1 filter=207 channel=69
    -7, -17, -7, -10, -18, -6, -21, 5, -22,
    -- layer=1 filter=207 channel=70
    13, 11, 0, 16, 0, 1, 4, 14, -4,
    -- layer=1 filter=207 channel=71
    -14, -12, -8, -21, -10, -15, -22, -23, -15,
    -- layer=1 filter=207 channel=72
    -3, -1, -13, -4, 7, -12, -7, 6, -2,
    -- layer=1 filter=207 channel=73
    1, 5, -6, 1, 3, -5, -5, 5, 0,
    -- layer=1 filter=207 channel=74
    -9, -15, 0, -12, -7, -13, -7, 5, -11,
    -- layer=1 filter=207 channel=75
    7, -10, -5, -13, -11, -6, -20, -16, -17,
    -- layer=1 filter=207 channel=76
    1, 1, -18, -10, 2, -9, 1, -1, -11,
    -- layer=1 filter=207 channel=77
    -17, -4, -17, -20, -24, -19, -23, -5, -5,
    -- layer=1 filter=207 channel=78
    -2, -8, 3, -6, 4, 6, -7, -3, -2,
    -- layer=1 filter=207 channel=79
    -12, -13, -13, -13, -23, -7, -7, -9, -9,
    -- layer=1 filter=207 channel=80
    9, 7, 7, 0, 7, -4, 6, -8, 10,
    -- layer=1 filter=207 channel=81
    -22, -13, -18, -18, -3, -12, -23, -14, -17,
    -- layer=1 filter=207 channel=82
    -10, -26, -28, -22, -26, -23, -21, -11, -20,
    -- layer=1 filter=207 channel=83
    0, -1, -2, 0, -7, -15, -10, 1, -8,
    -- layer=1 filter=207 channel=84
    -15, -6, -19, -13, -12, -18, -24, -17, -6,
    -- layer=1 filter=207 channel=85
    -3, -20, -17, -5, -12, -16, -19, -17, -22,
    -- layer=1 filter=207 channel=86
    11, -7, 7, -2, 8, -5, 7, 4, 0,
    -- layer=1 filter=207 channel=87
    1, 0, 3, -12, 5, 5, -1, -11, 0,
    -- layer=1 filter=207 channel=88
    -6, -11, -8, -21, -18, -17, -23, -10, -22,
    -- layer=1 filter=207 channel=89
    -24, -24, -27, -7, -14, -8, -26, -1, -16,
    -- layer=1 filter=207 channel=90
    -20, -4, -11, -13, -9, -11, -9, -10, -15,
    -- layer=1 filter=207 channel=91
    1, -16, -22, 3, -18, -13, -3, -22, -6,
    -- layer=1 filter=207 channel=92
    -11, 5, 7, 0, -13, -10, 3, 1, -4,
    -- layer=1 filter=207 channel=93
    0, -16, -2, -17, -17, -3, -11, -5, -8,
    -- layer=1 filter=207 channel=94
    5, -10, -15, -10, 2, -14, 2, 3, -1,
    -- layer=1 filter=207 channel=95
    -4, -9, -13, -15, -9, -15, -23, -15, -4,
    -- layer=1 filter=207 channel=96
    -8, -10, -9, -1, -11, -2, -7, 8, -6,
    -- layer=1 filter=207 channel=97
    1, -9, -2, -1, 4, 0, 0, -11, -8,
    -- layer=1 filter=207 channel=98
    -16, -11, -9, -14, -5, -10, 2, -22, -9,
    -- layer=1 filter=207 channel=99
    -19, -4, -13, -17, -19, -8, -14, -16, -11,
    -- layer=1 filter=207 channel=100
    -8, -4, 1, 5, -14, 2, 2, 0, -5,
    -- layer=1 filter=207 channel=101
    -2, -24, -16, -23, -7, -15, -13, -9, -22,
    -- layer=1 filter=207 channel=102
    0, -7, -11, -15, 3, -14, 5, 1, -2,
    -- layer=1 filter=207 channel=103
    -5, -4, -1, -11, -12, -4, 9, -5, 11,
    -- layer=1 filter=207 channel=104
    -8, -3, -7, 8, 4, 2, 3, 3, -9,
    -- layer=1 filter=207 channel=105
    -3, -13, -5, 3, 2, -10, -3, -14, -2,
    -- layer=1 filter=207 channel=106
    -15, -2, -19, -5, -25, -18, -17, -20, -3,
    -- layer=1 filter=207 channel=107
    -8, 2, 6, 7, 0, 7, 0, 1, -5,
    -- layer=1 filter=207 channel=108
    -13, -8, -20, -14, -20, -25, -10, -17, -1,
    -- layer=1 filter=207 channel=109
    0, 0, -9, -7, 8, -7, 4, 1, -1,
    -- layer=1 filter=207 channel=110
    0, 6, -9, 7, 4, -1, 8, -3, -5,
    -- layer=1 filter=207 channel=111
    -1, -13, -25, -25, -3, -9, -20, -9, -10,
    -- layer=1 filter=207 channel=112
    -19, -8, -13, -9, -14, -15, -4, -11, -2,
    -- layer=1 filter=207 channel=113
    3, -20, -16, -4, -5, 3, 9, 11, 6,
    -- layer=1 filter=207 channel=114
    15, -9, 0, -9, -15, -16, -7, 1, -15,
    -- layer=1 filter=207 channel=115
    -10, -2, 2, -14, -5, 0, 3, -2, 6,
    -- layer=1 filter=207 channel=116
    0, -5, 2, -10, 10, 0, 0, 6, -6,
    -- layer=1 filter=207 channel=117
    1, -2, -10, -11, 0, 1, -21, -11, 11,
    -- layer=1 filter=207 channel=118
    -13, -16, -22, -4, -22, -15, -17, -16, -14,
    -- layer=1 filter=207 channel=119
    -9, -2, -14, -11, -5, -16, -16, -3, -13,
    -- layer=1 filter=207 channel=120
    -7, -26, -19, -9, -21, -16, -10, -6, -28,
    -- layer=1 filter=207 channel=121
    6, -12, -10, -15, 1, -17, -13, 6, -2,
    -- layer=1 filter=207 channel=122
    -1, -8, 7, -8, 3, 5, 0, 1, -4,
    -- layer=1 filter=207 channel=123
    -16, 2, -13, -8, 2, -12, 2, 0, -4,
    -- layer=1 filter=207 channel=124
    -9, -3, 2, -1, -3, 0, 4, 3, -10,
    -- layer=1 filter=207 channel=125
    0, 6, 9, 8, 8, 10, 3, 0, 6,
    -- layer=1 filter=207 channel=126
    -9, -17, -22, -14, -3, -4, -12, -11, -18,
    -- layer=1 filter=207 channel=127
    -5, -4, -24, -24, -16, -13, -27, -10, -16,
    -- layer=1 filter=208 channel=0
    2, 3, -7, -5, -3, 1, 8, -7, -3,
    -- layer=1 filter=208 channel=1
    3, -4, 2, 8, 0, -4, -9, 3, -2,
    -- layer=1 filter=208 channel=2
    -7, 5, 0, 1, 10, -5, -8, 0, 2,
    -- layer=1 filter=208 channel=3
    -1, 2, 0, 5, 0, -8, -11, 5, 1,
    -- layer=1 filter=208 channel=4
    -7, 4, 2, 6, -6, -12, 5, 2, 3,
    -- layer=1 filter=208 channel=5
    -4, -10, 1, 1, -3, 0, -5, 9, -9,
    -- layer=1 filter=208 channel=6
    7, 4, -1, -8, 5, 7, 3, -11, -2,
    -- layer=1 filter=208 channel=7
    9, 6, 0, 1, 7, 2, 5, -3, 0,
    -- layer=1 filter=208 channel=8
    3, 0, 2, -6, -4, 3, 8, 0, -3,
    -- layer=1 filter=208 channel=9
    6, 2, -11, 5, -4, 5, -7, 2, -4,
    -- layer=1 filter=208 channel=10
    7, 0, -3, 5, 2, -7, 7, -2, -1,
    -- layer=1 filter=208 channel=11
    -9, -1, -3, -3, -6, -1, 0, 6, -8,
    -- layer=1 filter=208 channel=12
    -5, -10, -10, 0, 3, -8, -6, -2, 6,
    -- layer=1 filter=208 channel=13
    5, 6, -2, -5, 1, -11, 3, 6, -8,
    -- layer=1 filter=208 channel=14
    -1, -1, -9, -1, 6, -5, -6, -5, -11,
    -- layer=1 filter=208 channel=15
    4, 0, 5, -2, 5, -1, 3, -7, 0,
    -- layer=1 filter=208 channel=16
    -8, -2, 4, -11, -6, -7, 4, -4, 7,
    -- layer=1 filter=208 channel=17
    3, 1, -6, -2, -7, 0, -4, -1, -4,
    -- layer=1 filter=208 channel=18
    0, 1, 4, -7, 5, 7, -2, -3, 7,
    -- layer=1 filter=208 channel=19
    -3, 8, 0, 9, 7, -8, 6, 8, -12,
    -- layer=1 filter=208 channel=20
    -7, 7, -11, 5, -5, -8, -2, -9, 4,
    -- layer=1 filter=208 channel=21
    5, 0, -2, -6, -9, -5, -8, -3, 2,
    -- layer=1 filter=208 channel=22
    -11, -5, -8, 7, 1, 4, -8, -7, 2,
    -- layer=1 filter=208 channel=23
    0, -5, -9, -4, -6, -2, -4, -1, 2,
    -- layer=1 filter=208 channel=24
    -9, -1, -7, 5, -6, -4, -2, -2, -12,
    -- layer=1 filter=208 channel=25
    2, 2, -6, 2, 0, -5, 11, -10, -4,
    -- layer=1 filter=208 channel=26
    1, 7, -7, 1, -12, -3, -4, -8, -2,
    -- layer=1 filter=208 channel=27
    0, -11, -9, -10, -3, 4, -1, -9, -2,
    -- layer=1 filter=208 channel=28
    -3, -7, 8, 1, 1, 2, -5, -12, -4,
    -- layer=1 filter=208 channel=29
    -10, 3, 2, -7, -10, -8, 8, 3, 9,
    -- layer=1 filter=208 channel=30
    -5, 0, -1, -3, 1, -11, -7, -6, 1,
    -- layer=1 filter=208 channel=31
    5, 1, 7, -4, 7, -6, -6, -5, -4,
    -- layer=1 filter=208 channel=32
    -12, -4, 0, 4, 5, -1, -11, -4, -5,
    -- layer=1 filter=208 channel=33
    8, 9, 4, 3, -6, 9, -2, 10, 1,
    -- layer=1 filter=208 channel=34
    -12, -12, -6, 7, 0, -3, -4, 1, 4,
    -- layer=1 filter=208 channel=35
    -12, -8, -4, -1, -9, -8, -11, -10, 4,
    -- layer=1 filter=208 channel=36
    0, -6, -5, 8, 0, 3, 7, -2, -6,
    -- layer=1 filter=208 channel=37
    7, -7, 1, -5, -3, 4, -10, -1, -8,
    -- layer=1 filter=208 channel=38
    -3, 7, -7, -3, -8, 1, -11, -10, 4,
    -- layer=1 filter=208 channel=39
    -8, 5, 1, -11, 8, 3, -10, -2, 3,
    -- layer=1 filter=208 channel=40
    1, -3, 2, -1, -3, 0, 1, -2, -4,
    -- layer=1 filter=208 channel=41
    -3, 0, 5, 6, 10, -6, -7, 5, -7,
    -- layer=1 filter=208 channel=42
    -4, 5, 6, 1, 11, 6, -5, 0, -9,
    -- layer=1 filter=208 channel=43
    -2, 6, -7, -5, 5, 6, 7, -9, -7,
    -- layer=1 filter=208 channel=44
    3, -8, 5, 0, 6, 1, 4, 10, -1,
    -- layer=1 filter=208 channel=45
    8, -4, 4, -10, 6, 0, 6, 5, 6,
    -- layer=1 filter=208 channel=46
    -11, -8, 4, -8, -5, -8, 1, -1, -5,
    -- layer=1 filter=208 channel=47
    -8, -9, -9, 5, 2, -7, 0, 7, -10,
    -- layer=1 filter=208 channel=48
    -9, -11, 2, 0, 6, -8, -2, -9, -8,
    -- layer=1 filter=208 channel=49
    0, -6, -7, -3, -4, -3, -7, -1, -3,
    -- layer=1 filter=208 channel=50
    -1, -10, -4, -7, -11, 5, 4, 2, -9,
    -- layer=1 filter=208 channel=51
    2, -8, -11, -8, -7, 4, -4, -8, -1,
    -- layer=1 filter=208 channel=52
    5, 8, 3, 0, 7, 0, -9, 3, -9,
    -- layer=1 filter=208 channel=53
    -9, 1, -3, -1, 8, 5, 4, 0, -2,
    -- layer=1 filter=208 channel=54
    -5, 0, -8, 5, -10, 3, 2, -11, 5,
    -- layer=1 filter=208 channel=55
    7, 5, -5, -3, -1, 9, 2, 3, -3,
    -- layer=1 filter=208 channel=56
    -3, 2, 6, 1, 6, -5, -8, 6, 1,
    -- layer=1 filter=208 channel=57
    7, 0, 5, 0, -3, 7, -8, 3, 8,
    -- layer=1 filter=208 channel=58
    0, -4, 1, -2, -7, 4, 8, -9, -11,
    -- layer=1 filter=208 channel=59
    -8, 0, -9, 0, -1, 1, 6, 7, -1,
    -- layer=1 filter=208 channel=60
    8, 1, 11, -2, -9, 6, -2, 10, -4,
    -- layer=1 filter=208 channel=61
    -8, -4, -6, 1, 4, -9, -1, -6, 0,
    -- layer=1 filter=208 channel=62
    -3, -8, -6, -16, -11, 0, 6, -11, 6,
    -- layer=1 filter=208 channel=63
    0, 0, 5, -2, 5, 0, -4, 7, -8,
    -- layer=1 filter=208 channel=64
    -8, -3, 8, -4, 5, -1, 0, -1, -7,
    -- layer=1 filter=208 channel=65
    5, 2, -7, 8, -4, 3, 2, 7, -7,
    -- layer=1 filter=208 channel=66
    -8, -6, 6, -6, 0, -1, -9, 6, -4,
    -- layer=1 filter=208 channel=67
    8, 9, -6, 2, 0, -7, 5, -9, -8,
    -- layer=1 filter=208 channel=68
    2, -5, -4, 6, 1, 1, -11, -10, 7,
    -- layer=1 filter=208 channel=69
    0, 8, 0, 0, -7, -5, -3, 7, 1,
    -- layer=1 filter=208 channel=70
    2, -5, 9, 5, -7, 2, -8, 5, 9,
    -- layer=1 filter=208 channel=71
    -14, -6, 0, -2, -6, -8, 0, 6, -13,
    -- layer=1 filter=208 channel=72
    8, 7, 6, -2, -4, 5, 0, -10, 2,
    -- layer=1 filter=208 channel=73
    -2, 0, 6, 5, 0, 0, 1, 0, -7,
    -- layer=1 filter=208 channel=74
    0, 9, -6, 3, 5, -9, -8, -9, 8,
    -- layer=1 filter=208 channel=75
    -16, -7, -6, -3, -4, -4, 8, 0, -4,
    -- layer=1 filter=208 channel=76
    7, -1, -3, -6, 2, 4, -3, 7, 0,
    -- layer=1 filter=208 channel=77
    -5, 5, -3, -11, -6, -6, 2, -3, -6,
    -- layer=1 filter=208 channel=78
    0, -2, -2, -10, 2, 2, 5, -1, -10,
    -- layer=1 filter=208 channel=79
    -4, -1, 4, -10, -14, 3, 5, 1, -5,
    -- layer=1 filter=208 channel=80
    2, -2, -5, -8, -9, 8, -6, -4, 0,
    -- layer=1 filter=208 channel=81
    6, -12, 0, -11, 6, -9, -5, -3, 5,
    -- layer=1 filter=208 channel=82
    -5, -2, 1, 0, -2, -10, 2, -3, -4,
    -- layer=1 filter=208 channel=83
    0, -4, -1, -10, -6, 3, 0, 6, -9,
    -- layer=1 filter=208 channel=84
    6, 4, -4, -5, -6, -8, -1, -9, 0,
    -- layer=1 filter=208 channel=85
    -10, -10, -12, -5, 0, -6, 6, -10, 6,
    -- layer=1 filter=208 channel=86
    6, -10, -6, 8, -5, -2, 6, 2, 1,
    -- layer=1 filter=208 channel=87
    0, -1, 6, 9, -5, 6, -2, 3, 7,
    -- layer=1 filter=208 channel=88
    6, -9, -1, 3, 2, 9, 2, 6, -3,
    -- layer=1 filter=208 channel=89
    -7, -12, 1, 2, 5, 2, -10, -12, 0,
    -- layer=1 filter=208 channel=90
    -7, -3, -4, -11, -2, 0, 0, -6, -8,
    -- layer=1 filter=208 channel=91
    -9, -8, 2, 0, -8, -2, -4, 3, -5,
    -- layer=1 filter=208 channel=92
    -11, 8, 7, -7, 5, -11, 4, -7, -7,
    -- layer=1 filter=208 channel=93
    -5, -4, -2, -1, 5, -1, -2, 4, -2,
    -- layer=1 filter=208 channel=94
    -8, 5, 5, 0, -6, 4, -5, 0, 6,
    -- layer=1 filter=208 channel=95
    -13, -2, 1, -4, -7, -12, -9, -9, -6,
    -- layer=1 filter=208 channel=96
    -4, -7, 1, -7, -5, 4, 5, 0, -1,
    -- layer=1 filter=208 channel=97
    6, -8, -8, -7, 2, -2, -5, -3, 3,
    -- layer=1 filter=208 channel=98
    5, -8, 6, -4, -12, -7, -7, -4, 7,
    -- layer=1 filter=208 channel=99
    6, -6, 0, -9, 7, -1, -9, 0, 0,
    -- layer=1 filter=208 channel=100
    -10, -1, -1, -8, 5, 4, 5, 6, 8,
    -- layer=1 filter=208 channel=101
    -3, 0, -5, 5, -11, 5, 1, -8, 2,
    -- layer=1 filter=208 channel=102
    -1, 3, -4, 2, -7, 5, -5, 2, -4,
    -- layer=1 filter=208 channel=103
    -3, 2, 6, 5, 10, -3, 0, 2, -2,
    -- layer=1 filter=208 channel=104
    0, -3, 9, 8, -7, -7, 6, -2, -7,
    -- layer=1 filter=208 channel=105
    -8, -6, 1, 3, -2, -11, 5, 0, 7,
    -- layer=1 filter=208 channel=106
    -8, -9, -2, -5, 5, -6, -9, 0, 7,
    -- layer=1 filter=208 channel=107
    -1, 9, 5, 9, 3, -8, 0, 6, 8,
    -- layer=1 filter=208 channel=108
    -10, -1, 0, 3, -1, -10, -7, -10, -14,
    -- layer=1 filter=208 channel=109
    3, 2, 0, -9, -7, -9, 2, -4, -3,
    -- layer=1 filter=208 channel=110
    0, -1, 1, -1, -5, 3, -6, 0, -7,
    -- layer=1 filter=208 channel=111
    2, -11, -3, -3, 0, 1, -4, 5, -1,
    -- layer=1 filter=208 channel=112
    -10, 2, 0, -1, -3, -11, -2, -3, -7,
    -- layer=1 filter=208 channel=113
    -12, 2, -11, 0, 0, 1, 2, -11, -8,
    -- layer=1 filter=208 channel=114
    -6, -1, -3, 3, -8, 4, -8, 6, 2,
    -- layer=1 filter=208 channel=115
    -3, -10, -9, -3, 0, 3, -9, 8, -6,
    -- layer=1 filter=208 channel=116
    9, 9, 5, -5, -3, 6, -10, 0, 2,
    -- layer=1 filter=208 channel=117
    0, 2, -5, 10, -2, 4, -5, -2, -6,
    -- layer=1 filter=208 channel=118
    0, -13, -5, 6, -8, 8, -10, 0, 6,
    -- layer=1 filter=208 channel=119
    -2, -6, 3, -15, -6, 1, -4, -2, -6,
    -- layer=1 filter=208 channel=120
    -3, 7, -2, -6, -4, -8, -2, 3, -2,
    -- layer=1 filter=208 channel=121
    -6, 4, 5, -4, -9, -4, -7, 0, 2,
    -- layer=1 filter=208 channel=122
    3, -1, -3, 3, -5, -5, 0, 2, 6,
    -- layer=1 filter=208 channel=123
    -8, -10, -4, -9, 6, -6, 1, -5, 3,
    -- layer=1 filter=208 channel=124
    2, -5, -6, 8, 0, -6, -1, -5, -7,
    -- layer=1 filter=208 channel=125
    1, 7, -1, -6, 1, 0, -3, 8, 8,
    -- layer=1 filter=208 channel=126
    -5, 4, -9, -9, 1, 2, 4, -5, -8,
    -- layer=1 filter=208 channel=127
    -1, 0, 2, 2, 3, -11, 1, -11, -9,
    -- layer=1 filter=209 channel=0
    -9, 1, -5, -12, -2, -7, -6, -5, -11,
    -- layer=1 filter=209 channel=1
    -20, -15, -49, -12, -18, -6, -44, -43, 41,
    -- layer=1 filter=209 channel=2
    39, 32, 50, 38, 27, 38, 34, 29, 28,
    -- layer=1 filter=209 channel=3
    -7, -11, 4, 9, -8, 0, 9, 2, 6,
    -- layer=1 filter=209 channel=4
    15, 4, 7, -5, 3, -15, -3, -8, -10,
    -- layer=1 filter=209 channel=5
    -6, -12, -17, -42, -26, 13, -30, -10, 36,
    -- layer=1 filter=209 channel=6
    13, -18, -17, 12, 0, -9, 12, 2, -33,
    -- layer=1 filter=209 channel=7
    -41, -51, -124, -36, -52, -31, -84, 36, -17,
    -- layer=1 filter=209 channel=8
    -16, -38, -55, -39, -39, 6, -76, -19, 23,
    -- layer=1 filter=209 channel=9
    41, 40, 68, 54, 43, 50, 57, 60, 61,
    -- layer=1 filter=209 channel=10
    -36, -70, -101, -33, -32, -6, -58, 46, -6,
    -- layer=1 filter=209 channel=11
    -28, -37, -27, -21, -20, -27, -28, -42, -40,
    -- layer=1 filter=209 channel=12
    40, 40, 0, 68, 38, 33, 75, 56, 51,
    -- layer=1 filter=209 channel=13
    -5, -8, 2, -22, -12, -16, -13, -27, 7,
    -- layer=1 filter=209 channel=14
    1, -1, -68, 5, -11, -5, 14, 3, 6,
    -- layer=1 filter=209 channel=15
    46, 47, 52, 15, 29, 51, 32, -3, 53,
    -- layer=1 filter=209 channel=16
    1, -21, -32, -37, -2, 42, -64, 6, 18,
    -- layer=1 filter=209 channel=17
    -11, -18, -25, -18, -18, -31, -11, -39, -1,
    -- layer=1 filter=209 channel=18
    -8, -28, -41, 6, 9, -9, -4, -42, -19,
    -- layer=1 filter=209 channel=19
    38, -11, 26, 1, 0, 26, -31, 47, -14,
    -- layer=1 filter=209 channel=20
    -19, -11, -24, -15, -26, -19, -53, -29, 8,
    -- layer=1 filter=209 channel=21
    -9, -14, -4, -9, -15, -8, 0, -5, -5,
    -- layer=1 filter=209 channel=22
    -9, -15, -26, -16, -13, -5, -40, -21, 1,
    -- layer=1 filter=209 channel=23
    -37, -35, -84, -43, -37, -39, -20, -6, -24,
    -- layer=1 filter=209 channel=24
    -11, 0, 8, -4, -4, 0, -2, 5, -4,
    -- layer=1 filter=209 channel=25
    1, -39, -61, -16, -28, 0, -65, 26, -11,
    -- layer=1 filter=209 channel=26
    5, -16, 6, -9, -12, -4, -16, -27, 34,
    -- layer=1 filter=209 channel=27
    8, 32, 37, 27, 32, 42, 29, 15, 38,
    -- layer=1 filter=209 channel=28
    -27, -56, -104, -38, -50, -1, -93, 23, -3,
    -- layer=1 filter=209 channel=29
    -55, -44, -35, -53, -43, -49, -38, -62, -47,
    -- layer=1 filter=209 channel=30
    17, -22, -38, -4, -15, -12, -29, -55, -29,
    -- layer=1 filter=209 channel=31
    16, 22, 0, 33, 25, 5, 35, 5, 20,
    -- layer=1 filter=209 channel=32
    3, -22, 1, -24, -20, 6, -34, -51, 16,
    -- layer=1 filter=209 channel=33
    -17, -24, -22, 0, -8, -27, -12, -21, -20,
    -- layer=1 filter=209 channel=34
    0, -9, -33, 12, -16, -31, -8, -23, -41,
    -- layer=1 filter=209 channel=35
    6, 14, 3, 5, 2, -7, -1, -12, 7,
    -- layer=1 filter=209 channel=36
    -35, -57, -50, -28, -22, -22, -28, -41, -31,
    -- layer=1 filter=209 channel=37
    24, -6, 5, -21, 1, 26, -39, 33, 9,
    -- layer=1 filter=209 channel=38
    4, -12, -1, -8, -7, -11, -15, 2, -2,
    -- layer=1 filter=209 channel=39
    -17, 2, -10, -5, -21, -13, -18, -3, 8,
    -- layer=1 filter=209 channel=40
    1, 0, -20, 29, 0, -6, 25, 2, -13,
    -- layer=1 filter=209 channel=41
    7, 3, 34, 7, 3, 20, 34, 9, 31,
    -- layer=1 filter=209 channel=42
    31, 26, 47, 30, 35, 42, 36, 29, 35,
    -- layer=1 filter=209 channel=43
    -9, -47, -72, -53, -23, 2, -80, 11, 14,
    -- layer=1 filter=209 channel=44
    -32, -45, -30, -60, -49, -18, -41, -94, 14,
    -- layer=1 filter=209 channel=45
    -12, 9, -20, -20, -12, -1, -17, -42, 18,
    -- layer=1 filter=209 channel=46
    41, 28, 58, 31, 5, 24, 11, 34, 29,
    -- layer=1 filter=209 channel=47
    11, 21, 8, 3, 17, 31, 18, 34, 10,
    -- layer=1 filter=209 channel=48
    -22, -29, -30, -19, -20, -23, -15, 4, -28,
    -- layer=1 filter=209 channel=49
    18, 18, 22, 20, 24, 16, 30, 20, 29,
    -- layer=1 filter=209 channel=50
    -3, 8, -16, -16, -30, 5, -19, -24, -20,
    -- layer=1 filter=209 channel=51
    -11, -26, -40, 0, -1, -17, -16, 24, 3,
    -- layer=1 filter=209 channel=52
    -7, -20, 4, 6, -4, 0, -22, -34, 1,
    -- layer=1 filter=209 channel=53
    -15, 3, 2, 4, 8, -3, 1, 20, 9,
    -- layer=1 filter=209 channel=54
    2, -15, -3, 11, 5, 21, -16, 50, -1,
    -- layer=1 filter=209 channel=55
    -13, -10, 10, -11, -2, 2, 7, -3, -3,
    -- layer=1 filter=209 channel=56
    4, -8, 9, -5, 7, 1, 2, 8, 4,
    -- layer=1 filter=209 channel=57
    -19, -19, -38, -9, 1, 10, -10, 47, -8,
    -- layer=1 filter=209 channel=58
    -28, -29, -78, -23, -31, -10, -25, 42, -56,
    -- layer=1 filter=209 channel=59
    -3, -8, 1, 0, -5, 0, -5, -12, 0,
    -- layer=1 filter=209 channel=60
    7, -7, 9, -6, 14, 21, 0, -4, 4,
    -- layer=1 filter=209 channel=61
    -4, 6, -11, 12, 6, -9, 0, 9, -3,
    -- layer=1 filter=209 channel=62
    -22, -67, -65, -60, -32, 23, -81, 16, 19,
    -- layer=1 filter=209 channel=63
    -34, -47, -37, -30, -36, -21, -40, -59, -34,
    -- layer=1 filter=209 channel=64
    -12, -12, -9, 0, -9, -13, -15, -7, -3,
    -- layer=1 filter=209 channel=65
    -16, -8, -7, 6, 7, 1, -1, -3, -3,
    -- layer=1 filter=209 channel=66
    -19, -7, -18, -19, -22, -19, -19, -6, 1,
    -- layer=1 filter=209 channel=67
    -10, 0, -16, 28, -10, -4, 8, 39, 20,
    -- layer=1 filter=209 channel=68
    -27, -54, -23, -43, -49, -18, -38, -75, 8,
    -- layer=1 filter=209 channel=69
    18, 3, 22, -14, 12, 20, -26, -9, 28,
    -- layer=1 filter=209 channel=70
    -42, -30, -27, 21, 8, -30, 38, 10, -15,
    -- layer=1 filter=209 channel=71
    -14, -10, -25, -19, -23, -15, -19, -6, -21,
    -- layer=1 filter=209 channel=72
    39, -5, 20, 2, -10, 7, -19, 32, -3,
    -- layer=1 filter=209 channel=73
    5, -4, -10, 5, -12, -9, -1, 2, -4,
    -- layer=1 filter=209 channel=74
    5, -32, -18, -40, -5, -31, 5, -9, -5,
    -- layer=1 filter=209 channel=75
    2, 5, -32, 18, 1, 2, 40, 10, 17,
    -- layer=1 filter=209 channel=76
    13, -15, -21, -20, -3, 5, -16, -7, -11,
    -- layer=1 filter=209 channel=77
    -17, -23, -14, -29, -9, -19, -42, -19, -14,
    -- layer=1 filter=209 channel=78
    -13, -24, -19, -22, -9, -13, -37, 22, -13,
    -- layer=1 filter=209 channel=79
    -11, -21, -28, -36, -19, 22, -62, 9, 11,
    -- layer=1 filter=209 channel=80
    28, 5, 11, 2, 5, 37, 18, 12, 23,
    -- layer=1 filter=209 channel=81
    -15, -13, -15, -25, -21, -15, -20, -5, -25,
    -- layer=1 filter=209 channel=82
    -13, -14, -25, -16, -17, -15, -21, -18, -10,
    -- layer=1 filter=209 channel=83
    -18, -23, -35, -46, 0, -27, -31, -58, 11,
    -- layer=1 filter=209 channel=84
    -2, -46, -45, -15, -13, -3, -24, -50, 5,
    -- layer=1 filter=209 channel=85
    -1, 20, -28, -5, -13, 32, -10, 48, -13,
    -- layer=1 filter=209 channel=86
    -29, -15, -22, -25, -37, -15, -19, -25, 6,
    -- layer=1 filter=209 channel=87
    59, 19, 75, 33, 29, 40, 31, 65, 33,
    -- layer=1 filter=209 channel=88
    23, 9, 31, 33, 25, 26, 24, 23, 20,
    -- layer=1 filter=209 channel=89
    -20, -15, -16, -13, -12, -15, -14, -13, -14,
    -- layer=1 filter=209 channel=90
    -31, -33, -29, -63, -60, -36, -43, -90, 16,
    -- layer=1 filter=209 channel=91
    -4, -12, -42, 8, -4, -16, -13, -6, -21,
    -- layer=1 filter=209 channel=92
    31, 44, 76, 23, 46, 71, 45, 25, 69,
    -- layer=1 filter=209 channel=93
    -26, -27, -27, -23, -25, -23, -23, -15, -9,
    -- layer=1 filter=209 channel=94
    3, -18, -13, -4, -18, -13, -15, -11, -3,
    -- layer=1 filter=209 channel=95
    -1, -47, -54, -27, -17, -11, -16, -41, -3,
    -- layer=1 filter=209 channel=96
    15, 30, 43, 35, 37, 54, 52, 50, 36,
    -- layer=1 filter=209 channel=97
    -24, -16, -5, -12, -12, -25, -14, -13, 15,
    -- layer=1 filter=209 channel=98
    -4, -35, -41, -24, -1, 16, -76, 27, 18,
    -- layer=1 filter=209 channel=99
    -29, -31, -30, -43, -6, -8, -52, 52, 17,
    -- layer=1 filter=209 channel=100
    -18, -42, -31, -27, -10, -4, -18, -54, -18,
    -- layer=1 filter=209 channel=101
    -23, -29, -38, -23, -10, -28, -23, -24, -20,
    -- layer=1 filter=209 channel=102
    0, -19, -19, -24, -3, -19, -18, -28, -21,
    -- layer=1 filter=209 channel=103
    -17, -10, -12, 9, 0, 9, 0, -4, -28,
    -- layer=1 filter=209 channel=104
    14, 29, -13, -6, 3, -17, 5, 23, -2,
    -- layer=1 filter=209 channel=105
    -20, -16, -19, -16, -20, -14, -19, 6, 10,
    -- layer=1 filter=209 channel=106
    -2, -2, -9, -3, -15, -17, -3, -34, 10,
    -- layer=1 filter=209 channel=107
    -13, -6, -7, -1, 2, -15, -9, -11, -2,
    -- layer=1 filter=209 channel=108
    0, -13, -16, -37, -28, -7, -18, -45, 14,
    -- layer=1 filter=209 channel=109
    -1, -4, -5, -5, -7, -7, -4, -6, 0,
    -- layer=1 filter=209 channel=110
    4, -13, -4, 0, -8, 3, -6, -15, 4,
    -- layer=1 filter=209 channel=111
    -8, -34, -43, 0, -17, -14, -9, -40, -5,
    -- layer=1 filter=209 channel=112
    -55, -67, -91, -17, -4, -12, -43, -46, -23,
    -- layer=1 filter=209 channel=113
    35, 22, 24, 38, 25, 36, 28, 40, 29,
    -- layer=1 filter=209 channel=114
    -4, -4, 0, -16, -3, 30, -35, -14, 19,
    -- layer=1 filter=209 channel=115
    -21, -34, -56, -12, -23, -1, -50, 15, 9,
    -- layer=1 filter=209 channel=116
    -8, -9, -8, -5, 2, 5, -2, -4, -3,
    -- layer=1 filter=209 channel=117
    -64, -55, -111, 2, -22, -39, -29, -35, -52,
    -- layer=1 filter=209 channel=118
    6, -34, -17, 0, -4, -7, -31, -38, -18,
    -- layer=1 filter=209 channel=119
    -4, -41, -23, -36, -30, -15, -29, -69, 4,
    -- layer=1 filter=209 channel=120
    -15, -6, -20, -11, -5, 5, -31, 20, -5,
    -- layer=1 filter=209 channel=121
    15, -6, 1, 8, 9, -16, 6, -11, -4,
    -- layer=1 filter=209 channel=122
    9, 8, 3, 5, -6, -9, 3, -9, 4,
    -- layer=1 filter=209 channel=123
    -18, 0, -16, -9, -12, -23, -3, 0, -9,
    -- layer=1 filter=209 channel=124
    19, 3, 14, 18, 19, 4, 25, 27, 23,
    -- layer=1 filter=209 channel=125
    -6, -14, -7, 28, 17, 2, 33, 26, 0,
    -- layer=1 filter=209 channel=126
    -20, -8, -45, -30, -2, 3, -68, -22, 22,
    -- layer=1 filter=209 channel=127
    -1, -30, -35, -2, -7, -8, -31, -37, -22,
    -- layer=1 filter=210 channel=0
    -12, -9, -9, -15, -2, -11, -13, -10, -8,
    -- layer=1 filter=210 channel=1
    1, -1, 0, 5, -5, -7, 3, -8, -4,
    -- layer=1 filter=210 channel=2
    7, -8, -2, -4, -5, -1, -7, 0, -8,
    -- layer=1 filter=210 channel=3
    1, 1, 4, -2, -7, 0, 0, 6, -3,
    -- layer=1 filter=210 channel=4
    7, -6, -9, 0, -1, 1, -6, 4, -7,
    -- layer=1 filter=210 channel=5
    -2, -8, -10, -4, -6, -7, -7, -5, 0,
    -- layer=1 filter=210 channel=6
    0, -5, -10, 4, -5, -2, 1, 4, 0,
    -- layer=1 filter=210 channel=7
    2, -6, 10, -14, -8, 2, -16, 4, 13,
    -- layer=1 filter=210 channel=8
    2, -6, -5, -2, 5, -16, -1, -10, 2,
    -- layer=1 filter=210 channel=9
    -4, 9, -8, -2, 2, -4, -3, 6, -9,
    -- layer=1 filter=210 channel=10
    -9, -4, -7, -9, 0, -3, 0, -7, 10,
    -- layer=1 filter=210 channel=11
    4, -4, -4, -5, -11, 4, 9, 0, 7,
    -- layer=1 filter=210 channel=12
    2, 1, 0, -4, 0, -4, -4, 6, -6,
    -- layer=1 filter=210 channel=13
    -9, -1, -4, -6, -7, 3, -9, 11, -6,
    -- layer=1 filter=210 channel=14
    -7, 3, -5, -8, -11, 2, 0, 4, 5,
    -- layer=1 filter=210 channel=15
    0, 5, 8, 4, -6, -7, 5, -7, -8,
    -- layer=1 filter=210 channel=16
    -13, 8, -7, -11, -2, -17, -6, -3, -4,
    -- layer=1 filter=210 channel=17
    8, 8, -8, 7, -2, -2, -10, 4, 8,
    -- layer=1 filter=210 channel=18
    -14, 3, -6, -11, -16, -9, -11, -9, -5,
    -- layer=1 filter=210 channel=19
    4, 7, 1, 4, 2, -5, 6, 6, 0,
    -- layer=1 filter=210 channel=20
    -1, -13, -1, 3, -3, 5, -11, 0, -12,
    -- layer=1 filter=210 channel=21
    1, 4, -3, -2, 1, 7, -15, -15, -10,
    -- layer=1 filter=210 channel=22
    2, 0, -4, -5, 3, 4, -2, 4, -4,
    -- layer=1 filter=210 channel=23
    3, -4, -1, 3, -7, -2, -8, -10, -8,
    -- layer=1 filter=210 channel=24
    6, 0, 6, 3, 3, -5, 0, -7, -7,
    -- layer=1 filter=210 channel=25
    1, 2, -7, -11, 2, -10, 5, -12, 0,
    -- layer=1 filter=210 channel=26
    0, -15, -4, -5, -16, -7, 0, 0, 3,
    -- layer=1 filter=210 channel=27
    1, 6, -11, 5, -2, -13, -5, -15, -9,
    -- layer=1 filter=210 channel=28
    -2, 5, 4, 0, -5, -3, -12, -5, 10,
    -- layer=1 filter=210 channel=29
    -10, -2, -4, -9, -5, -9, -10, 4, -5,
    -- layer=1 filter=210 channel=30
    5, 0, 1, -14, -15, 6, 13, 8, -11,
    -- layer=1 filter=210 channel=31
    -13, -4, -11, -1, -5, 4, -7, 3, 4,
    -- layer=1 filter=210 channel=32
    3, -4, -7, 3, -11, -4, -3, -3, -10,
    -- layer=1 filter=210 channel=33
    -7, 5, -3, 2, 8, 9, -3, 7, 5,
    -- layer=1 filter=210 channel=34
    -5, 0, 2, -6, -4, -7, 1, -4, 4,
    -- layer=1 filter=210 channel=35
    -8, -11, 7, 0, 1, -10, -10, -7, 0,
    -- layer=1 filter=210 channel=36
    -5, -5, 4, 3, 0, -13, 7, -9, 3,
    -- layer=1 filter=210 channel=37
    -12, -9, -18, -15, -13, -3, -5, 1, 11,
    -- layer=1 filter=210 channel=38
    6, -2, 7, -6, 5, 3, -5, 9, -4,
    -- layer=1 filter=210 channel=39
    -9, -1, -6, -3, 4, -9, -4, -3, 0,
    -- layer=1 filter=210 channel=40
    0, -1, -4, 5, -10, -3, 2, 0, 5,
    -- layer=1 filter=210 channel=41
    -1, 2, -6, 8, 0, 6, 0, 5, -5,
    -- layer=1 filter=210 channel=42
    -6, -5, -2, 6, 4, 1, -9, -4, 0,
    -- layer=1 filter=210 channel=43
    -5, -10, 5, 8, -5, 0, 6, -14, 2,
    -- layer=1 filter=210 channel=44
    -8, -15, 1, -5, 3, 0, 4, -1, 2,
    -- layer=1 filter=210 channel=45
    -11, 3, 1, 0, -6, 3, 0, 3, 4,
    -- layer=1 filter=210 channel=46
    8, -10, -10, -2, -10, 2, 4, 3, -3,
    -- layer=1 filter=210 channel=47
    6, 4, 2, 4, 1, 7, 0, 7, 5,
    -- layer=1 filter=210 channel=48
    -13, 2, -12, -8, 2, 0, 4, -4, -13,
    -- layer=1 filter=210 channel=49
    5, -7, 4, -2, 0, 3, -9, -7, 1,
    -- layer=1 filter=210 channel=50
    3, 5, -9, 0, 0, -7, -2, 9, 9,
    -- layer=1 filter=210 channel=51
    -2, -5, 7, -2, 5, -8, -7, -12, -7,
    -- layer=1 filter=210 channel=52
    -7, -6, -5, -9, 0, -5, 3, 7, 1,
    -- layer=1 filter=210 channel=53
    -5, 3, 5, -1, 5, -3, -5, -10, 2,
    -- layer=1 filter=210 channel=54
    -16, 2, -12, 1, -20, -4, 0, -3, 0,
    -- layer=1 filter=210 channel=55
    -9, 2, 3, -5, -3, -10, 4, -13, 5,
    -- layer=1 filter=210 channel=56
    6, 2, -4, 8, -4, 8, 5, -1, -8,
    -- layer=1 filter=210 channel=57
    -1, -2, -9, -10, -2, 1, 7, -6, 8,
    -- layer=1 filter=210 channel=58
    5, -16, 0, 0, 0, -5, -7, 4, 18,
    -- layer=1 filter=210 channel=59
    5, -3, -11, -6, -10, -3, 2, -11, 4,
    -- layer=1 filter=210 channel=60
    6, -9, 8, 3, 0, 9, -11, -10, 5,
    -- layer=1 filter=210 channel=61
    2, 12, 7, 0, 11, -2, 2, 3, -11,
    -- layer=1 filter=210 channel=62
    -3, 1, -5, -1, -21, -16, -3, -9, 6,
    -- layer=1 filter=210 channel=63
    0, -8, -7, -16, -4, -6, -1, -4, -17,
    -- layer=1 filter=210 channel=64
    1, -6, 4, -2, -3, -6, 4, -9, -8,
    -- layer=1 filter=210 channel=65
    -8, -13, -10, -8, -6, -4, 2, -9, -15,
    -- layer=1 filter=210 channel=66
    -2, -9, -1, 0, 0, -18, -1, 1, -7,
    -- layer=1 filter=210 channel=67
    12, 15, 5, 0, 16, 7, 0, -3, -8,
    -- layer=1 filter=210 channel=68
    4, -3, -2, -3, -14, -7, -3, 4, 3,
    -- layer=1 filter=210 channel=69
    -5, -1, 12, 4, -5, -19, -7, -4, 2,
    -- layer=1 filter=210 channel=70
    3, -10, 1, -8, -8, 6, 12, 0, -8,
    -- layer=1 filter=210 channel=71
    1, -14, -5, -11, -2, 1, -15, -2, -14,
    -- layer=1 filter=210 channel=72
    -5, -5, 0, -10, -11, -12, 5, 6, -14,
    -- layer=1 filter=210 channel=73
    4, -8, 0, 5, -1, -9, -6, 5, 3,
    -- layer=1 filter=210 channel=74
    -3, -10, 2, 3, 6, 7, 10, -8, -8,
    -- layer=1 filter=210 channel=75
    -12, -8, 1, -11, -11, 14, -7, 0, -2,
    -- layer=1 filter=210 channel=76
    -5, -8, -4, -3, -5, -14, 1, -8, -7,
    -- layer=1 filter=210 channel=77
    -10, 6, 0, -8, -8, -1, -7, -9, -6,
    -- layer=1 filter=210 channel=78
    0, -9, -4, 5, -5, -4, -8, 8, -4,
    -- layer=1 filter=210 channel=79
    -6, -7, 3, 9, -5, -19, -9, -1, -4,
    -- layer=1 filter=210 channel=80
    -4, -2, -8, 2, 6, -1, 2, -7, -6,
    -- layer=1 filter=210 channel=81
    -1, 4, 0, -7, -13, 2, -17, 1, -6,
    -- layer=1 filter=210 channel=82
    3, 6, -5, 6, -7, 5, -8, -3, -3,
    -- layer=1 filter=210 channel=83
    -3, -5, -11, -4, 5, 4, -11, -8, 7,
    -- layer=1 filter=210 channel=84
    -9, -5, -11, -5, -12, 7, 4, -2, 2,
    -- layer=1 filter=210 channel=85
    7, -8, 7, -8, -15, 9, -14, -5, 5,
    -- layer=1 filter=210 channel=86
    -3, -13, -7, -11, -10, -3, 3, 7, 0,
    -- layer=1 filter=210 channel=87
    -3, 4, 6, 0, 7, 7, -4, -4, -7,
    -- layer=1 filter=210 channel=88
    -9, -7, 8, -7, -5, -6, -2, 3, -6,
    -- layer=1 filter=210 channel=89
    -9, 6, 1, -8, -3, 1, -2, -13, -10,
    -- layer=1 filter=210 channel=90
    -12, -10, -6, -8, 4, -10, 6, -4, -9,
    -- layer=1 filter=210 channel=91
    1, 8, -2, 2, -7, 0, 6, -1, 4,
    -- layer=1 filter=210 channel=92
    0, 9, -8, 4, 2, -1, -7, 5, -10,
    -- layer=1 filter=210 channel=93
    3, 4, 0, -13, -11, -5, -2, -4, -14,
    -- layer=1 filter=210 channel=94
    -9, -13, 0, -8, -7, -16, -6, -11, -8,
    -- layer=1 filter=210 channel=95
    -7, -16, -4, -2, -5, -10, 0, -13, -2,
    -- layer=1 filter=210 channel=96
    -8, -11, 0, 0, -3, 0, 0, 6, -9,
    -- layer=1 filter=210 channel=97
    -8, 3, 0, -7, -8, -17, -11, -7, -17,
    -- layer=1 filter=210 channel=98
    -2, 0, 2, -8, 0, -10, -1, 7, 6,
    -- layer=1 filter=210 channel=99
    7, 0, -9, -13, -1, -12, -10, 0, 4,
    -- layer=1 filter=210 channel=100
    2, 0, -3, -5, 1, -9, 8, -11, -4,
    -- layer=1 filter=210 channel=101
    1, 2, -8, -1, 0, 7, -13, -12, -10,
    -- layer=1 filter=210 channel=102
    -5, 1, -8, 5, 3, -4, 4, -8, -2,
    -- layer=1 filter=210 channel=103
    -13, -8, -12, -8, -11, -10, -12, 0, -1,
    -- layer=1 filter=210 channel=104
    -7, -7, -4, -8, 8, 9, 8, -9, -2,
    -- layer=1 filter=210 channel=105
    -8, -6, 3, -11, -5, -8, -15, -9, 0,
    -- layer=1 filter=210 channel=106
    -6, 3, 2, 5, -2, 8, 9, 2, -2,
    -- layer=1 filter=210 channel=107
    -6, -1, 7, 8, -2, 9, -7, 2, -9,
    -- layer=1 filter=210 channel=108
    -11, 0, -7, 10, -9, -13, 5, -9, 6,
    -- layer=1 filter=210 channel=109
    10, 9, 8, -8, 0, -5, -4, 3, 4,
    -- layer=1 filter=210 channel=110
    -1, -10, -8, -9, -4, -12, -6, -3, -8,
    -- layer=1 filter=210 channel=111
    -11, -9, -8, -15, -6, -6, 9, -4, 5,
    -- layer=1 filter=210 channel=112
    -5, -1, -10, 5, -2, -8, 2, 2, -1,
    -- layer=1 filter=210 channel=113
    9, -2, -3, 6, 8, 2, 9, 8, 2,
    -- layer=1 filter=210 channel=114
    1, -13, 5, 3, -14, -9, 6, -10, -2,
    -- layer=1 filter=210 channel=115
    -5, -2, -13, -7, -3, 2, -2, -1, 2,
    -- layer=1 filter=210 channel=116
    -1, 10, -10, -4, 7, -2, -10, 8, -7,
    -- layer=1 filter=210 channel=117
    -13, -10, 4, -2, 6, 0, -2, 7, 7,
    -- layer=1 filter=210 channel=118
    -9, 1, -7, -13, 0, 5, 6, 8, -7,
    -- layer=1 filter=210 channel=119
    -3, 0, -16, -1, -11, 1, 0, -10, -11,
    -- layer=1 filter=210 channel=120
    3, 0, 3, 6, -4, -3, -3, -2, -2,
    -- layer=1 filter=210 channel=121
    -16, -10, -13, -14, -5, -12, 6, 10, -8,
    -- layer=1 filter=210 channel=122
    -2, 3, 8, 4, -1, -9, -8, -6, -1,
    -- layer=1 filter=210 channel=123
    4, 0, -3, -2, -9, -9, -1, -8, 3,
    -- layer=1 filter=210 channel=124
    -7, 0, -5, 0, -6, -3, 0, 7, -5,
    -- layer=1 filter=210 channel=125
    -1, -5, -12, 5, -4, 2, 0, 0, 11,
    -- layer=1 filter=210 channel=126
    -8, 13, 10, -7, -10, -3, 0, 9, -2,
    -- layer=1 filter=210 channel=127
    -2, 2, -13, -7, -10, 9, -5, 3, 4,
    -- layer=1 filter=211 channel=0
    2, -1, -10, -9, -11, -11, 4, 0, 0,
    -- layer=1 filter=211 channel=1
    6, -5, -6, -3, 6, 1, 5, -2, -9,
    -- layer=1 filter=211 channel=2
    -8, -8, -7, -5, -9, -11, 6, -15, -7,
    -- layer=1 filter=211 channel=3
    4, -1, 4, 6, 3, 7, -1, -4, -7,
    -- layer=1 filter=211 channel=4
    4, 4, 1, -7, 8, -3, 0, -4, -8,
    -- layer=1 filter=211 channel=5
    -2, -1, -12, -1, -2, 0, -1, -15, -9,
    -- layer=1 filter=211 channel=6
    -2, -2, 2, 2, 12, -3, -6, -1, 3,
    -- layer=1 filter=211 channel=7
    6, -10, -15, 1, -2, 0, -7, -21, -7,
    -- layer=1 filter=211 channel=8
    -10, 9, 4, 5, -4, 9, -1, -1, -9,
    -- layer=1 filter=211 channel=9
    -2, -7, -5, 2, 0, 8, 0, -12, -10,
    -- layer=1 filter=211 channel=10
    -7, 7, -6, 0, -12, -8, 0, -13, -9,
    -- layer=1 filter=211 channel=11
    -11, 0, 1, -8, -9, -2, 0, -9, 3,
    -- layer=1 filter=211 channel=12
    -6, -1, -5, 8, 6, 4, 3, 0, -5,
    -- layer=1 filter=211 channel=13
    -4, -6, -11, -5, 4, -2, -5, -1, 8,
    -- layer=1 filter=211 channel=14
    8, 3, -4, 3, 1, 5, -7, 4, 5,
    -- layer=1 filter=211 channel=15
    -3, 5, -1, 0, 4, 3, 1, -14, 4,
    -- layer=1 filter=211 channel=16
    -9, 7, 8, -8, 4, 3, 1, 2, 1,
    -- layer=1 filter=211 channel=17
    0, 0, 7, -7, 0, 7, 5, 4, 8,
    -- layer=1 filter=211 channel=18
    1, 5, -8, -10, -8, -3, -7, 2, -2,
    -- layer=1 filter=211 channel=19
    -5, -3, -12, -10, 0, -1, 1, -1, -11,
    -- layer=1 filter=211 channel=20
    0, -7, 7, -1, -4, 5, -10, -10, -4,
    -- layer=1 filter=211 channel=21
    -11, -6, -5, -10, 0, 7, 4, 5, 0,
    -- layer=1 filter=211 channel=22
    -10, 0, -9, 4, -1, -7, 6, 2, 7,
    -- layer=1 filter=211 channel=23
    6, 8, -3, -13, -7, 3, -6, 0, -12,
    -- layer=1 filter=211 channel=24
    -2, -3, -4, -6, -3, 0, 0, 0, 5,
    -- layer=1 filter=211 channel=25
    6, 4, 3, -5, -15, -5, -10, -13, 0,
    -- layer=1 filter=211 channel=26
    7, -8, 0, -4, -12, 7, 2, 5, -6,
    -- layer=1 filter=211 channel=27
    -10, 5, 7, 0, 5, 6, 1, -7, -11,
    -- layer=1 filter=211 channel=28
    4, 10, -10, -1, -10, -10, 2, 7, 0,
    -- layer=1 filter=211 channel=29
    7, 8, 0, 6, -5, -7, -3, -10, -7,
    -- layer=1 filter=211 channel=30
    0, 5, 6, -4, -11, -12, -13, -5, 1,
    -- layer=1 filter=211 channel=31
    -9, 0, -5, 3, 4, 0, 0, -6, 10,
    -- layer=1 filter=211 channel=32
    4, -5, -8, -7, -2, -4, -5, -9, 4,
    -- layer=1 filter=211 channel=33
    1, 0, 4, 7, -1, 13, -7, 5, -6,
    -- layer=1 filter=211 channel=34
    -9, -2, -9, 5, -6, 2, -5, 0, 5,
    -- layer=1 filter=211 channel=35
    1, 1, 4, 5, -7, -7, -7, -7, 2,
    -- layer=1 filter=211 channel=36
    1, 6, 0, 8, -3, -9, -6, -1, 8,
    -- layer=1 filter=211 channel=37
    -11, 7, 6, 3, -1, 0, -14, -9, -10,
    -- layer=1 filter=211 channel=38
    -3, 1, -3, 5, 6, -2, 7, -10, -5,
    -- layer=1 filter=211 channel=39
    -3, -6, 0, -2, 7, 8, -1, -11, -1,
    -- layer=1 filter=211 channel=40
    -9, -11, -6, 0, -2, 8, -2, 0, -9,
    -- layer=1 filter=211 channel=41
    2, 0, -6, -5, 8, 1, 1, -3, 6,
    -- layer=1 filter=211 channel=42
    8, -4, 5, -7, 1, -14, -9, 2, -9,
    -- layer=1 filter=211 channel=43
    -4, -9, -6, -1, 0, -8, 0, -1, 5,
    -- layer=1 filter=211 channel=44
    9, -5, -8, 1, -1, 2, -9, -5, 6,
    -- layer=1 filter=211 channel=45
    -2, 1, 0, 7, 4, 4, -12, -6, -5,
    -- layer=1 filter=211 channel=46
    12, -1, -9, 4, -6, -4, -9, 0, -3,
    -- layer=1 filter=211 channel=47
    -7, 0, -9, -10, -8, 8, 1, -3, 5,
    -- layer=1 filter=211 channel=48
    6, -11, -2, -4, 0, -2, -5, -4, -5,
    -- layer=1 filter=211 channel=49
    0, -5, 3, -5, 8, 4, -3, 1, 7,
    -- layer=1 filter=211 channel=50
    3, 6, -7, -5, 4, -4, -8, -8, 0,
    -- layer=1 filter=211 channel=51
    0, -6, 1, 5, 0, -9, 3, 8, 1,
    -- layer=1 filter=211 channel=52
    -4, -2, 2, -5, -10, 5, 2, -10, 8,
    -- layer=1 filter=211 channel=53
    1, -7, 5, -7, -9, 8, 5, -9, -8,
    -- layer=1 filter=211 channel=54
    -1, 0, 6, -6, 0, -5, 7, 0, -13,
    -- layer=1 filter=211 channel=55
    2, -6, -7, 1, 4, -13, -11, 6, -5,
    -- layer=1 filter=211 channel=56
    0, 2, -1, 4, -8, -2, -7, 8, -1,
    -- layer=1 filter=211 channel=57
    -5, -8, 7, -5, 2, 6, -9, -1, 0,
    -- layer=1 filter=211 channel=58
    -6, 1, -3, -6, -6, -9, 8, 2, 0,
    -- layer=1 filter=211 channel=59
    -11, -1, -4, 6, 8, -12, -3, -5, -6,
    -- layer=1 filter=211 channel=60
    -1, -2, 3, 5, -7, 6, -7, 3, 1,
    -- layer=1 filter=211 channel=61
    2, 6, 0, -5, -7, 4, -6, 6, 3,
    -- layer=1 filter=211 channel=62
    -4, -10, -14, 3, 0, -9, -14, -13, -8,
    -- layer=1 filter=211 channel=63
    0, 4, 5, -7, -11, 0, 5, -12, 7,
    -- layer=1 filter=211 channel=64
    -11, -5, -3, -3, 1, 0, 2, 6, 3,
    -- layer=1 filter=211 channel=65
    0, -5, -7, 8, -2, 2, 4, -2, 8,
    -- layer=1 filter=211 channel=66
    1, 2, -8, -4, -8, 4, -11, 4, 1,
    -- layer=1 filter=211 channel=67
    1, -8, 11, -1, -8, -7, -8, -4, 11,
    -- layer=1 filter=211 channel=68
    6, -9, 10, -1, 5, -2, 3, 3, 2,
    -- layer=1 filter=211 channel=69
    7, 3, -9, -12, -12, -17, -5, -5, -6,
    -- layer=1 filter=211 channel=70
    5, -5, 0, -1, -8, -9, -3, -2, -4,
    -- layer=1 filter=211 channel=71
    9, 8, 4, -5, -6, -9, 3, -2, -11,
    -- layer=1 filter=211 channel=72
    7, 3, -11, 2, -6, -11, -2, -1, 8,
    -- layer=1 filter=211 channel=73
    4, -3, 7, 3, 9, 0, -5, -5, 1,
    -- layer=1 filter=211 channel=74
    8, -9, 5, -2, 7, 6, 4, -5, -5,
    -- layer=1 filter=211 channel=75
    -12, -1, -9, -9, -2, 0, -2, -2, -12,
    -- layer=1 filter=211 channel=76
    2, 2, -7, 7, 4, 7, 3, 1, -4,
    -- layer=1 filter=211 channel=77
    -9, -6, -12, 4, -3, 5, -8, -5, 6,
    -- layer=1 filter=211 channel=78
    -11, 5, -3, -10, 8, -7, 5, 8, -9,
    -- layer=1 filter=211 channel=79
    8, 0, 8, -3, -1, 5, -2, -11, 0,
    -- layer=1 filter=211 channel=80
    -1, 0, 0, -8, 6, -4, -1, -1, 2,
    -- layer=1 filter=211 channel=81
    -3, 4, 4, -3, 4, 1, 6, 0, 5,
    -- layer=1 filter=211 channel=82
    1, -1, -3, -5, -11, 2, 1, 6, -2,
    -- layer=1 filter=211 channel=83
    -8, -10, 2, 2, 2, -3, 6, 0, -9,
    -- layer=1 filter=211 channel=84
    -9, -10, -6, -9, 2, 0, -7, 1, 6,
    -- layer=1 filter=211 channel=85
    -3, -2, -10, 1, -10, 0, -6, -1, -9,
    -- layer=1 filter=211 channel=86
    0, -14, 4, -10, -11, 0, 1, -1, -9,
    -- layer=1 filter=211 channel=87
    -2, 0, -6, -6, -6, -8, -7, -4, -8,
    -- layer=1 filter=211 channel=88
    8, -8, 6, -12, 6, -10, -3, 9, 0,
    -- layer=1 filter=211 channel=89
    0, -7, 6, 7, 0, -8, -12, -1, 1,
    -- layer=1 filter=211 channel=90
    3, 6, 4, -1, 6, 4, -11, -11, 4,
    -- layer=1 filter=211 channel=91
    5, 1, 1, -8, -12, -6, 7, 8, -1,
    -- layer=1 filter=211 channel=92
    2, -4, -11, -7, -4, 0, -1, 1, 7,
    -- layer=1 filter=211 channel=93
    0, -1, -6, -1, 6, -4, 2, -9, 0,
    -- layer=1 filter=211 channel=94
    8, -1, -7, 8, -6, 2, -11, 1, 0,
    -- layer=1 filter=211 channel=95
    5, 8, -2, 9, 9, -2, 4, -10, 0,
    -- layer=1 filter=211 channel=96
    4, 0, -6, -10, 0, -9, -3, 2, 8,
    -- layer=1 filter=211 channel=97
    -10, 0, -10, 2, 5, -5, -10, 1, -4,
    -- layer=1 filter=211 channel=98
    -1, -7, -3, -4, -5, -5, 1, -12, -7,
    -- layer=1 filter=211 channel=99
    8, 9, 1, 0, -11, -1, -6, -3, -10,
    -- layer=1 filter=211 channel=100
    -9, 3, -1, -10, -8, 4, 3, -7, -3,
    -- layer=1 filter=211 channel=101
    -3, 3, -5, 0, 8, -5, -11, 4, -11,
    -- layer=1 filter=211 channel=102
    -2, 0, 0, 3, -9, -5, -3, 4, -2,
    -- layer=1 filter=211 channel=103
    0, 5, -7, -5, -7, -9, -1, 0, -2,
    -- layer=1 filter=211 channel=104
    -4, 8, -5, 0, -7, 7, 1, -10, 8,
    -- layer=1 filter=211 channel=105
    3, 5, -8, 0, 4, -10, -2, -4, -5,
    -- layer=1 filter=211 channel=106
    -2, 0, 4, 1, 3, 7, 5, 4, 5,
    -- layer=1 filter=211 channel=107
    -5, 8, 4, 10, -6, -10, 4, 3, 6,
    -- layer=1 filter=211 channel=108
    -4, -13, 6, -17, -8, -7, -16, 0, -10,
    -- layer=1 filter=211 channel=109
    2, 11, -6, 1, 6, 2, -1, 9, -2,
    -- layer=1 filter=211 channel=110
    -6, 2, 2, 3, -1, 3, -4, -1, 0,
    -- layer=1 filter=211 channel=111
    6, 6, -2, 2, -6, 4, 6, -9, -13,
    -- layer=1 filter=211 channel=112
    4, -8, -7, 4, 1, -11, -3, 1, 4,
    -- layer=1 filter=211 channel=113
    5, -1, -9, -3, 2, -5, 5, -5, -3,
    -- layer=1 filter=211 channel=114
    4, 3, -3, -13, -2, -9, -6, 0, 4,
    -- layer=1 filter=211 channel=115
    7, -2, -10, -7, -7, -8, -8, -2, 2,
    -- layer=1 filter=211 channel=116
    2, -10, -2, -2, -10, 4, 8, -2, -3,
    -- layer=1 filter=211 channel=117
    -5, -9, -9, -14, -5, -16, -7, 2, -1,
    -- layer=1 filter=211 channel=118
    -8, 10, 9, -6, -8, 0, -3, 10, -3,
    -- layer=1 filter=211 channel=119
    -9, 0, 2, -9, -4, -13, -7, 2, 4,
    -- layer=1 filter=211 channel=120
    -3, 1, 0, 1, 0, -3, -11, 0, 6,
    -- layer=1 filter=211 channel=121
    -10, 0, -1, -6, -8, 0, 1, -15, -8,
    -- layer=1 filter=211 channel=122
    6, -8, 1, -3, 3, -10, -2, -3, 4,
    -- layer=1 filter=211 channel=123
    -1, 1, 4, 7, -10, 5, 5, -1, 2,
    -- layer=1 filter=211 channel=124
    -3, 0, -6, 1, -3, -3, -9, 6, -8,
    -- layer=1 filter=211 channel=125
    -6, -6, -7, -7, -6, -8, -4, -3, -1,
    -- layer=1 filter=211 channel=126
    3, -2, 8, -6, -5, 8, 7, 5, 9,
    -- layer=1 filter=211 channel=127
    -10, -7, -6, 8, -2, 2, -2, 6, -3,
    -- layer=1 filter=212 channel=0
    -9, 6, 5, 0, 6, 0, -1, -3, 5,
    -- layer=1 filter=212 channel=1
    4, 4, -10, -5, -2, 8, -3, 0, 5,
    -- layer=1 filter=212 channel=2
    -11, -12, -18, 5, 2, 12, -2, 8, -8,
    -- layer=1 filter=212 channel=3
    3, 0, 0, -2, 8, 2, 8, 9, 1,
    -- layer=1 filter=212 channel=4
    -10, -9, -4, 4, -11, 8, -11, -4, 4,
    -- layer=1 filter=212 channel=5
    -10, 5, -10, -3, -3, -6, 0, 2, -6,
    -- layer=1 filter=212 channel=6
    -10, 7, -9, 4, -13, -10, 2, -2, -3,
    -- layer=1 filter=212 channel=7
    -7, 2, -7, 0, 1, 8, 7, -4, -1,
    -- layer=1 filter=212 channel=8
    -7, 0, 1, 0, 0, -1, -12, -13, 6,
    -- layer=1 filter=212 channel=9
    -15, 4, -3, 4, 12, -8, 6, -2, 0,
    -- layer=1 filter=212 channel=10
    5, 12, -6, 2, 4, -5, -2, 8, -13,
    -- layer=1 filter=212 channel=11
    5, 0, -5, 0, -4, 4, 3, 4, -7,
    -- layer=1 filter=212 channel=12
    -9, 1, 2, 0, -7, 7, 6, -10, -9,
    -- layer=1 filter=212 channel=13
    1, -3, -1, -9, -9, -3, -8, -11, 1,
    -- layer=1 filter=212 channel=14
    1, -4, -6, 9, 7, -9, -11, -1, 3,
    -- layer=1 filter=212 channel=15
    -9, 5, 7, 7, -11, -6, -5, -8, -9,
    -- layer=1 filter=212 channel=16
    2, 1, 0, -9, -10, 0, 0, 0, -9,
    -- layer=1 filter=212 channel=17
    -9, 5, -11, -4, 3, -11, 3, -6, 8,
    -- layer=1 filter=212 channel=18
    -6, -1, 2, -3, -10, 7, -7, -5, -1,
    -- layer=1 filter=212 channel=19
    -4, -7, -5, -4, -6, 3, -5, 4, -4,
    -- layer=1 filter=212 channel=20
    0, -3, 0, -2, 4, -6, -11, -7, -12,
    -- layer=1 filter=212 channel=21
    3, -7, -4, -1, 8, -4, 0, -13, -10,
    -- layer=1 filter=212 channel=22
    -9, 2, -2, -11, -6, -9, -7, -4, -4,
    -- layer=1 filter=212 channel=23
    -5, -10, -1, -11, -3, -5, -2, -7, -10,
    -- layer=1 filter=212 channel=24
    -18, -14, -4, -14, -4, -15, -7, -2, -5,
    -- layer=1 filter=212 channel=25
    -2, 2, 3, 5, -1, 4, 5, -5, 9,
    -- layer=1 filter=212 channel=26
    -6, -3, -13, -11, -2, -12, -17, -7, -3,
    -- layer=1 filter=212 channel=27
    2, 4, -3, 7, 10, -3, 0, 6, 6,
    -- layer=1 filter=212 channel=28
    -1, -9, -9, 0, -8, -11, 0, 6, 1,
    -- layer=1 filter=212 channel=29
    -7, -7, 11, 8, 8, 8, 3, 5, 6,
    -- layer=1 filter=212 channel=30
    -2, -11, -6, 0, -2, 4, 6, 8, 0,
    -- layer=1 filter=212 channel=31
    2, -14, 7, -9, 0, -8, -6, -7, 4,
    -- layer=1 filter=212 channel=32
    -2, 4, 2, -9, 3, -14, -2, 6, -4,
    -- layer=1 filter=212 channel=33
    -9, -7, 9, 0, 2, -10, 8, 9, 0,
    -- layer=1 filter=212 channel=34
    3, -8, 3, -9, -2, 2, -11, -6, 6,
    -- layer=1 filter=212 channel=35
    0, -6, -6, -11, -5, -10, 4, 0, -1,
    -- layer=1 filter=212 channel=36
    -7, 6, -10, -2, 3, -6, -4, -3, 6,
    -- layer=1 filter=212 channel=37
    -13, 0, 5, -6, -3, -15, 2, 7, -5,
    -- layer=1 filter=212 channel=38
    4, 3, -2, -3, -12, -14, 6, -4, 9,
    -- layer=1 filter=212 channel=39
    -2, -1, -9, 5, -8, -3, -9, -5, -1,
    -- layer=1 filter=212 channel=40
    -15, 1, -5, 2, -13, 0, -5, -1, 1,
    -- layer=1 filter=212 channel=41
    0, -4, -10, 3, 2, 2, -6, 0, -10,
    -- layer=1 filter=212 channel=42
    0, -15, 4, -2, 7, -6, 1, 6, 9,
    -- layer=1 filter=212 channel=43
    -4, 4, 0, -5, -11, 6, -5, 4, -10,
    -- layer=1 filter=212 channel=44
    7, 6, -12, 1, 8, 1, 5, 1, 2,
    -- layer=1 filter=212 channel=45
    -5, 5, -6, -7, -3, 6, -10, -13, 5,
    -- layer=1 filter=212 channel=46
    -8, -8, -6, 8, -2, -5, 11, -1, 2,
    -- layer=1 filter=212 channel=47
    4, 0, 0, 4, 2, 7, -7, 5, 11,
    -- layer=1 filter=212 channel=48
    -7, 7, -7, -4, -12, -7, -11, 0, 3,
    -- layer=1 filter=212 channel=49
    5, 6, -6, 3, 1, -7, -7, -11, -3,
    -- layer=1 filter=212 channel=50
    1, 1, 1, 8, -10, -6, -8, 8, -7,
    -- layer=1 filter=212 channel=51
    0, -8, -11, -3, -6, -9, -8, 2, 2,
    -- layer=1 filter=212 channel=52
    7, -10, -6, 0, -6, 6, -8, 8, -2,
    -- layer=1 filter=212 channel=53
    -1, 8, 3, 4, -10, -8, -7, 2, -8,
    -- layer=1 filter=212 channel=54
    -10, -10, 0, -1, -3, 0, -7, 7, 8,
    -- layer=1 filter=212 channel=55
    7, -1, 9, 1, -9, 2, 1, 4, -12,
    -- layer=1 filter=212 channel=56
    1, -7, -1, -8, 7, 7, 3, -1, -4,
    -- layer=1 filter=212 channel=57
    -3, -6, 8, 0, 0, 1, -1, 2, -3,
    -- layer=1 filter=212 channel=58
    -4, 7, 12, 9, -4, -10, -2, -1, -13,
    -- layer=1 filter=212 channel=59
    -5, 2, -1, 3, 0, -3, 7, 0, 5,
    -- layer=1 filter=212 channel=60
    4, 2, 3, -11, 4, -5, 1, 4, 0,
    -- layer=1 filter=212 channel=61
    6, -1, 0, -2, -4, 8, -8, -9, -7,
    -- layer=1 filter=212 channel=62
    3, -1, 6, 6, -11, -5, -2, 9, -1,
    -- layer=1 filter=212 channel=63
    -3, -8, 0, -8, -3, 7, -2, 8, -4,
    -- layer=1 filter=212 channel=64
    7, -10, -5, 6, 7, 5, 0, 8, -9,
    -- layer=1 filter=212 channel=65
    0, -9, -9, -11, -6, 2, 2, 2, 3,
    -- layer=1 filter=212 channel=66
    -5, 4, -4, -9, -8, 3, -9, -2, -3,
    -- layer=1 filter=212 channel=67
    -12, -1, -3, 1, 6, -1, 4, -8, -10,
    -- layer=1 filter=212 channel=68
    2, -11, -18, -6, 3, 8, -3, -5, -11,
    -- layer=1 filter=212 channel=69
    -5, -13, -6, 0, -9, -5, 1, 10, 8,
    -- layer=1 filter=212 channel=70
    5, -6, 0, 2, 0, 4, -8, 5, 0,
    -- layer=1 filter=212 channel=71
    -8, -2, -9, 0, -6, 0, -8, -10, -4,
    -- layer=1 filter=212 channel=72
    0, 6, -1, -7, 3, -12, 0, 0, -6,
    -- layer=1 filter=212 channel=73
    6, 2, -11, 5, -6, -8, -6, 4, -8,
    -- layer=1 filter=212 channel=74
    -9, 8, -7, -11, 0, 2, 5, -7, -1,
    -- layer=1 filter=212 channel=75
    -7, -12, 8, -2, 8, 14, 8, -9, -8,
    -- layer=1 filter=212 channel=76
    0, -11, -3, 6, 3, -1, 0, 6, 3,
    -- layer=1 filter=212 channel=77
    0, 1, -2, -7, 2, -5, -12, -2, 1,
    -- layer=1 filter=212 channel=78
    -5, -4, -10, 2, 8, -2, -10, 0, 3,
    -- layer=1 filter=212 channel=79
    -9, -2, 8, -12, -12, -10, 3, 3, -2,
    -- layer=1 filter=212 channel=80
    -4, 1, 7, -5, -6, -4, -1, 3, 9,
    -- layer=1 filter=212 channel=81
    5, -8, 3, -2, -4, 4, 3, -4, -2,
    -- layer=1 filter=212 channel=82
    -7, -7, -8, 4, -3, 3, -9, -15, 1,
    -- layer=1 filter=212 channel=83
    5, 2, 4, -7, 4, -5, -4, 5, 3,
    -- layer=1 filter=212 channel=84
    -2, -8, 3, -11, -8, -3, -7, -9, 8,
    -- layer=1 filter=212 channel=85
    -6, -5, 3, 6, 5, 3, -11, -5, -6,
    -- layer=1 filter=212 channel=86
    -13, -12, -1, -4, -8, -5, -2, -5, -10,
    -- layer=1 filter=212 channel=87
    8, -8, 3, 0, 8, 0, -12, 6, 1,
    -- layer=1 filter=212 channel=88
    -6, -3, 0, -10, -11, -13, -9, -7, -11,
    -- layer=1 filter=212 channel=89
    7, -12, -4, -7, -10, 7, 8, 0, -10,
    -- layer=1 filter=212 channel=90
    -8, -4, -5, 6, 0, 0, -5, -4, -9,
    -- layer=1 filter=212 channel=91
    -3, -7, 1, 3, -12, 5, -11, -11, -6,
    -- layer=1 filter=212 channel=92
    -4, 4, -3, -1, -11, -4, -6, 2, 6,
    -- layer=1 filter=212 channel=93
    2, -12, -11, -1, -6, 1, -1, -7, 0,
    -- layer=1 filter=212 channel=94
    -5, -11, 0, -7, -5, 3, 6, 7, -6,
    -- layer=1 filter=212 channel=95
    1, 0, -5, 2, 8, 6, 11, -8, -9,
    -- layer=1 filter=212 channel=96
    1, -3, -4, -5, -1, -2, -2, 7, -6,
    -- layer=1 filter=212 channel=97
    3, 0, 0, -11, -1, 4, -10, 4, 2,
    -- layer=1 filter=212 channel=98
    8, -8, -1, 4, -9, -13, -14, -3, -5,
    -- layer=1 filter=212 channel=99
    3, 3, -4, -10, 3, 7, -2, 7, 7,
    -- layer=1 filter=212 channel=100
    -8, -1, 5, 2, 8, -5, -8, -8, -6,
    -- layer=1 filter=212 channel=101
    0, -3, -4, -6, -6, -8, 8, 5, 5,
    -- layer=1 filter=212 channel=102
    7, 8, 1, -9, 1, 0, 0, 1, -6,
    -- layer=1 filter=212 channel=103
    -1, 5, -8, -9, -14, -9, 7, 0, -5,
    -- layer=1 filter=212 channel=104
    0, -4, 2, -2, 7, -1, 3, 8, -4,
    -- layer=1 filter=212 channel=105
    7, 6, 5, -9, 1, -12, 5, -5, -5,
    -- layer=1 filter=212 channel=106
    -1, -11, -11, 4, -16, 7, -12, 6, -9,
    -- layer=1 filter=212 channel=107
    7, 0, 2, -5, -10, -10, -8, 1, -9,
    -- layer=1 filter=212 channel=108
    0, 0, 0, -19, -6, -14, -6, -10, 0,
    -- layer=1 filter=212 channel=109
    -2, -7, -10, 7, 5, 2, 6, -5, 4,
    -- layer=1 filter=212 channel=110
    -1, 9, -3, 1, 8, 0, 2, 3, 8,
    -- layer=1 filter=212 channel=111
    -5, -2, 10, -13, 0, -1, 0, 3, -8,
    -- layer=1 filter=212 channel=112
    8, -3, -6, -2, -10, 6, -7, -6, 0,
    -- layer=1 filter=212 channel=113
    -8, -8, 7, -6, -4, 7, 5, -7, 2,
    -- layer=1 filter=212 channel=114
    4, 6, 2, -3, 3, -14, -4, -1, 8,
    -- layer=1 filter=212 channel=115
    -4, -11, 2, 0, 8, -1, 4, -12, 0,
    -- layer=1 filter=212 channel=116
    -2, 5, -4, -5, -7, 0, 9, -5, 6,
    -- layer=1 filter=212 channel=117
    1, -6, 5, -4, -8, 5, 6, 7, -12,
    -- layer=1 filter=212 channel=118
    -6, -8, -9, -12, 7, 1, 3, -1, -6,
    -- layer=1 filter=212 channel=119
    -7, -1, -5, -5, -8, -4, -11, -11, 9,
    -- layer=1 filter=212 channel=120
    -10, 0, -10, -3, -2, -12, 0, 0, 1,
    -- layer=1 filter=212 channel=121
    0, -12, -8, 12, 0, -1, 1, -9, -4,
    -- layer=1 filter=212 channel=122
    0, 7, -8, -2, 8, 0, -10, 5, 8,
    -- layer=1 filter=212 channel=123
    0, 1, -8, 7, -6, 3, -10, -6, -11,
    -- layer=1 filter=212 channel=124
    2, -4, -8, -8, 4, 9, -7, -5, 0,
    -- layer=1 filter=212 channel=125
    -1, -8, 0, 0, -5, -6, -1, -11, -3,
    -- layer=1 filter=212 channel=126
    -10, -2, 4, 2, -1, -1, -12, -11, 0,
    -- layer=1 filter=212 channel=127
    -9, 6, -1, -10, 1, 8, -1, -7, -1,
    -- layer=1 filter=213 channel=0
    7, 3, -3, -1, 5, -5, 4, -2, -10,
    -- layer=1 filter=213 channel=1
    2, -1, 2, 5, -2, 0, 3, 6, -9,
    -- layer=1 filter=213 channel=2
    2, -1, -12, -1, -1, -4, 1, 2, -7,
    -- layer=1 filter=213 channel=3
    9, 8, -8, -7, 5, 5, 6, -6, 7,
    -- layer=1 filter=213 channel=4
    -1, 1, -4, -10, -6, -9, 8, -9, -6,
    -- layer=1 filter=213 channel=5
    -15, 2, -6, -7, -9, 6, 1, -13, 2,
    -- layer=1 filter=213 channel=6
    -1, 6, 5, 0, -12, -18, -13, -12, -8,
    -- layer=1 filter=213 channel=7
    -17, 0, -9, -14, -7, -14, -6, -3, -12,
    -- layer=1 filter=213 channel=8
    -8, -10, 3, 1, 3, 3, 3, -3, 4,
    -- layer=1 filter=213 channel=9
    -5, -7, -4, 4, 1, -2, -10, -2, -4,
    -- layer=1 filter=213 channel=10
    -13, -1, -10, -8, -10, 0, 0, 2, 0,
    -- layer=1 filter=213 channel=11
    -2, -8, -2, -15, -13, -12, -6, 6, -8,
    -- layer=1 filter=213 channel=12
    -4, -6, 1, -8, -5, -7, 0, 2, -12,
    -- layer=1 filter=213 channel=13
    1, -6, -11, -2, 7, -7, -7, -8, -9,
    -- layer=1 filter=213 channel=14
    2, 1, 3, -3, 7, 3, 5, -17, -15,
    -- layer=1 filter=213 channel=15
    -9, 0, -8, -3, 6, -10, -5, 4, -11,
    -- layer=1 filter=213 channel=16
    6, 5, -3, -12, -7, -8, 2, -12, -4,
    -- layer=1 filter=213 channel=17
    -1, 3, -4, -8, 0, 0, 8, -2, -4,
    -- layer=1 filter=213 channel=18
    0, -5, -9, -11, -17, 5, 1, 1, -2,
    -- layer=1 filter=213 channel=19
    0, -2, 5, 2, -3, -2, -10, 1, 3,
    -- layer=1 filter=213 channel=20
    1, -1, -6, -10, 2, 9, 8, -7, -8,
    -- layer=1 filter=213 channel=21
    -7, -1, 0, -3, -5, -10, -23, 2, -2,
    -- layer=1 filter=213 channel=22
    4, -9, -5, -2, -11, 5, -4, -1, 1,
    -- layer=1 filter=213 channel=23
    1, -2, 5, 0, -1, -4, 7, -3, -9,
    -- layer=1 filter=213 channel=24
    1, -8, 5, -1, -1, -13, -18, -17, -3,
    -- layer=1 filter=213 channel=25
    -16, -3, -11, -11, -8, -6, -4, -12, 2,
    -- layer=1 filter=213 channel=26
    -14, -3, 5, -1, -4, -3, -23, -9, 3,
    -- layer=1 filter=213 channel=27
    4, 11, 16, -24, -2, 9, -3, -1, -10,
    -- layer=1 filter=213 channel=28
    -7, 2, -10, 7, 6, -10, -2, 0, -6,
    -- layer=1 filter=213 channel=29
    1, 13, 0, 0, 2, 1, 6, -4, 16,
    -- layer=1 filter=213 channel=30
    -20, -5, -5, 5, -1, 0, -2, 2, -15,
    -- layer=1 filter=213 channel=31
    7, 8, 0, -14, -6, -5, 10, 1, -8,
    -- layer=1 filter=213 channel=32
    -11, -8, -7, -11, 0, -16, -7, -10, -3,
    -- layer=1 filter=213 channel=33
    -9, 2, -7, -10, -2, -7, -4, 7, -1,
    -- layer=1 filter=213 channel=34
    3, -6, -6, -5, 3, -3, 7, -10, 3,
    -- layer=1 filter=213 channel=35
    -11, -11, -3, 6, 9, 8, 5, -7, -5,
    -- layer=1 filter=213 channel=36
    -4, 4, -10, 0, 2, 4, -4, -12, -11,
    -- layer=1 filter=213 channel=37
    -9, 0, 1, -11, -1, 3, -6, -12, -7,
    -- layer=1 filter=213 channel=38
    -10, 6, 0, -6, -17, -9, -1, 4, -16,
    -- layer=1 filter=213 channel=39
    1, -8, 6, 0, -8, -10, 8, 2, 0,
    -- layer=1 filter=213 channel=40
    -17, -3, 0, 2, -10, -12, -11, -6, 0,
    -- layer=1 filter=213 channel=41
    3, -3, 3, 0, -1, -1, -7, -11, 8,
    -- layer=1 filter=213 channel=42
    3, 0, -11, -14, -5, 3, 6, -9, -17,
    -- layer=1 filter=213 channel=43
    2, 4, -3, 2, 4, -11, 2, -1, -7,
    -- layer=1 filter=213 channel=44
    0, -1, -9, 3, 2, 0, -9, 2, -11,
    -- layer=1 filter=213 channel=45
    -4, -8, 0, -8, 6, -3, -10, 1, -7,
    -- layer=1 filter=213 channel=46
    -13, 8, 0, 9, 0, -4, -11, -21, -8,
    -- layer=1 filter=213 channel=47
    -17, -9, -6, -2, 4, 6, -3, 1, 3,
    -- layer=1 filter=213 channel=48
    0, 4, 0, -6, -11, -1, 9, -4, -9,
    -- layer=1 filter=213 channel=49
    -8, -8, -1, 0, 3, 4, -8, -2, -13,
    -- layer=1 filter=213 channel=50
    8, -10, 10, -9, 4, -7, 2, 6, -2,
    -- layer=1 filter=213 channel=51
    -12, 0, 0, 0, 1, -8, 0, 0, -7,
    -- layer=1 filter=213 channel=52
    -6, 2, 2, 6, -8, -2, 0, -7, -4,
    -- layer=1 filter=213 channel=53
    -2, 8, 2, 8, 4, 9, -8, -8, 7,
    -- layer=1 filter=213 channel=54
    6, -7, -6, 0, 0, 0, 0, 4, -3,
    -- layer=1 filter=213 channel=55
    -4, 10, 4, -17, -7, 1, -9, -9, 0,
    -- layer=1 filter=213 channel=56
    -3, 11, -4, 7, -1, -10, 6, -5, -10,
    -- layer=1 filter=213 channel=57
    -11, -10, -3, -1, 5, 0, 3, 4, -4,
    -- layer=1 filter=213 channel=58
    -14, -7, -5, -12, -1, -15, -7, -15, -5,
    -- layer=1 filter=213 channel=59
    -8, -4, 0, -10, -9, -8, -5, 7, 7,
    -- layer=1 filter=213 channel=60
    9, 2, 0, 9, 0, -12, -9, 0, 3,
    -- layer=1 filter=213 channel=61
    -4, 5, 2, -11, -7, 8, -3, 0, -6,
    -- layer=1 filter=213 channel=62
    8, -9, -6, -2, 2, -5, -5, -9, 0,
    -- layer=1 filter=213 channel=63
    5, 10, 0, -4, -1, 0, -2, -9, 5,
    -- layer=1 filter=213 channel=64
    2, -6, -3, 2, -5, -6, 0, 0, -4,
    -- layer=1 filter=213 channel=65
    -9, -9, 9, 6, 6, 8, -8, 3, 9,
    -- layer=1 filter=213 channel=66
    0, -10, 3, -8, -3, -8, -4, 4, 0,
    -- layer=1 filter=213 channel=67
    0, -4, 4, 5, -2, -7, 4, -10, 3,
    -- layer=1 filter=213 channel=68
    4, 4, 3, -11, 4, -4, -12, -5, -7,
    -- layer=1 filter=213 channel=69
    -7, -3, -8, -17, -8, -3, -26, -16, -9,
    -- layer=1 filter=213 channel=70
    5, -1, -2, -2, 1, -9, -9, -11, -7,
    -- layer=1 filter=213 channel=71
    -3, -10, 1, -9, 0, 1, -14, -9, -13,
    -- layer=1 filter=213 channel=72
    4, -4, -7, -5, -12, 8, -3, 9, -4,
    -- layer=1 filter=213 channel=73
    2, 6, 1, 1, 9, 8, 5, 5, 7,
    -- layer=1 filter=213 channel=74
    1, -2, 5, 6, 2, -6, 6, 0, 5,
    -- layer=1 filter=213 channel=75
    4, -10, -8, -12, -3, -5, 4, -7, 0,
    -- layer=1 filter=213 channel=76
    -6, -1, 8, 2, 2, 3, 4, -10, 1,
    -- layer=1 filter=213 channel=77
    1, -5, 3, 2, 4, 6, 8, -5, -2,
    -- layer=1 filter=213 channel=78
    5, -8, 7, -2, 4, -9, -2, -3, 8,
    -- layer=1 filter=213 channel=79
    -5, 2, 6, -13, -5, -1, 5, -10, -7,
    -- layer=1 filter=213 channel=80
    0, 0, 1, 8, -9, -11, -5, 5, 0,
    -- layer=1 filter=213 channel=81
    6, -2, -2, 6, 7, 4, 4, 0, 2,
    -- layer=1 filter=213 channel=82
    -15, -7, -3, 0, -14, 1, -10, 4, -13,
    -- layer=1 filter=213 channel=83
    -10, 2, -3, -1, 6, 9, 6, -1, -9,
    -- layer=1 filter=213 channel=84
    1, -4, -2, -8, -15, 2, -4, -1, -3,
    -- layer=1 filter=213 channel=85
    -9, -5, 12, -11, -4, 4, -2, -10, -12,
    -- layer=1 filter=213 channel=86
    -1, -14, -3, 0, -2, -9, -9, 0, -3,
    -- layer=1 filter=213 channel=87
    7, 3, -8, 5, 4, 0, -1, -9, -5,
    -- layer=1 filter=213 channel=88
    -3, 1, -7, 5, -10, -4, -14, -19, -18,
    -- layer=1 filter=213 channel=89
    -4, -6, -8, -14, -6, -13, -10, -8, 3,
    -- layer=1 filter=213 channel=90
    -4, 0, 4, 0, 1, -5, -9, -8, 2,
    -- layer=1 filter=213 channel=91
    -19, -4, -8, -5, -14, -15, -7, 0, -5,
    -- layer=1 filter=213 channel=92
    -3, 9, 2, -9, -1, 8, -3, 0, 8,
    -- layer=1 filter=213 channel=93
    -12, 0, -11, 2, 5, -12, 0, -2, -10,
    -- layer=1 filter=213 channel=94
    -3, -3, -1, -11, -8, -2, 7, -9, -5,
    -- layer=1 filter=213 channel=95
    0, 6, -5, -13, 0, 6, -1, 3, 0,
    -- layer=1 filter=213 channel=96
    7, 3, 9, -10, -9, 1, -6, 0, -6,
    -- layer=1 filter=213 channel=97
    -8, 7, 4, -2, -10, 2, -3, 9, 4,
    -- layer=1 filter=213 channel=98
    -3, -11, 0, -23, -9, -10, -5, -4, 8,
    -- layer=1 filter=213 channel=99
    -4, -2, -9, -1, 5, 5, 7, -7, -3,
    -- layer=1 filter=213 channel=100
    4, -8, 9, 1, -7, -2, 8, -10, -5,
    -- layer=1 filter=213 channel=101
    -1, -8, -2, -5, 6, -11, -10, -7, -2,
    -- layer=1 filter=213 channel=102
    -4, 2, -8, 3, 2, 1, -7, -3, -1,
    -- layer=1 filter=213 channel=103
    1, 8, 4, 5, -15, 3, -9, 6, -11,
    -- layer=1 filter=213 channel=104
    3, -10, -7, -11, 6, 0, -10, 0, -5,
    -- layer=1 filter=213 channel=105
    3, -1, 3, 3, 0, -4, -1, -8, 0,
    -- layer=1 filter=213 channel=106
    -8, -12, -11, -20, -11, -14, -15, 0, -10,
    -- layer=1 filter=213 channel=107
    0, -7, 5, -3, -6, 1, 0, -3, 3,
    -- layer=1 filter=213 channel=108
    -17, 1, 0, -3, -6, -14, -17, -4, 4,
    -- layer=1 filter=213 channel=109
    1, -8, 3, -8, -6, -7, 3, -1, 4,
    -- layer=1 filter=213 channel=110
    3, -5, 4, -2, -2, 0, -9, -5, -7,
    -- layer=1 filter=213 channel=111
    -2, -1, 5, 2, -11, 6, -15, -9, -10,
    -- layer=1 filter=213 channel=112
    -4, -2, 7, -8, -5, -4, 3, 3, 9,
    -- layer=1 filter=213 channel=113
    -11, -5, -9, 6, 3, 0, 0, -8, -9,
    -- layer=1 filter=213 channel=114
    -11, -18, 0, -4, -14, 2, -11, -16, -2,
    -- layer=1 filter=213 channel=115
    -12, 0, 9, -10, -1, 2, 9, -10, -4,
    -- layer=1 filter=213 channel=116
    -10, 8, -9, -8, 0, -6, 0, 1, 2,
    -- layer=1 filter=213 channel=117
    -2, -7, -8, -15, -2, 4, 3, -6, -1,
    -- layer=1 filter=213 channel=118
    -10, 4, -12, -7, -11, 0, -15, -12, -11,
    -- layer=1 filter=213 channel=119
    -18, 4, -6, 4, -3, -13, -7, 0, -11,
    -- layer=1 filter=213 channel=120
    -13, 0, 1, -3, -13, 5, -4, 1, -1,
    -- layer=1 filter=213 channel=121
    -9, -7, 8, -10, -4, 10, -4, -8, -7,
    -- layer=1 filter=213 channel=122
    -7, 10, 8, -9, 1, 8, -9, 0, 0,
    -- layer=1 filter=213 channel=123
    -5, -2, 9, -7, -9, -4, -1, 3, 2,
    -- layer=1 filter=213 channel=124
    4, 7, -3, 3, -2, -9, 5, 5, -2,
    -- layer=1 filter=213 channel=125
    1, -8, 1, 0, 5, -1, 0, 6, -7,
    -- layer=1 filter=213 channel=126
    -10, -11, 1, -8, -11, 4, 4, 3, 10,
    -- layer=1 filter=213 channel=127
    2, -3, -11, -5, -2, 4, -12, -1, -5,
    -- layer=1 filter=214 channel=0
    -8, 6, 0, -5, 1, 3, -10, -3, -10,
    -- layer=1 filter=214 channel=1
    -11, -5, 2, -4, 5, -6, 7, -6, 3,
    -- layer=1 filter=214 channel=2
    -3, 1, -1, 9, 6, 12, 2, 17, 11,
    -- layer=1 filter=214 channel=3
    -2, 0, -8, 7, -5, -4, 4, -9, -5,
    -- layer=1 filter=214 channel=4
    0, -7, 5, 9, 0, -3, -10, 5, 4,
    -- layer=1 filter=214 channel=5
    -3, -6, -14, 0, -1, 9, -6, -4, 1,
    -- layer=1 filter=214 channel=6
    0, 5, 8, -6, -6, -4, -8, 2, -7,
    -- layer=1 filter=214 channel=7
    -11, -8, -3, -6, -1, 13, 1, 5, 0,
    -- layer=1 filter=214 channel=8
    -11, -2, -3, 9, 6, 2, -11, 0, -4,
    -- layer=1 filter=214 channel=9
    5, 0, -12, -10, 0, -6, -1, -3, -7,
    -- layer=1 filter=214 channel=10
    -5, -11, 7, 2, -2, 7, 4, -8, 0,
    -- layer=1 filter=214 channel=11
    3, -5, -10, 4, -7, 6, -8, 1, -5,
    -- layer=1 filter=214 channel=12
    -6, 9, 2, -4, 3, 6, 1, 0, 4,
    -- layer=1 filter=214 channel=13
    3, -9, -9, 3, 5, 0, 3, -5, 4,
    -- layer=1 filter=214 channel=14
    0, 1, -12, -5, -9, 0, -3, -5, 5,
    -- layer=1 filter=214 channel=15
    -10, -11, -1, 5, -8, 5, -9, 6, -4,
    -- layer=1 filter=214 channel=16
    -15, 2, -5, 0, -2, -10, -4, 4, -4,
    -- layer=1 filter=214 channel=17
    6, 2, 6, -3, 1, -1, 0, -4, -9,
    -- layer=1 filter=214 channel=18
    -5, 0, -10, 4, -1, -8, 2, -4, 6,
    -- layer=1 filter=214 channel=19
    0, 0, 6, -7, 1, -3, 6, 0, -11,
    -- layer=1 filter=214 channel=20
    -11, 7, -10, -7, -3, -5, -4, -6, -9,
    -- layer=1 filter=214 channel=21
    -13, 5, 0, 0, -6, -5, 0, 3, -9,
    -- layer=1 filter=214 channel=22
    -4, -10, -8, -5, -7, -5, -9, 7, -8,
    -- layer=1 filter=214 channel=23
    -12, 4, 3, -2, -7, 1, -1, -8, 2,
    -- layer=1 filter=214 channel=24
    5, 3, -6, -12, 2, -11, -1, -3, 0,
    -- layer=1 filter=214 channel=25
    4, -15, 1, -7, 1, -1, -4, 5, 1,
    -- layer=1 filter=214 channel=26
    5, -12, 3, 0, 0, -8, -10, 2, 4,
    -- layer=1 filter=214 channel=27
    -1, 12, 11, -7, 10, 7, 10, -7, 5,
    -- layer=1 filter=214 channel=28
    -2, -6, -15, 1, -10, -10, 2, -10, -13,
    -- layer=1 filter=214 channel=29
    2, 5, 8, 5, -4, -6, -9, 5, -6,
    -- layer=1 filter=214 channel=30
    -18, -1, -13, -5, -14, -11, -9, -17, -14,
    -- layer=1 filter=214 channel=31
    0, 0, -14, -10, -1, -15, -16, 0, 2,
    -- layer=1 filter=214 channel=32
    -2, -13, -1, 0, -9, 6, -1, -1, -2,
    -- layer=1 filter=214 channel=33
    -2, -1, 3, 12, 6, -1, -3, -7, -6,
    -- layer=1 filter=214 channel=34
    6, -4, -10, -9, -10, -5, -10, -8, -9,
    -- layer=1 filter=214 channel=35
    1, -3, 7, 1, 7, -10, -11, -3, 5,
    -- layer=1 filter=214 channel=36
    -4, 1, 0, -4, 5, -5, -3, 1, -7,
    -- layer=1 filter=214 channel=37
    -4, -17, -16, 1, -2, 8, -12, 2, 8,
    -- layer=1 filter=214 channel=38
    3, 6, -9, -6, 0, 3, -4, 5, -9,
    -- layer=1 filter=214 channel=39
    4, -11, -2, -7, -7, -7, -12, 0, 0,
    -- layer=1 filter=214 channel=40
    -20, -4, -12, -18, -20, -16, -9, -5, 9,
    -- layer=1 filter=214 channel=41
    6, -1, 9, -6, -6, -3, -6, 1, -4,
    -- layer=1 filter=214 channel=42
    0, 1, 5, 0, 8, 11, 8, 14, 7,
    -- layer=1 filter=214 channel=43
    -6, 8, -11, -2, -8, 1, -2, 9, -12,
    -- layer=1 filter=214 channel=44
    -4, 6, -7, 6, 1, -3, 5, -2, 2,
    -- layer=1 filter=214 channel=45
    -3, -11, -11, 0, 0, -13, -4, 0, -8,
    -- layer=1 filter=214 channel=46
    -13, -4, -7, -4, 14, 14, -15, 11, 0,
    -- layer=1 filter=214 channel=47
    3, -6, 8, -6, -4, 1, -8, 8, 5,
    -- layer=1 filter=214 channel=48
    -11, -7, 1, 1, 3, 0, 1, -9, -5,
    -- layer=1 filter=214 channel=49
    -8, -5, -2, -11, 2, -3, 5, -5, 3,
    -- layer=1 filter=214 channel=50
    -11, 4, -4, 3, -4, -4, -12, -9, 0,
    -- layer=1 filter=214 channel=51
    4, 0, -7, -6, -8, -3, 5, 3, -1,
    -- layer=1 filter=214 channel=52
    -7, -5, -7, 5, -7, -7, 5, -2, 12,
    -- layer=1 filter=214 channel=53
    -8, -8, 7, 8, 4, -10, 0, -8, 7,
    -- layer=1 filter=214 channel=54
    4, -11, 6, 3, 4, 8, -11, 6, 3,
    -- layer=1 filter=214 channel=55
    -7, 7, 7, -4, 2, -10, 5, -5, 7,
    -- layer=1 filter=214 channel=56
    5, 4, -1, -7, -2, 0, 0, 7, 4,
    -- layer=1 filter=214 channel=57
    -8, -4, -13, -6, -1, -7, 0, 7, 2,
    -- layer=1 filter=214 channel=58
    -8, -10, 0, 4, 0, -7, -4, 10, 5,
    -- layer=1 filter=214 channel=59
    4, 4, -7, 7, -5, -5, -7, 6, -8,
    -- layer=1 filter=214 channel=60
    6, -2, 8, 0, 9, -7, -4, 3, -2,
    -- layer=1 filter=214 channel=61
    -5, -6, -8, -11, 3, -6, 5, 4, 2,
    -- layer=1 filter=214 channel=62
    -9, -4, -18, -11, 1, 8, -3, 9, -1,
    -- layer=1 filter=214 channel=63
    -8, -9, 0, 4, -3, 1, -5, -5, -7,
    -- layer=1 filter=214 channel=64
    -5, -2, 4, -8, -11, 2, -2, -9, -8,
    -- layer=1 filter=214 channel=65
    -9, -2, 6, -4, 0, 2, 2, 4, 4,
    -- layer=1 filter=214 channel=66
    -1, 0, 4, 1, 8, 0, 5, 4, 0,
    -- layer=1 filter=214 channel=67
    -7, -16, -14, 1, 5, 3, -9, -6, 6,
    -- layer=1 filter=214 channel=68
    -5, 0, -6, -9, -10, 7, 3, 4, -8,
    -- layer=1 filter=214 channel=69
    -11, 2, -11, 8, 12, 7, -12, -3, 7,
    -- layer=1 filter=214 channel=70
    -11, -13, -11, -11, 0, -4, -10, -6, -7,
    -- layer=1 filter=214 channel=71
    -12, -10, 3, -2, -9, -4, -3, -7, 0,
    -- layer=1 filter=214 channel=72
    -2, 8, -6, 0, 8, 4, 6, 0, 7,
    -- layer=1 filter=214 channel=73
    8, -5, 6, 7, -4, 6, -2, 5, -10,
    -- layer=1 filter=214 channel=74
    3, 0, 0, -12, -10, 4, 2, -6, -8,
    -- layer=1 filter=214 channel=75
    -3, 2, -12, 3, -8, -16, -12, -5, -6,
    -- layer=1 filter=214 channel=76
    3, -8, 3, -8, -1, 3, 0, 4, -9,
    -- layer=1 filter=214 channel=77
    6, 0, 0, -8, 6, -7, 5, -5, -8,
    -- layer=1 filter=214 channel=78
    -6, -2, -1, -5, 1, 6, 7, -9, -3,
    -- layer=1 filter=214 channel=79
    -10, 4, 0, -3, 3, 0, 1, 0, -13,
    -- layer=1 filter=214 channel=80
    9, -2, -4, -7, 1, 2, 1, 2, 9,
    -- layer=1 filter=214 channel=81
    -10, 5, -11, -10, -9, 0, -5, 3, -2,
    -- layer=1 filter=214 channel=82
    2, 2, -8, 5, -2, -9, -3, -3, 1,
    -- layer=1 filter=214 channel=83
    -9, 4, 0, -5, 3, -9, 6, 5, 3,
    -- layer=1 filter=214 channel=84
    -9, 5, -8, -14, -15, -14, -4, 2, 11,
    -- layer=1 filter=214 channel=85
    10, 1, -2, 0, 8, 3, 10, -8, -9,
    -- layer=1 filter=214 channel=86
    0, 6, -4, 0, -8, -7, 4, -8, -2,
    -- layer=1 filter=214 channel=87
    10, 2, -6, -9, 1, 11, 6, 0, 6,
    -- layer=1 filter=214 channel=88
    -13, 2, 0, -2, -4, -15, -4, -10, 0,
    -- layer=1 filter=214 channel=89
    -3, -2, 2, -5, -2, -10, -2, -12, 0,
    -- layer=1 filter=214 channel=90
    5, 3, 8, 0, 1, 1, -8, 7, -11,
    -- layer=1 filter=214 channel=91
    -6, -4, -9, -8, 5, -14, 2, -13, -12,
    -- layer=1 filter=214 channel=92
    -6, 5, -6, -5, -7, 9, -2, -5, 5,
    -- layer=1 filter=214 channel=93
    0, 2, 5, -8, -5, 0, -12, -13, -8,
    -- layer=1 filter=214 channel=94
    6, -2, -7, 5, -10, -7, 7, -7, -8,
    -- layer=1 filter=214 channel=95
    -8, -13, 4, 2, -7, -11, -10, -10, -7,
    -- layer=1 filter=214 channel=96
    -2, -1, -7, -11, -4, 9, 4, -5, -6,
    -- layer=1 filter=214 channel=97
    5, -11, 0, 0, 4, -5, -3, -7, 1,
    -- layer=1 filter=214 channel=98
    0, 3, -6, -16, 4, -13, -4, -3, -14,
    -- layer=1 filter=214 channel=99
    -7, 0, 3, 2, 9, -5, 0, -3, 1,
    -- layer=1 filter=214 channel=100
    0, -10, 3, -3, -4, 5, -11, 0, -5,
    -- layer=1 filter=214 channel=101
    4, 0, -6, 3, 4, -2, -2, -1, 6,
    -- layer=1 filter=214 channel=102
    -9, -2, -12, -8, -2, 1, 0, -4, 0,
    -- layer=1 filter=214 channel=103
    -2, 4, -9, -13, 0, 7, -5, -7, 3,
    -- layer=1 filter=214 channel=104
    7, -7, 5, -3, 6, 8, 9, 7, -8,
    -- layer=1 filter=214 channel=105
    4, 8, -6, -10, 2, -4, -10, 8, -5,
    -- layer=1 filter=214 channel=106
    -3, -7, -11, -8, -1, 2, 3, -10, -3,
    -- layer=1 filter=214 channel=107
    -8, 1, 11, -2, 4, 0, 7, -9, -3,
    -- layer=1 filter=214 channel=108
    -8, 5, -1, 1, -1, -1, 6, -4, 0,
    -- layer=1 filter=214 channel=109
    0, 0, -6, -3, -9, -3, 10, 4, -4,
    -- layer=1 filter=214 channel=110
    -6, 4, -7, 2, -7, -9, -11, 8, -3,
    -- layer=1 filter=214 channel=111
    -11, 4, -6, 6, 5, -2, -5, 7, 6,
    -- layer=1 filter=214 channel=112
    -1, -10, -2, -8, 4, 2, 4, 7, -8,
    -- layer=1 filter=214 channel=113
    7, -12, 4, 3, -11, -11, 6, -4, -10,
    -- layer=1 filter=214 channel=114
    -8, -5, 2, -7, -8, 12, -15, -8, 5,
    -- layer=1 filter=214 channel=115
    5, -4, 0, -10, 5, -2, -2, 0, 5,
    -- layer=1 filter=214 channel=116
    -4, 0, -4, -9, 5, 0, 4, 1, -9,
    -- layer=1 filter=214 channel=117
    0, -6, -4, -7, -6, 1, -2, -4, -1,
    -- layer=1 filter=214 channel=118
    -10, -7, 0, -8, -4, -11, -15, -11, -8,
    -- layer=1 filter=214 channel=119
    4, -16, -7, -3, 0, -15, 3, 8, 9,
    -- layer=1 filter=214 channel=120
    5, 0, -13, -10, -6, 3, 6, -1, 2,
    -- layer=1 filter=214 channel=121
    -5, 3, 3, -2, -2, 4, 6, -8, 11,
    -- layer=1 filter=214 channel=122
    0, -7, -6, -8, -7, -6, -3, 9, -6,
    -- layer=1 filter=214 channel=123
    0, 0, 7, 3, -8, 2, -12, -11, 0,
    -- layer=1 filter=214 channel=124
    2, 9, 1, 2, 5, -6, 10, 13, 10,
    -- layer=1 filter=214 channel=125
    4, -19, -5, -3, 9, 6, -1, 0, 8,
    -- layer=1 filter=214 channel=126
    6, 9, 0, -2, 3, -8, 5, 4, 1,
    -- layer=1 filter=214 channel=127
    -11, -6, -6, 1, -7, -11, -17, 1, -4,
    -- layer=1 filter=215 channel=0
    -20, 24, 11, -19, 25, 19, -14, -7, 19,
    -- layer=1 filter=215 channel=1
    -11, -4, 17, 5, -29, 3, -16, -10, -11,
    -- layer=1 filter=215 channel=2
    -11, -25, -38, -19, -11, -26, 9, 0, -5,
    -- layer=1 filter=215 channel=3
    -7, -6, 11, -5, -6, 2, 6, 6, 7,
    -- layer=1 filter=215 channel=4
    10, 10, -5, -3, -5, 3, -3, 8, 9,
    -- layer=1 filter=215 channel=5
    -11, 15, 34, 23, -8, 14, 10, 16, 1,
    -- layer=1 filter=215 channel=6
    74, 11, 1, 85, -19, -61, 80, -53, -51,
    -- layer=1 filter=215 channel=7
    45, 64, 43, 33, 68, 44, 12, 66, 50,
    -- layer=1 filter=215 channel=8
    -17, 21, 26, 11, -11, 15, -20, 14, -9,
    -- layer=1 filter=215 channel=9
    -48, -62, -43, -17, -69, -19, 7, 40, -1,
    -- layer=1 filter=215 channel=10
    39, 65, 40, 17, 56, 38, 3, 57, 51,
    -- layer=1 filter=215 channel=11
    -8, 10, 16, -23, 0, 18, -9, 3, 13,
    -- layer=1 filter=215 channel=12
    32, 58, 25, -32, -6, -12, -28, 0, -44,
    -- layer=1 filter=215 channel=13
    3, -12, -12, 24, -23, -8, 16, -43, -22,
    -- layer=1 filter=215 channel=14
    13, 42, 38, 14, 62, 40, -48, 46, 12,
    -- layer=1 filter=215 channel=15
    -41, -24, 30, 15, -35, 39, -37, -20, -22,
    -- layer=1 filter=215 channel=16
    -19, 7, 9, -4, 5, 2, -8, 24, -15,
    -- layer=1 filter=215 channel=17
    -11, 24, 28, -35, -5, 20, -18, -28, 17,
    -- layer=1 filter=215 channel=18
    9, 20, -10, -41, 24, 49, 3, 32, 20,
    -- layer=1 filter=215 channel=19
    -34, -86, -39, -52, -30, -24, -15, -18, -12,
    -- layer=1 filter=215 channel=20
    -5, -21, -3, -7, -28, -4, -20, -34, -34,
    -- layer=1 filter=215 channel=21
    11, -18, -30, 21, -44, -41, 4, -28, -32,
    -- layer=1 filter=215 channel=22
    6, -2, -10, 35, -33, -11, -9, -34, -44,
    -- layer=1 filter=215 channel=23
    -33, -32, 43, -19, 1, 26, -48, 13, 5,
    -- layer=1 filter=215 channel=24
    -36, -25, -19, -36, -31, -13, -9, -37, 2,
    -- layer=1 filter=215 channel=25
    17, 23, 33, 12, 27, -6, -6, 25, 11,
    -- layer=1 filter=215 channel=26
    -76, -32, 14, -30, -54, 20, -24, -49, 12,
    -- layer=1 filter=215 channel=27
    -13, 7, 10, -11, -10, 11, 8, 13, 14,
    -- layer=1 filter=215 channel=28
    8, 42, 6, 13, 45, 18, 6, 41, 27,
    -- layer=1 filter=215 channel=29
    -29, 0, 11, -34, -17, 6, -18, -4, -1,
    -- layer=1 filter=215 channel=30
    13, -20, -35, -50, 23, 27, 7, 1, 0,
    -- layer=1 filter=215 channel=31
    -15, 9, -38, -18, 7, -7, 6, -23, -34,
    -- layer=1 filter=215 channel=32
    -65, -64, 10, -51, -112, 16, -28, -54, -13,
    -- layer=1 filter=215 channel=33
    30, 10, -15, 32, 6, -1, 20, 10, 5,
    -- layer=1 filter=215 channel=34
    94, 35, 6, 78, 43, 1, 40, -18, 7,
    -- layer=1 filter=215 channel=35
    -7, -12, 4, -17, -23, -9, -9, -14, -19,
    -- layer=1 filter=215 channel=36
    -9, 33, 18, -25, 37, 29, -12, 25, 43,
    -- layer=1 filter=215 channel=37
    -5, 20, -4, 5, -9, 8, 5, 27, 12,
    -- layer=1 filter=215 channel=38
    16, -8, -19, 7, -25, -19, 10, -35, -26,
    -- layer=1 filter=215 channel=39
    -21, 3, 25, 6, 21, 0, -2, -1, 0,
    -- layer=1 filter=215 channel=40
    -9, -14, -60, -7, 3, -32, -1, -3, -38,
    -- layer=1 filter=215 channel=41
    -19, -75, -14, -37, -78, 4, 2, -11, 0,
    -- layer=1 filter=215 channel=42
    1, -10, -22, -16, 10, -24, -28, -8, -28,
    -- layer=1 filter=215 channel=43
    -13, 24, 33, 18, -4, 15, 3, 28, -6,
    -- layer=1 filter=215 channel=44
    -104, -39, 41, -42, -69, 43, -39, -50, 19,
    -- layer=1 filter=215 channel=45
    -10, -5, 5, -9, -40, 21, -11, -28, -22,
    -- layer=1 filter=215 channel=46
    -13, -60, -8, -40, -4, -3, 21, 0, 29,
    -- layer=1 filter=215 channel=47
    -10, -31, 34, -10, -13, 5, -14, -16, -37,
    -- layer=1 filter=215 channel=48
    9, -7, -14, 0, -7, -22, 3, -22, -7,
    -- layer=1 filter=215 channel=49
    20, -12, -30, 27, -11, -23, 33, -18, -28,
    -- layer=1 filter=215 channel=50
    -2, -13, -36, -4, 7, 8, 7, -19, 7,
    -- layer=1 filter=215 channel=51
    22, 5, 19, 7, -8, -7, 2, -12, -18,
    -- layer=1 filter=215 channel=52
    -8, -25, -26, 10, 18, 34, 10, -4, -11,
    -- layer=1 filter=215 channel=53
    6, 0, -8, -12, -2, -15, -5, -17, -11,
    -- layer=1 filter=215 channel=54
    -14, 9, 14, -15, 25, -14, -4, 49, 17,
    -- layer=1 filter=215 channel=55
    -11, -1, 8, 5, 1, 7, -2, 5, 12,
    -- layer=1 filter=215 channel=56
    7, 7, 8, -2, -3, -10, -1, 0, -6,
    -- layer=1 filter=215 channel=57
    13, 42, 17, 6, 44, 11, 3, 26, 26,
    -- layer=1 filter=215 channel=58
    2, -8, 29, -13, 19, 17, -28, 29, 33,
    -- layer=1 filter=215 channel=59
    5, -1, 13, 15, -2, -13, 12, -9, 5,
    -- layer=1 filter=215 channel=60
    18, 15, 20, 3, 4, 19, 3, 20, 18,
    -- layer=1 filter=215 channel=61
    -3, 8, -6, -2, -1, 9, -4, 7, -8,
    -- layer=1 filter=215 channel=62
    -26, 5, 19, -11, -17, 15, -11, 13, -18,
    -- layer=1 filter=215 channel=63
    4, -3, 5, -22, 26, 26, -1, 28, 18,
    -- layer=1 filter=215 channel=64
    17, 8, 23, 7, -4, -2, -4, -4, -4,
    -- layer=1 filter=215 channel=65
    1, -20, 0, 1, -19, -18, -13, -11, -11,
    -- layer=1 filter=215 channel=66
    -5, 24, 19, -10, 10, 17, -1, 11, 23,
    -- layer=1 filter=215 channel=67
    -11, -10, -3, -12, -89, -76, 14, -86, -74,
    -- layer=1 filter=215 channel=68
    -106, -1, 18, -67, -69, 32, -53, -28, 25,
    -- layer=1 filter=215 channel=69
    -28, 0, 22, -12, -11, 7, -24, -7, -20,
    -- layer=1 filter=215 channel=70
    30, 26, 6, 76, -21, -47, 51, -29, -71,
    -- layer=1 filter=215 channel=71
    -13, -6, -14, -8, -26, -10, -2, 7, 2,
    -- layer=1 filter=215 channel=72
    15, -55, -11, -47, -28, -5, -4, -8, 7,
    -- layer=1 filter=215 channel=73
    -7, 6, 11, 8, 7, -4, 11, 9, 7,
    -- layer=1 filter=215 channel=74
    -50, 0, -28, -72, -36, 10, -39, -12, -6,
    -- layer=1 filter=215 channel=75
    37, 21, 27, 6, 42, 44, 14, 23, 3,
    -- layer=1 filter=215 channel=76
    -31, -19, 0, -37, -14, 22, -12, -13, -5,
    -- layer=1 filter=215 channel=77
    -2, -3, -23, 5, -16, -13, 27, -6, -5,
    -- layer=1 filter=215 channel=78
    0, 21, -3, -23, 8, 7, -5, 9, 16,
    -- layer=1 filter=215 channel=79
    -16, -5, 3, -2, -14, -4, -13, -3, -21,
    -- layer=1 filter=215 channel=80
    -2, -4, 0, -1, 2, 5, -4, -7, -7,
    -- layer=1 filter=215 channel=81
    9, -11, -8, 5, -6, -14, 17, 16, 3,
    -- layer=1 filter=215 channel=82
    15, -29, -10, 16, -30, -28, 21, -36, -40,
    -- layer=1 filter=215 channel=83
    -34, 0, 39, -1, -22, 31, -14, -22, 4,
    -- layer=1 filter=215 channel=84
    -31, -28, -32, -62, -26, 0, 0, -4, -1,
    -- layer=1 filter=215 channel=85
    10, -41, 25, -32, -2, -5, -36, 4, 3,
    -- layer=1 filter=215 channel=86
    -24, 10, 25, -20, 17, 14, -28, 6, 16,
    -- layer=1 filter=215 channel=87
    11, -55, -43, -46, -57, -25, 33, 18, -16,
    -- layer=1 filter=215 channel=88
    1, -15, -2, 23, -9, -12, 22, 7, -15,
    -- layer=1 filter=215 channel=89
    -2, -36, -23, 11, -43, -21, 4, -9, -43,
    -- layer=1 filter=215 channel=90
    -78, 5, 11, -44, -31, 33, -32, -62, 31,
    -- layer=1 filter=215 channel=91
    18, 2, -23, 14, -3, -33, 16, -19, -23,
    -- layer=1 filter=215 channel=92
    -34, -20, -5, 10, -68, 23, -53, -66, -56,
    -- layer=1 filter=215 channel=93
    -1, -5, 8, -10, -6, 2, -20, -10, 3,
    -- layer=1 filter=215 channel=94
    0, 22, 10, -9, 39, 25, -17, 18, 12,
    -- layer=1 filter=215 channel=95
    -15, -13, -18, -29, 5, 39, -2, 18, -12,
    -- layer=1 filter=215 channel=96
    9, 0, -8, 3, 17, 4, 8, 21, 13,
    -- layer=1 filter=215 channel=97
    -13, 13, 22, -4, 6, 13, -4, -9, 17,
    -- layer=1 filter=215 channel=98
    -3, 20, 21, 7, -5, 3, -22, -1, -18,
    -- layer=1 filter=215 channel=99
    -40, 58, -14, -62, 27, 39, -34, 24, 65,
    -- layer=1 filter=215 channel=100
    -7, -13, 3, -32, -7, -1, -4, 2, 1,
    -- layer=1 filter=215 channel=101
    -6, -9, -14, 10, -27, -22, 0, -22, -36,
    -- layer=1 filter=215 channel=102
    -3, 13, 15, -17, 10, 10, -19, 0, 1,
    -- layer=1 filter=215 channel=103
    15, 19, 27, -16, 0, 4, 1, 12, 12,
    -- layer=1 filter=215 channel=104
    -15, -27, 44, -50, -26, 30, -28, 4, 32,
    -- layer=1 filter=215 channel=105
    -10, 23, 27, -11, 16, 20, -22, 2, 20,
    -- layer=1 filter=215 channel=106
    -22, -30, -9, -7, -91, -14, -2, -41, -29,
    -- layer=1 filter=215 channel=107
    12, 2, -3, 0, 4, 13, 13, 12, 20,
    -- layer=1 filter=215 channel=108
    -90, -73, 18, -27, -78, 43, -39, -88, 0,
    -- layer=1 filter=215 channel=109
    3, 8, 4, -3, -3, -11, 3, 0, -5,
    -- layer=1 filter=215 channel=110
    -5, 20, 19, 6, 3, 1, -13, 11, 9,
    -- layer=1 filter=215 channel=111
    -10, 19, -9, -39, 19, 33, -1, 29, 8,
    -- layer=1 filter=215 channel=112
    -3, -10, -7, -10, 8, 18, -1, -4, -22,
    -- layer=1 filter=215 channel=113
    21, -7, -55, 19, 10, -70, -7, -27, -58,
    -- layer=1 filter=215 channel=114
    -7, 6, 31, 14, 19, 19, 17, 36, 11,
    -- layer=1 filter=215 channel=115
    -1, 36, 18, -18, 18, 24, -15, 14, 9,
    -- layer=1 filter=215 channel=116
    5, -10, 4, -4, 9, 1, 4, 2, -10,
    -- layer=1 filter=215 channel=117
    -6, 33, 22, -38, 19, 32, 21, 7, 13,
    -- layer=1 filter=215 channel=118
    -27, -19, -14, -62, -40, 19, -8, -2, 3,
    -- layer=1 filter=215 channel=119
    -77, -41, 12, -63, -68, 16, -37, -59, 13,
    -- layer=1 filter=215 channel=120
    31, -9, -11, 19, -14, -40, 19, -9, -13,
    -- layer=1 filter=215 channel=121
    -5, -22, -26, -7, 4, 9, 23, 24, 11,
    -- layer=1 filter=215 channel=122
    0, 1, 2, 8, -7, 0, -2, 2, 5,
    -- layer=1 filter=215 channel=123
    11, -2, 0, -11, 5, 11, -4, 17, 10,
    -- layer=1 filter=215 channel=124
    -8, -14, -10, 5, -2, 4, 3, -8, -3,
    -- layer=1 filter=215 channel=125
    24, 32, -27, 39, -33, -64, 54, -23, -56,
    -- layer=1 filter=215 channel=126
    1, 33, 15, 30, -6, 1, -8, -28, -35,
    -- layer=1 filter=215 channel=127
    -9, -11, -21, -33, 14, 31, 0, 18, -7,
    -- layer=1 filter=216 channel=0
    -5, -1, 0, -14, -11, -35, -19, -31, -10,
    -- layer=1 filter=216 channel=1
    -3, -15, -1, 6, 11, -2, -14, 13, 1,
    -- layer=1 filter=216 channel=2
    -16, -20, 6, 0, 11, 10, 49, 41, 49,
    -- layer=1 filter=216 channel=3
    6, 8, -1, -2, 5, -7, 0, -8, -1,
    -- layer=1 filter=216 channel=4
    -3, -7, 2, 4, 18, -2, 1, 0, 3,
    -- layer=1 filter=216 channel=5
    -18, -25, 0, 2, -6, 0, -9, 9, -4,
    -- layer=1 filter=216 channel=6
    74, 40, 12, -15, -18, -13, 10, 0, -14,
    -- layer=1 filter=216 channel=7
    26, -7, 5, 50, 14, 8, -7, -21, 14,
    -- layer=1 filter=216 channel=8
    -30, -34, -21, -6, -27, -11, -6, 18, 9,
    -- layer=1 filter=216 channel=9
    9, 60, 49, 63, 67, 100, 98, 116, 94,
    -- layer=1 filter=216 channel=10
    29, 17, 13, 31, 22, 28, -21, -25, 5,
    -- layer=1 filter=216 channel=11
    3, 3, 2, 0, -8, 2, -13, -1, -17,
    -- layer=1 filter=216 channel=12
    35, 18, 11, 19, 37, 33, 64, 81, 89,
    -- layer=1 filter=216 channel=13
    -2, 4, -5, -14, -37, -3, -6, -8, -5,
    -- layer=1 filter=216 channel=14
    13, -5, -6, 59, 51, 26, 41, 50, 22,
    -- layer=1 filter=216 channel=15
    -33, -32, -52, -20, -20, -25, 7, 8, -26,
    -- layer=1 filter=216 channel=16
    -30, -23, -6, -14, -15, 2, 16, 17, 10,
    -- layer=1 filter=216 channel=17
    -29, -25, -34, -37, -46, -42, -31, -27, -23,
    -- layer=1 filter=216 channel=18
    4, -22, -16, 0, 12, 2, 26, 24, 8,
    -- layer=1 filter=216 channel=19
    44, 72, 38, 57, 67, 83, 79, 72, 85,
    -- layer=1 filter=216 channel=20
    -8, -21, -9, -37, -46, -18, -35, -14, -13,
    -- layer=1 filter=216 channel=21
    43, 13, 13, 22, -4, -11, -17, -9, -8,
    -- layer=1 filter=216 channel=22
    10, -6, -3, -21, -33, -23, -30, -4, -6,
    -- layer=1 filter=216 channel=23
    61, 68, 47, 34, 45, 20, -24, -29, -47,
    -- layer=1 filter=216 channel=24
    8, 35, 3, 1, 17, 29, 12, 3, -7,
    -- layer=1 filter=216 channel=25
    34, 37, 27, 38, 38, 40, 4, 5, 39,
    -- layer=1 filter=216 channel=26
    -16, 13, 2, 0, 11, 12, 10, -11, -6,
    -- layer=1 filter=216 channel=27
    20, 8, 19, -9, -10, 8, -14, -16, -3,
    -- layer=1 filter=216 channel=28
    23, 6, 25, 22, 15, 14, 1, 10, 24,
    -- layer=1 filter=216 channel=29
    28, 12, 40, 33, 18, 24, 12, 2, 13,
    -- layer=1 filter=216 channel=30
    0, 0, -23, 2, 4, 20, 40, 58, 10,
    -- layer=1 filter=216 channel=31
    0, -39, -46, -11, -31, -42, -4, -20, -21,
    -- layer=1 filter=216 channel=32
    -9, 22, 10, 17, 40, 53, 11, 17, -17,
    -- layer=1 filter=216 channel=33
    25, 7, 23, -19, -16, -14, -17, -17, -20,
    -- layer=1 filter=216 channel=34
    63, 19, -7, -1, -21, -34, -38, -30, -13,
    -- layer=1 filter=216 channel=35
    -11, -18, -27, -7, -31, -20, -2, -16, -25,
    -- layer=1 filter=216 channel=36
    -2, 9, 17, -1, -15, 8, -13, -23, -13,
    -- layer=1 filter=216 channel=37
    -4, 3, 2, 22, 14, 18, 6, 8, 16,
    -- layer=1 filter=216 channel=38
    11, -7, -17, -20, -27, -12, -18, -19, -20,
    -- layer=1 filter=216 channel=39
    2, -20, -33, -14, -29, -19, -18, -21, -8,
    -- layer=1 filter=216 channel=40
    -16, -24, -42, -2, -5, -26, -2, 1, -29,
    -- layer=1 filter=216 channel=41
    -17, 32, 6, 31, 47, 71, 34, 60, 14,
    -- layer=1 filter=216 channel=42
    -18, -17, -3, 17, 12, 18, 55, 49, 54,
    -- layer=1 filter=216 channel=43
    0, -5, -2, -7, 9, 1, -4, 15, 35,
    -- layer=1 filter=216 channel=44
    3, 28, 22, 35, 25, 39, -9, -7, -27,
    -- layer=1 filter=216 channel=45
    9, 8, 11, 14, -8, 0, 10, 4, -11,
    -- layer=1 filter=216 channel=46
    43, 10, -13, 21, 20, 11, 74, 56, 53,
    -- layer=1 filter=216 channel=47
    4, 59, 24, 36, 26, 2, -35, -24, -60,
    -- layer=1 filter=216 channel=48
    17, 14, -4, 5, 0, -10, -17, -24, -30,
    -- layer=1 filter=216 channel=49
    35, 45, 27, 31, 16, 0, -2, 17, -21,
    -- layer=1 filter=216 channel=50
    10, -2, 1, 16, -11, 12, -1, 2, -9,
    -- layer=1 filter=216 channel=51
    27, 5, -15, -8, -3, -2, -19, -19, -24,
    -- layer=1 filter=216 channel=52
    7, 13, 3, 12, 27, 24, 3, 14, 0,
    -- layer=1 filter=216 channel=53
    -1, 11, -11, -4, 9, 0, -2, 7, 19,
    -- layer=1 filter=216 channel=54
    30, 40, 34, 24, 46, 48, 21, 1, 52,
    -- layer=1 filter=216 channel=55
    15, 27, 31, 2, 10, 3, -4, -12, -16,
    -- layer=1 filter=216 channel=56
    5, -7, 6, 10, 11, -3, 7, -3, 2,
    -- layer=1 filter=216 channel=57
    25, -7, 0, 3, 1, 12, -48, -41, -3,
    -- layer=1 filter=216 channel=58
    73, 63, 38, 65, 48, 50, -32, -36, -19,
    -- layer=1 filter=216 channel=59
    -9, 24, -31, -17, -29, -11, 21, 15, 2,
    -- layer=1 filter=216 channel=60
    -6, 14, -1, 26, 27, 4, -26, 6, -2,
    -- layer=1 filter=216 channel=61
    -13, 13, -7, 10, 4, 8, -1, 4, 5,
    -- layer=1 filter=216 channel=62
    0, -6, -13, 0, -1, 18, 5, 16, 10,
    -- layer=1 filter=216 channel=63
    5, 0, 13, -18, 0, 7, -15, -13, -17,
    -- layer=1 filter=216 channel=64
    14, -4, 7, 9, 14, -1, -15, 17, 0,
    -- layer=1 filter=216 channel=65
    9, 8, 1, -3, -18, -23, -23, -22, -16,
    -- layer=1 filter=216 channel=66
    0, 7, 18, -1, -13, -21, -28, -23, -16,
    -- layer=1 filter=216 channel=67
    118, 95, 81, 51, 56, 16, 58, 61, 30,
    -- layer=1 filter=216 channel=68
    3, 35, 11, 26, 20, 45, 1, -21, -13,
    -- layer=1 filter=216 channel=69
    -5, 4, -10, 2, 8, 1, 14, 21, -6,
    -- layer=1 filter=216 channel=70
    60, 22, 19, 42, 13, -29, 6, -8, -31,
    -- layer=1 filter=216 channel=71
    27, 19, 15, -4, 0, -6, -2, -22, -4,
    -- layer=1 filter=216 channel=72
    17, 20, -2, 33, 19, 44, 69, 60, 46,
    -- layer=1 filter=216 channel=73
    -2, -3, 3, 7, 9, 7, 6, -13, -5,
    -- layer=1 filter=216 channel=74
    7, 8, -3, 7, 16, 31, -19, 22, 23,
    -- layer=1 filter=216 channel=75
    23, 7, 4, 31, 51, 8, 64, 68, 48,
    -- layer=1 filter=216 channel=76
    -8, 3, -14, -5, -3, 32, -13, 1, -1,
    -- layer=1 filter=216 channel=77
    19, 32, 15, 1, -9, -11, -14, -30, -12,
    -- layer=1 filter=216 channel=78
    15, 29, -2, 1, 29, 13, 3, -11, -8,
    -- layer=1 filter=216 channel=79
    -20, -5, -7, -10, -1, -4, 8, 5, 14,
    -- layer=1 filter=216 channel=80
    2, 6, 4, -1, -18, -16, 7, 12, 12,
    -- layer=1 filter=216 channel=81
    13, 14, -1, -12, -5, -14, -12, -24, -9,
    -- layer=1 filter=216 channel=82
    18, 17, 2, 7, -5, -16, -17, -23, -32,
    -- layer=1 filter=216 channel=83
    -4, -13, -29, -5, -5, -23, -26, 7, -44,
    -- layer=1 filter=216 channel=84
    -3, 21, 9, 22, 42, 49, 48, 50, 42,
    -- layer=1 filter=216 channel=85
    42, 62, 40, 56, 50, 54, -2, -17, 1,
    -- layer=1 filter=216 channel=86
    -8, -8, 1, -10, -29, -9, -27, -28, -5,
    -- layer=1 filter=216 channel=87
    -18, 21, -5, 74, 27, 63, 33, 77, 50,
    -- layer=1 filter=216 channel=88
    25, 23, 18, 4, 21, 4, 8, 15, 7,
    -- layer=1 filter=216 channel=89
    15, 18, 8, 1, 6, -7, -20, -22, -39,
    -- layer=1 filter=216 channel=90
    -3, 8, 8, 22, -5, 26, 4, 0, -40,
    -- layer=1 filter=216 channel=91
    -8, -11, -38, -17, -21, -44, -36, -38, -38,
    -- layer=1 filter=216 channel=92
    -21, 14, 17, -2, 16, 47, -16, 37, -6,
    -- layer=1 filter=216 channel=93
    7, 5, 8, -11, 0, -16, -18, -10, -28,
    -- layer=1 filter=216 channel=94
    -26, -28, -21, -26, -21, -38, -27, -33, -23,
    -- layer=1 filter=216 channel=95
    13, 3, 9, 5, 30, 34, 37, 53, 10,
    -- layer=1 filter=216 channel=96
    4, 2, 8, 1, 11, 11, 0, -4, -24,
    -- layer=1 filter=216 channel=97
    -3, -5, 3, -22, -9, -24, -25, -18, -29,
    -- layer=1 filter=216 channel=98
    9, 14, -6, -1, -5, -8, 5, 6, 34,
    -- layer=1 filter=216 channel=99
    40, 47, 29, 51, 34, 19, -22, -26, -10,
    -- layer=1 filter=216 channel=100
    21, 8, 24, -15, -13, 0, -14, 3, -21,
    -- layer=1 filter=216 channel=101
    7, -26, -22, -12, -30, -21, -35, -31, -30,
    -- layer=1 filter=216 channel=102
    -30, -52, -31, -54, -43, -35, -38, -33, -46,
    -- layer=1 filter=216 channel=103
    12, 14, 3, -24, -2, 4, -8, 11, 6,
    -- layer=1 filter=216 channel=104
    -20, 10, 5, 25, 24, 9, 6, 14, -16,
    -- layer=1 filter=216 channel=105
    2, -11, -20, -20, -14, -9, -24, -33, -25,
    -- layer=1 filter=216 channel=106
    -11, 0, -1, -16, 5, -3, -25, -30, -39,
    -- layer=1 filter=216 channel=107
    -16, -11, -7, -6, -6, -8, -14, -9, -7,
    -- layer=1 filter=216 channel=108
    -21, 34, 2, 14, 12, 29, 8, 20, -27,
    -- layer=1 filter=216 channel=109
    -1, -4, 5, 7, 0, -4, -7, -3, -8,
    -- layer=1 filter=216 channel=110
    1, 4, -12, 10, 9, 6, -15, -10, -15,
    -- layer=1 filter=216 channel=111
    5, -17, -28, 10, 15, 13, 41, 40, 3,
    -- layer=1 filter=216 channel=112
    1, 4, 13, 11, 46, 10, 30, 40, 38,
    -- layer=1 filter=216 channel=113
    38, 0, -27, -12, -30, -47, -26, -45, -25,
    -- layer=1 filter=216 channel=114
    -20, -32, -32, 3, 8, -8, 3, 7, 2,
    -- layer=1 filter=216 channel=115
    0, -27, -27, -11, -6, -12, -30, -35, -6,
    -- layer=1 filter=216 channel=116
    -5, 9, 0, 2, -7, 0, -8, -2, -6,
    -- layer=1 filter=216 channel=117
    36, 3, -15, 75, 60, 35, 70, 63, 34,
    -- layer=1 filter=216 channel=118
    -2, 8, 4, 11, 13, 19, 30, 41, 31,
    -- layer=1 filter=216 channel=119
    -26, 21, 8, 18, 22, 46, 9, 7, -8,
    -- layer=1 filter=216 channel=120
    19, 29, -2, 7, -5, -2, -3, -5, 0,
    -- layer=1 filter=216 channel=121
    22, 11, 1, 16, 13, 6, 33, 49, 20,
    -- layer=1 filter=216 channel=122
    6, -2, -9, 8, 0, 5, 8, 4, -2,
    -- layer=1 filter=216 channel=123
    6, 18, 13, 1, 8, 0, -11, 21, -7,
    -- layer=1 filter=216 channel=124
    17, 5, -6, 3, 6, -13, 13, 22, -6,
    -- layer=1 filter=216 channel=125
    87, 50, 37, 77, 30, -2, -16, -40, -37,
    -- layer=1 filter=216 channel=126
    16, 22, -22, 10, -16, -23, 2, 0, -6,
    -- layer=1 filter=216 channel=127
    -12, -11, -1, 9, 10, 3, 40, 51, 13,
    -- layer=1 filter=217 channel=0
    -10, 0, -12, -14, 0, -9, 1, -16, -8,
    -- layer=1 filter=217 channel=1
    -15, 3, -17, 6, -5, -3, 1, -6, -13,
    -- layer=1 filter=217 channel=2
    -5, -4, -6, -3, -10, -9, 10, 0, -4,
    -- layer=1 filter=217 channel=3
    -7, 2, 9, -7, -8, 1, 9, 9, -1,
    -- layer=1 filter=217 channel=4
    1, -1, -3, 8, 0, 7, -5, -4, -3,
    -- layer=1 filter=217 channel=5
    -2, -1, -14, -16, -7, -14, -14, 2, -5,
    -- layer=1 filter=217 channel=6
    -5, 3, -2, 0, -3, -7, 1, -10, 10,
    -- layer=1 filter=217 channel=7
    -13, -4, -6, -1, 0, -7, -1, -11, -4,
    -- layer=1 filter=217 channel=8
    -5, -7, -9, 4, -9, 5, -17, -12, -9,
    -- layer=1 filter=217 channel=9
    0, -18, -7, 1, -1, 8, 7, -9, -4,
    -- layer=1 filter=217 channel=10
    0, -10, -17, -12, -11, -10, -9, -11, -4,
    -- layer=1 filter=217 channel=11
    -2, -9, 3, -11, 5, -6, -6, -2, 4,
    -- layer=1 filter=217 channel=12
    2, -10, 5, 7, 12, 3, -15, 0, -13,
    -- layer=1 filter=217 channel=13
    3, -6, -12, 0, -3, 0, 3, 3, 0,
    -- layer=1 filter=217 channel=14
    -4, -3, -14, 4, 3, -5, -5, 5, -7,
    -- layer=1 filter=217 channel=15
    2, -4, -6, -2, -16, -9, 1, 5, 1,
    -- layer=1 filter=217 channel=16
    -1, 0, -4, -4, 0, -9, -13, -2, -10,
    -- layer=1 filter=217 channel=17
    1, -10, -9, 0, -9, -5, 3, -10, -4,
    -- layer=1 filter=217 channel=18
    0, -13, -2, 4, -7, -11, -1, -8, 5,
    -- layer=1 filter=217 channel=19
    8, 11, -5, 0, -5, 5, 1, 6, 4,
    -- layer=1 filter=217 channel=20
    -7, 5, -7, 2, 4, 1, -9, -1, -11,
    -- layer=1 filter=217 channel=21
    -9, 5, 6, -1, -6, 0, 6, 3, -9,
    -- layer=1 filter=217 channel=22
    -6, -1, -9, 0, 9, -8, 2, 4, 4,
    -- layer=1 filter=217 channel=23
    -17, 0, 0, -12, -5, 2, -23, -13, 0,
    -- layer=1 filter=217 channel=24
    -3, -7, -1, -5, -1, 5, -1, -12, 1,
    -- layer=1 filter=217 channel=25
    -14, 5, -10, -2, -3, -13, -2, -13, 2,
    -- layer=1 filter=217 channel=26
    1, -14, 3, -15, 0, -9, -1, 5, 5,
    -- layer=1 filter=217 channel=27
    -10, 6, 2, -7, -1, -6, -10, 5, 2,
    -- layer=1 filter=217 channel=28
    -1, 0, -15, 0, 0, -14, 1, -4, 1,
    -- layer=1 filter=217 channel=29
    4, 0, -8, -14, -14, -5, 0, 2, -12,
    -- layer=1 filter=217 channel=30
    -12, -12, -1, -15, -2, -9, -5, 0, 5,
    -- layer=1 filter=217 channel=31
    -1, -6, 13, -3, 12, 9, -3, 3, -1,
    -- layer=1 filter=217 channel=32
    -4, 0, -1, -3, 1, 7, -17, -1, 5,
    -- layer=1 filter=217 channel=33
    9, 0, 0, -1, 11, 0, 3, -8, 5,
    -- layer=1 filter=217 channel=34
    -6, -7, 4, -2, 3, -6, -1, 7, 6,
    -- layer=1 filter=217 channel=35
    5, -9, -1, -6, -12, -1, 7, -2, -2,
    -- layer=1 filter=217 channel=36
    -5, -17, -3, -5, -3, -5, 2, -4, -12,
    -- layer=1 filter=217 channel=37
    0, 5, -6, 5, -15, -5, 3, -2, 8,
    -- layer=1 filter=217 channel=38
    -2, 3, -8, 0, -5, -9, -1, 5, 2,
    -- layer=1 filter=217 channel=39
    -10, 0, -12, -2, -13, 4, -8, -9, -14,
    -- layer=1 filter=217 channel=40
    6, -13, -11, 8, 9, 5, 5, 0, -7,
    -- layer=1 filter=217 channel=41
    -3, -15, -11, -3, -3, 5, -18, 3, 17,
    -- layer=1 filter=217 channel=42
    2, 5, -12, 5, -11, 0, -4, 3, 14,
    -- layer=1 filter=217 channel=43
    -14, 2, -8, -4, -4, 1, -2, -12, -2,
    -- layer=1 filter=217 channel=44
    -3, 0, -3, -15, -17, 2, -17, -7, -3,
    -- layer=1 filter=217 channel=45
    8, -10, 5, 7, -2, -5, -1, -4, -10,
    -- layer=1 filter=217 channel=46
    1, -6, -6, 8, -13, -18, 0, 10, 3,
    -- layer=1 filter=217 channel=47
    -1, -17, -10, -1, 7, 13, -12, 4, -4,
    -- layer=1 filter=217 channel=48
    1, 8, -11, -8, -6, 5, 1, 2, -8,
    -- layer=1 filter=217 channel=49
    -10, 5, 6, -6, 6, 7, -1, -1, -2,
    -- layer=1 filter=217 channel=50
    5, 1, 6, -6, 0, -2, 7, 0, 12,
    -- layer=1 filter=217 channel=51
    -4, -7, 4, 4, 6, 0, 6, -3, 9,
    -- layer=1 filter=217 channel=52
    -7, 10, 3, -9, 8, 0, 2, -4, -4,
    -- layer=1 filter=217 channel=53
    0, -1, -9, 7, -6, -6, -9, 2, 3,
    -- layer=1 filter=217 channel=54
    1, 6, -13, -7, -10, -20, -2, 5, 5,
    -- layer=1 filter=217 channel=55
    -10, -13, 6, 4, 0, 5, -7, 0, -2,
    -- layer=1 filter=217 channel=56
    0, 4, 3, -8, 9, 4, 7, -5, 9,
    -- layer=1 filter=217 channel=57
    -8, -2, -2, -2, -11, -8, -2, -9, -7,
    -- layer=1 filter=217 channel=58
    -11, -2, 3, -6, 1, -11, 2, -6, -3,
    -- layer=1 filter=217 channel=59
    -2, 7, -9, 0, 1, 0, -18, -15, 1,
    -- layer=1 filter=217 channel=60
    -6, -6, -9, 0, -6, -9, 9, -6, 9,
    -- layer=1 filter=217 channel=61
    0, -9, -4, 8, -2, -4, 0, -8, 0,
    -- layer=1 filter=217 channel=62
    5, 7, -17, 6, 1, 2, -4, -7, 7,
    -- layer=1 filter=217 channel=63
    0, -9, -4, 1, -6, 6, -9, -8, -11,
    -- layer=1 filter=217 channel=64
    -2, -6, 7, 2, 8, 5, 5, -9, -10,
    -- layer=1 filter=217 channel=65
    -10, -1, 8, 4, -5, 6, 5, 0, -9,
    -- layer=1 filter=217 channel=66
    -16, -3, -8, 3, -4, -6, -16, -7, -17,
    -- layer=1 filter=217 channel=67
    9, -3, -1, 5, 0, -2, 0, 0, 5,
    -- layer=1 filter=217 channel=68
    0, -3, -11, -12, -13, 5, -10, 2, -9,
    -- layer=1 filter=217 channel=69
    -1, 1, -10, -5, 0, -2, -2, 7, 6,
    -- layer=1 filter=217 channel=70
    12, 3, 2, 7, 10, 1, -4, 3, 3,
    -- layer=1 filter=217 channel=71
    6, -6, 6, -10, -16, -1, -2, -3, 9,
    -- layer=1 filter=217 channel=72
    -10, -4, -4, -11, -11, -11, -6, -3, 0,
    -- layer=1 filter=217 channel=73
    3, -7, -5, 1, -11, 6, 3, 3, -4,
    -- layer=1 filter=217 channel=74
    -8, 0, 7, -8, 3, 6, -4, 5, -6,
    -- layer=1 filter=217 channel=75
    -11, -4, 5, 1, 2, -13, 5, 10, -4,
    -- layer=1 filter=217 channel=76
    0, -8, -11, -14, -8, 5, -11, -5, 4,
    -- layer=1 filter=217 channel=77
    -5, -9, -10, -5, -2, -5, -6, -3, 2,
    -- layer=1 filter=217 channel=78
    0, -13, -14, -16, -14, -3, -12, -13, -16,
    -- layer=1 filter=217 channel=79
    -8, -6, -11, -4, -7, 3, -2, 0, -7,
    -- layer=1 filter=217 channel=80
    -16, 5, -7, 9, -19, 11, -2, 9, 3,
    -- layer=1 filter=217 channel=81
    -11, -4, -11, 3, 6, 1, -9, -1, 6,
    -- layer=1 filter=217 channel=82
    -12, -2, -9, 7, -9, -1, -11, -10, -7,
    -- layer=1 filter=217 channel=83
    3, -3, -15, -10, -7, -3, -18, -10, -14,
    -- layer=1 filter=217 channel=84
    5, -11, -8, -4, 1, -2, -4, 0, 2,
    -- layer=1 filter=217 channel=85
    6, 8, -2, 5, -13, -11, 0, -3, -4,
    -- layer=1 filter=217 channel=86
    -5, 2, -6, 0, -11, -11, -16, -9, -9,
    -- layer=1 filter=217 channel=87
    -5, 0, -6, -3, 6, 9, -15, -8, -7,
    -- layer=1 filter=217 channel=88
    -8, -8, 6, 8, -3, 7, 5, 4, -6,
    -- layer=1 filter=217 channel=89
    -11, -13, 2, 2, -7, -11, 3, 2, -2,
    -- layer=1 filter=217 channel=90
    -2, -1, -5, -6, -4, -5, -17, -1, 6,
    -- layer=1 filter=217 channel=91
    -1, 7, 7, 2, -7, -9, 4, 0, -2,
    -- layer=1 filter=217 channel=92
    -3, 2, -7, -23, -7, 4, -14, -1, 0,
    -- layer=1 filter=217 channel=93
    -11, 10, 0, 5, 0, -7, 5, -7, 5,
    -- layer=1 filter=217 channel=94
    -4, -12, -5, -11, -6, -12, -2, -13, -15,
    -- layer=1 filter=217 channel=95
    4, -12, -9, 0, -10, 6, -6, -7, -4,
    -- layer=1 filter=217 channel=96
    -13, -8, 8, -3, -9, 4, -10, 4, -7,
    -- layer=1 filter=217 channel=97
    -11, -3, -6, -12, 0, -9, 2, -8, -5,
    -- layer=1 filter=217 channel=98
    4, -1, -5, -9, -1, -12, 2, -2, -8,
    -- layer=1 filter=217 channel=99
    -11, -4, -9, -11, -2, 0, -5, 0, 3,
    -- layer=1 filter=217 channel=100
    -9, -6, -5, 2, -1, -3, -4, 0, 5,
    -- layer=1 filter=217 channel=101
    1, -5, -5, -9, -1, 8, 3, -6, 4,
    -- layer=1 filter=217 channel=102
    -10, 3, -13, -15, -13, -13, -2, -7, -7,
    -- layer=1 filter=217 channel=103
    4, -1, 2, -5, 4, 9, 1, 1, 2,
    -- layer=1 filter=217 channel=104
    -4, -10, 4, -12, 5, 0, 0, -5, 2,
    -- layer=1 filter=217 channel=105
    -17, 3, -11, 1, 2, -8, -7, -8, 3,
    -- layer=1 filter=217 channel=106
    -11, 1, 6, 0, 0, 3, 0, -7, -5,
    -- layer=1 filter=217 channel=107
    6, -5, 7, -8, 8, 6, -9, 6, 4,
    -- layer=1 filter=217 channel=108
    -6, -8, -15, -18, -2, 4, 0, 0, -2,
    -- layer=1 filter=217 channel=109
    -1, 6, 5, -10, 7, -6, 6, -3, 4,
    -- layer=1 filter=217 channel=110
    -20, -13, 2, -17, -11, 1, -3, 8, -11,
    -- layer=1 filter=217 channel=111
    -2, -5, -2, 0, 0, 0, -9, 5, -5,
    -- layer=1 filter=217 channel=112
    -5, -8, -8, 6, 11, -7, -6, -12, -9,
    -- layer=1 filter=217 channel=113
    8, 6, -9, 10, 8, 8, 0, -6, 18,
    -- layer=1 filter=217 channel=114
    -15, -13, -18, -1, -4, -12, -1, -11, 1,
    -- layer=1 filter=217 channel=115
    -16, 5, -14, -15, -7, -8, -4, -18, -12,
    -- layer=1 filter=217 channel=116
    0, -4, -2, -3, -8, 7, -10, 8, 4,
    -- layer=1 filter=217 channel=117
    -4, -11, -13, -7, 11, -6, -11, 3, -7,
    -- layer=1 filter=217 channel=118
    -1, -13, 0, 0, 0, 8, -6, 4, 5,
    -- layer=1 filter=217 channel=119
    -17, -13, -12, -9, -12, -3, -2, -16, 0,
    -- layer=1 filter=217 channel=120
    -8, -7, -10, -10, -4, -7, -2, -3, -6,
    -- layer=1 filter=217 channel=121
    -7, -10, 2, -11, -5, -2, 3, -2, -1,
    -- layer=1 filter=217 channel=122
    1, 0, 6, 0, 0, 2, -2, -4, -7,
    -- layer=1 filter=217 channel=123
    -12, -1, -3, -9, 0, -8, -5, -6, -1,
    -- layer=1 filter=217 channel=124
    -8, -3, 6, 6, 7, -1, 2, -2, -4,
    -- layer=1 filter=217 channel=125
    4, 13, 2, 12, -1, 9, 7, -1, 6,
    -- layer=1 filter=217 channel=126
    -13, 2, -11, 10, -4, -9, 2, 0, -8,
    -- layer=1 filter=217 channel=127
    3, -16, -1, -7, 5, -8, 0, 5, 2,
    -- layer=1 filter=218 channel=0
    26, 20, -2, -11, -9, -24, -22, -20, -9,
    -- layer=1 filter=218 channel=1
    27, 5, -30, 5, -9, 9, -15, 13, -3,
    -- layer=1 filter=218 channel=2
    3, -5, 0, -29, -37, -1, -33, -17, -3,
    -- layer=1 filter=218 channel=3
    7, 0, -5, -14, -12, -14, -6, 11, -8,
    -- layer=1 filter=218 channel=4
    -6, 6, 3, -1, -2, 3, 3, 9, -2,
    -- layer=1 filter=218 channel=5
    17, -17, -30, -12, -4, 18, -21, -14, -1,
    -- layer=1 filter=218 channel=6
    -52, -81, -39, -48, -36, -14, 5, -6, 14,
    -- layer=1 filter=218 channel=7
    -7, -66, -70, -111, -134, -65, -70, -57, -17,
    -- layer=1 filter=218 channel=8
    15, -23, -26, 29, 5, 36, 1, 22, 13,
    -- layer=1 filter=218 channel=9
    -11, -26, 62, -8, -42, -5, 4, -4, -13,
    -- layer=1 filter=218 channel=10
    -19, -108, -80, -119, -118, -63, -52, -43, -24,
    -- layer=1 filter=218 channel=11
    34, 41, 35, 16, 12, -8, -3, -28, -33,
    -- layer=1 filter=218 channel=12
    -71, -41, -57, -56, -59, -7, 3, 23, -48,
    -- layer=1 filter=218 channel=13
    -14, -41, -17, 0, 3, -1, 28, 17, 29,
    -- layer=1 filter=218 channel=14
    -71, -21, -45, -69, -85, -93, -73, -72, -53,
    -- layer=1 filter=218 channel=15
    3, -38, -85, -43, -5, 10, -17, -28, 6,
    -- layer=1 filter=218 channel=16
    11, -15, -36, 4, 1, 38, -4, 1, 1,
    -- layer=1 filter=218 channel=17
    16, -1, -14, 11, -6, -34, 9, -2, -15,
    -- layer=1 filter=218 channel=18
    11, 27, 33, 8, 7, 7, 44, -39, -48,
    -- layer=1 filter=218 channel=19
    55, 51, 56, 53, 33, 60, 45, 37, -49,
    -- layer=1 filter=218 channel=20
    -6, -32, -24, 8, -6, 12, 20, 40, 29,
    -- layer=1 filter=218 channel=21
    -22, -27, -10, -6, 8, 6, 23, 27, 51,
    -- layer=1 filter=218 channel=22
    -20, -20, -25, 8, 23, 21, 0, 33, 35,
    -- layer=1 filter=218 channel=23
    9, -15, -50, -65, -58, -89, -19, -39, -72,
    -- layer=1 filter=218 channel=24
    7, 0, 15, 13, 16, 21, 7, 32, 7,
    -- layer=1 filter=218 channel=25
    23, -40, -41, -37, -3, 13, 0, 1, -2,
    -- layer=1 filter=218 channel=26
    5, -1, 27, 30, 20, 27, 20, 0, -20,
    -- layer=1 filter=218 channel=27
    20, 46, 15, 3, -6, 0, -7, 23, 23,
    -- layer=1 filter=218 channel=28
    23, -37, -74, -20, -80, -25, -34, -17, 0,
    -- layer=1 filter=218 channel=29
    11, 6, -9, -26, -59, -44, -35, -20, -12,
    -- layer=1 filter=218 channel=30
    22, 14, 52, 13, 18, 39, 90, 17, -61,
    -- layer=1 filter=218 channel=31
    -40, -46, -25, -27, -13, -9, 16, 6, -11,
    -- layer=1 filter=218 channel=32
    32, -10, 48, 22, -2, -1, 30, -11, -52,
    -- layer=1 filter=218 channel=33
    0, 7, -9, -3, 2, -2, 8, 18, 13,
    -- layer=1 filter=218 channel=34
    -11, -46, 24, -22, -17, 13, 36, 49, 44,
    -- layer=1 filter=218 channel=35
    -12, -13, -9, -10, -9, 0, 4, -6, -9,
    -- layer=1 filter=218 channel=36
    36, 32, 38, 6, 11, -22, -15, -22, -30,
    -- layer=1 filter=218 channel=37
    28, -10, -36, -9, -15, 29, 0, 0, -1,
    -- layer=1 filter=218 channel=38
    -17, -24, -3, -12, 11, 18, 30, 30, 26,
    -- layer=1 filter=218 channel=39
    16, 0, -7, 0, -8, -4, 0, -1, -3,
    -- layer=1 filter=218 channel=40
    -40, -21, -6, -15, -6, -10, 40, -5, -3,
    -- layer=1 filter=218 channel=41
    56, 4, 37, 24, -26, -3, 50, -5, -87,
    -- layer=1 filter=218 channel=42
    -7, -14, -14, -27, -33, -20, -34, -44, -14,
    -- layer=1 filter=218 channel=43
    6, -23, -48, 17, 10, 31, 15, 7, 18,
    -- layer=1 filter=218 channel=44
    4, -5, 26, 40, 19, -21, -8, -37, -34,
    -- layer=1 filter=218 channel=45
    -13, -30, -29, -2, -7, 22, -5, 26, 26,
    -- layer=1 filter=218 channel=46
    13, 5, -12, 8, -23, -43, -22, -45, -63,
    -- layer=1 filter=218 channel=47
    18, -33, -41, -65, -57, -36, 19, -5, -32,
    -- layer=1 filter=218 channel=48
    -17, -15, -17, -18, -3, 7, 19, 9, 30,
    -- layer=1 filter=218 channel=49
    -3, -38, -9, -38, -24, 16, 26, 32, 46,
    -- layer=1 filter=218 channel=50
    -18, -18, 17, 2, 6, -8, 27, 17, -3,
    -- layer=1 filter=218 channel=51
    -31, -32, -36, -44, -19, 9, 7, 35, 14,
    -- layer=1 filter=218 channel=52
    -7, 18, 24, 11, -6, 0, 7, 29, 39,
    -- layer=1 filter=218 channel=53
    -1, -5, 0, -15, 11, -2, -3, -16, 7,
    -- layer=1 filter=218 channel=54
    47, -4, -9, -27, 8, 21, -3, -2, -9,
    -- layer=1 filter=218 channel=55
    25, 27, 24, -1, -14, -2, -27, -23, -11,
    -- layer=1 filter=218 channel=56
    -8, -7, 7, -8, -4, -4, 0, 1, -5,
    -- layer=1 filter=218 channel=57
    -23, -93, -93, -97, -84, -42, -21, -14, -11,
    -- layer=1 filter=218 channel=58
    -41, -108, -92, -114, -105, -65, -17, -39, -63,
    -- layer=1 filter=218 channel=59
    0, -2, -6, 1, 0, -7, -9, -2, 3,
    -- layer=1 filter=218 channel=60
    15, -3, -3, -1, 9, 7, 0, -9, -1,
    -- layer=1 filter=218 channel=61
    -1, 3, 3, -6, 3, -2, -3, 1, -4,
    -- layer=1 filter=218 channel=62
    43, -10, -23, 14, 18, 42, 6, 11, 18,
    -- layer=1 filter=218 channel=63
    44, 47, 37, 4, 1, -5, -10, -47, -49,
    -- layer=1 filter=218 channel=64
    -11, -13, -29, 5, 0, -3, -1, 17, 18,
    -- layer=1 filter=218 channel=65
    -18, -16, -10, 5, -4, 0, 7, 15, 15,
    -- layer=1 filter=218 channel=66
    32, 25, -2, 0, -26, -22, -25, -36, -26,
    -- layer=1 filter=218 channel=67
    -40, -39, -41, -45, -22, -3, -7, 21, 29,
    -- layer=1 filter=218 channel=68
    24, 16, 32, 33, 10, -2, -12, -24, -30,
    -- layer=1 filter=218 channel=69
    1, -14, -49, 14, -5, 14, -6, -2, -6,
    -- layer=1 filter=218 channel=70
    -69, -82, -64, -85, -77, 2, -10, 12, 12,
    -- layer=1 filter=218 channel=71
    -13, 2, -1, 5, -3, 10, 8, 4, 6,
    -- layer=1 filter=218 channel=72
    14, 14, 32, 64, 19, 34, 50, 3, -45,
    -- layer=1 filter=218 channel=73
    5, -2, 1, -4, -15, 1, -8, -10, -17,
    -- layer=1 filter=218 channel=74
    5, -2, 6, 7, 16, -26, 12, -46, -46,
    -- layer=1 filter=218 channel=75
    -47, -38, -14, -37, -26, -24, 8, -31, -38,
    -- layer=1 filter=218 channel=76
    9, 20, 24, 16, 12, -37, 21, -53, -72,
    -- layer=1 filter=218 channel=77
    -31, -17, -28, -11, -6, -2, 6, 19, 23,
    -- layer=1 filter=218 channel=78
    17, 7, 10, -14, -21, -24, -18, -21, 10,
    -- layer=1 filter=218 channel=79
    20, -6, -40, 14, 12, 29, 23, 9, 25,
    -- layer=1 filter=218 channel=80
    8, 3, -2, 4, 4, 5, -9, -2, -5,
    -- layer=1 filter=218 channel=81
    -30, -33, -32, -14, 5, 21, -11, 7, 28,
    -- layer=1 filter=218 channel=82
    -20, -25, -22, -5, 10, 8, 22, 41, 52,
    -- layer=1 filter=218 channel=83
    0, -33, -31, 16, -13, 1, 10, 0, 11,
    -- layer=1 filter=218 channel=84
    47, 59, 68, 51, 48, 24, 63, -35, -49,
    -- layer=1 filter=218 channel=85
    32, -36, -39, -32, -51, -63, -13, -16, -56,
    -- layer=1 filter=218 channel=86
    38, 45, 21, 6, -16, -16, -23, -33, -14,
    -- layer=1 filter=218 channel=87
    17, -33, 3, 48, -5, 11, -11, 22, -35,
    -- layer=1 filter=218 channel=88
    -31, -22, -21, -30, -10, 11, 8, 25, 30,
    -- layer=1 filter=218 channel=89
    -10, -2, 10, 11, 8, 11, 15, 9, 18,
    -- layer=1 filter=218 channel=90
    -17, -38, 0, 5, -20, -11, -22, -9, -23,
    -- layer=1 filter=218 channel=91
    -3, -25, -20, -11, 4, -5, 29, 17, 36,
    -- layer=1 filter=218 channel=92
    18, -75, -40, -33, -33, -26, -13, -28, -33,
    -- layer=1 filter=218 channel=93
    -7, -12, -17, 4, 12, 1, -2, 28, 22,
    -- layer=1 filter=218 channel=94
    29, 8, 10, 7, -28, -38, -10, -32, -43,
    -- layer=1 filter=218 channel=95
    43, 51, 65, 32, 55, 23, 76, -33, -51,
    -- layer=1 filter=218 channel=96
    7, 6, -7, -12, -22, -29, -16, -9, -4,
    -- layer=1 filter=218 channel=97
    12, 0, -7, 4, -5, -19, -10, -13, 1,
    -- layer=1 filter=218 channel=98
    15, -39, -26, 25, 22, 24, 3, 32, 31,
    -- layer=1 filter=218 channel=99
    -28, -46, -94, -84, -92, -100, -27, -44, -55,
    -- layer=1 filter=218 channel=100
    51, 49, 41, 7, 12, -21, 24, -11, -25,
    -- layer=1 filter=218 channel=101
    -1, -9, -11, -4, 6, -2, 22, 26, 32,
    -- layer=1 filter=218 channel=102
    23, 11, -4, -2, -26, -50, -5, -35, -24,
    -- layer=1 filter=218 channel=103
    23, 43, 42, 20, 5, 0, 11, 10, 7,
    -- layer=1 filter=218 channel=104
    19, 0, 7, 8, -7, -26, 17, 21, -43,
    -- layer=1 filter=218 channel=105
    28, 6, 1, 0, -24, -9, -8, -17, -15,
    -- layer=1 filter=218 channel=106
    -13, -4, 9, 4, 14, -8, 30, 14, 32,
    -- layer=1 filter=218 channel=107
    1, -4, 6, 5, 14, 16, 16, -1, 6,
    -- layer=1 filter=218 channel=108
    0, -27, 2, 31, -8, -18, 12, 7, -39,
    -- layer=1 filter=218 channel=109
    6, -8, 8, 0, -4, -5, -9, 0, -4,
    -- layer=1 filter=218 channel=110
    0, -2, 5, -6, -10, -1, -8, -2, -6,
    -- layer=1 filter=218 channel=111
    29, 16, 29, 19, 26, 19, 61, -33, -64,
    -- layer=1 filter=218 channel=112
    11, 17, 15, 10, 7, -14, 17, -38, 2,
    -- layer=1 filter=218 channel=113
    -19, -44, -40, -58, -49, -19, 8, -17, -19,
    -- layer=1 filter=218 channel=114
    -30, -6, -57, -11, -20, -3, -31, -26, -24,
    -- layer=1 filter=218 channel=115
    25, -4, -1, -20, -25, -20, -19, -22, -15,
    -- layer=1 filter=218 channel=116
    -1, 3, 4, 3, 1, -9, 0, 10, -4,
    -- layer=1 filter=218 channel=117
    1, 14, 14, 11, 0, -27, -11, -34, -8,
    -- layer=1 filter=218 channel=118
    31, 30, 40, 14, 27, 8, 56, -25, -42,
    -- layer=1 filter=218 channel=119
    13, 2, 30, 36, 4, -2, 28, -7, -26,
    -- layer=1 filter=218 channel=120
    -11, -34, -21, -40, -10, -3, 10, 24, 36,
    -- layer=1 filter=218 channel=121
    5, -8, 16, -2, -11, -11, 8, 0, -44,
    -- layer=1 filter=218 channel=122
    4, -4, -6, 0, 0, 0, 7, -5, 4,
    -- layer=1 filter=218 channel=123
    2, 21, 21, -2, -23, -5, 9, -21, -35,
    -- layer=1 filter=218 channel=124
    0, -5, -8, -18, -10, -7, -24, -25, -14,
    -- layer=1 filter=218 channel=125
    -76, -89, -103, -81, -90, -13, -17, 9, 0,
    -- layer=1 filter=218 channel=126
    -6, -36, -41, 43, 24, 50, 9, 28, 38,
    -- layer=1 filter=218 channel=127
    37, 36, 57, 28, 33, 33, 66, -17, -40,
    -- layer=1 filter=219 channel=0
    -12, 7, 2, -3, 5, 3, 0, -4, -3,
    -- layer=1 filter=219 channel=1
    4, -11, -4, 2, 7, -3, 7, 8, -8,
    -- layer=1 filter=219 channel=2
    -16, -2, 1, 6, -9, -15, -1, -14, -10,
    -- layer=1 filter=219 channel=3
    -7, -3, -9, -7, 6, -5, 6, 10, 0,
    -- layer=1 filter=219 channel=4
    3, -1, -10, 6, 5, -8, -3, -6, 5,
    -- layer=1 filter=219 channel=5
    2, 6, -4, -13, -1, -2, 2, 7, -8,
    -- layer=1 filter=219 channel=6
    4, 2, 6, -9, 8, -13, 7, 2, 0,
    -- layer=1 filter=219 channel=7
    -8, -4, -3, 1, -3, 4, -6, 6, 4,
    -- layer=1 filter=219 channel=8
    -4, 1, 0, 1, 1, -8, -2, -6, -6,
    -- layer=1 filter=219 channel=9
    -11, 6, 8, -2, -6, 2, -2, -7, -18,
    -- layer=1 filter=219 channel=10
    1, 5, -2, 6, 0, -2, 3, 7, -9,
    -- layer=1 filter=219 channel=11
    1, -2, 3, 4, -3, -4, -2, -11, 2,
    -- layer=1 filter=219 channel=12
    -1, -5, 6, 8, 7, -9, -6, -6, -2,
    -- layer=1 filter=219 channel=13
    2, 6, -4, -7, 5, 5, -2, 3, 2,
    -- layer=1 filter=219 channel=14
    6, 0, -2, 5, 4, 0, -2, 4, -5,
    -- layer=1 filter=219 channel=15
    -6, 11, -2, 6, 3, -4, -5, -5, -3,
    -- layer=1 filter=219 channel=16
    3, -8, 11, -11, -12, 11, -11, 6, 8,
    -- layer=1 filter=219 channel=17
    -11, -5, 0, 4, -2, 0, -9, -11, -10,
    -- layer=1 filter=219 channel=18
    -11, -11, -11, 0, -7, 2, 0, 11, 2,
    -- layer=1 filter=219 channel=19
    -7, -9, 7, 6, -8, -10, 6, 3, 5,
    -- layer=1 filter=219 channel=20
    3, -10, 0, 8, 2, -8, 0, 4, -8,
    -- layer=1 filter=219 channel=21
    -9, -11, -11, -14, 5, 3, 9, -11, -4,
    -- layer=1 filter=219 channel=22
    -5, 1, 7, -5, 1, 3, 0, 4, 3,
    -- layer=1 filter=219 channel=23
    0, 0, -10, -10, -3, 2, 8, -9, -2,
    -- layer=1 filter=219 channel=24
    -13, -9, -1, -9, 4, -14, -12, -9, -3,
    -- layer=1 filter=219 channel=25
    4, 5, 0, -5, -2, 3, -12, 0, -7,
    -- layer=1 filter=219 channel=26
    -13, -9, -6, 1, -4, 0, 9, 6, -13,
    -- layer=1 filter=219 channel=27
    -6, -1, -1, 3, 6, -2, 0, -7, -5,
    -- layer=1 filter=219 channel=28
    6, -9, -4, -10, 0, 2, 2, 0, -10,
    -- layer=1 filter=219 channel=29
    0, -5, 10, -4, -5, -3, 5, -2, -5,
    -- layer=1 filter=219 channel=30
    0, 0, -15, 0, -8, 3, 1, 7, -5,
    -- layer=1 filter=219 channel=31
    -8, -4, 0, 6, -9, -8, -6, 0, 5,
    -- layer=1 filter=219 channel=32
    -10, -9, 6, -3, -5, -8, -10, -2, 6,
    -- layer=1 filter=219 channel=33
    -3, -5, 6, 3, -7, 10, -3, -2, -1,
    -- layer=1 filter=219 channel=34
    -9, 3, -9, 5, 3, 4, 2, 0, -2,
    -- layer=1 filter=219 channel=35
    9, 1, 7, -5, 7, 4, -9, -7, 2,
    -- layer=1 filter=219 channel=36
    5, -6, -4, 0, -8, -1, 0, -10, -2,
    -- layer=1 filter=219 channel=37
    -3, -8, -5, 3, 2, -2, 0, 0, 3,
    -- layer=1 filter=219 channel=38
    -12, 0, -6, -13, 2, -6, 3, 0, 5,
    -- layer=1 filter=219 channel=39
    8, -7, -9, 8, 0, -5, 2, -6, -10,
    -- layer=1 filter=219 channel=40
    11, 7, -8, -3, 12, -5, -9, 1, -6,
    -- layer=1 filter=219 channel=41
    -4, 7, -9, -9, 0, -9, -2, -5, -12,
    -- layer=1 filter=219 channel=42
    -10, -2, 2, 8, 1, -11, 8, -8, 3,
    -- layer=1 filter=219 channel=43
    4, -6, 3, -4, -9, -1, -7, 4, 4,
    -- layer=1 filter=219 channel=44
    0, 6, 4, 5, 3, -1, 3, 1, 8,
    -- layer=1 filter=219 channel=45
    7, -3, 3, 2, 0, 4, -2, -4, -5,
    -- layer=1 filter=219 channel=46
    -14, 3, 3, -7, -10, -8, 0, -3, -4,
    -- layer=1 filter=219 channel=47
    -4, 0, -13, -8, -10, 5, -2, 2, -6,
    -- layer=1 filter=219 channel=48
    -6, 0, 6, -1, -3, -5, -8, 2, -3,
    -- layer=1 filter=219 channel=49
    5, 6, -8, -4, -10, 2, 6, 4, -8,
    -- layer=1 filter=219 channel=50
    6, -1, -4, 6, -3, -7, 5, 7, 8,
    -- layer=1 filter=219 channel=51
    4, -1, -6, -2, -8, -2, 1, -7, 2,
    -- layer=1 filter=219 channel=52
    -5, -1, 8, 4, 7, 7, 2, 10, -5,
    -- layer=1 filter=219 channel=53
    -10, -2, 5, 5, 3, 4, 0, -5, 2,
    -- layer=1 filter=219 channel=54
    7, -8, -2, 7, -4, 1, -17, 0, -1,
    -- layer=1 filter=219 channel=55
    -13, -8, 0, 0, -13, -1, 0, 2, -10,
    -- layer=1 filter=219 channel=56
    -11, -9, 5, -2, 1, 2, 6, 5, 6,
    -- layer=1 filter=219 channel=57
    7, -1, 1, -4, -5, -9, -10, -2, 1,
    -- layer=1 filter=219 channel=58
    -11, -10, -1, 14, -1, 5, -4, -8, 5,
    -- layer=1 filter=219 channel=59
    6, 0, -10, 7, -11, -4, -4, -1, -6,
    -- layer=1 filter=219 channel=60
    0, 8, 0, -5, 10, 2, -7, 6, -5,
    -- layer=1 filter=219 channel=61
    10, 3, 3, 9, -10, -9, -8, -5, 7,
    -- layer=1 filter=219 channel=62
    -6, -4, -8, -13, 2, -3, -6, -3, 5,
    -- layer=1 filter=219 channel=63
    3, -2, -8, -1, 6, -4, -6, 6, 5,
    -- layer=1 filter=219 channel=64
    -1, -2, -6, 0, -7, -4, -8, 0, 4,
    -- layer=1 filter=219 channel=65
    -9, -1, -8, -3, 3, 1, -8, 4, -7,
    -- layer=1 filter=219 channel=66
    5, -11, -2, 6, -5, 2, 7, 7, -8,
    -- layer=1 filter=219 channel=67
    9, -6, -4, -9, 0, -7, -9, -3, 2,
    -- layer=1 filter=219 channel=68
    -1, -2, -9, -11, 0, -9, -5, -4, 4,
    -- layer=1 filter=219 channel=69
    9, -3, -12, -2, -1, 0, -8, -12, -5,
    -- layer=1 filter=219 channel=70
    -3, -1, -7, 1, 3, 9, -8, -4, 7,
    -- layer=1 filter=219 channel=71
    1, 1, -2, -8, 0, -5, -2, 8, 0,
    -- layer=1 filter=219 channel=72
    -2, -3, -5, 5, -1, -7, -5, 7, 3,
    -- layer=1 filter=219 channel=73
    9, 6, 1, -2, 0, -2, 4, -2, 1,
    -- layer=1 filter=219 channel=74
    -2, 2, 6, 3, 4, 5, 1, -10, 7,
    -- layer=1 filter=219 channel=75
    -7, -5, -8, -8, -1, 0, 0, 3, -3,
    -- layer=1 filter=219 channel=76
    -8, -3, 3, 0, 8, -11, -3, 4, -3,
    -- layer=1 filter=219 channel=77
    -6, -10, 5, -3, -6, -7, 1, -5, -10,
    -- layer=1 filter=219 channel=78
    0, -10, 4, 9, -2, -11, -2, 0, 8,
    -- layer=1 filter=219 channel=79
    -5, 4, 3, 1, -13, -8, 8, -6, -3,
    -- layer=1 filter=219 channel=80
    4, -3, -7, 1, 6, -8, 9, 7, 10,
    -- layer=1 filter=219 channel=81
    3, -6, -8, 0, 2, -2, -3, -1, 8,
    -- layer=1 filter=219 channel=82
    -2, -7, -3, -9, 1, 3, 0, 8, -6,
    -- layer=1 filter=219 channel=83
    -2, 2, -10, -4, -8, -7, -3, -8, 4,
    -- layer=1 filter=219 channel=84
    7, 8, 7, -5, -8, 10, 0, -4, 2,
    -- layer=1 filter=219 channel=85
    2, 2, 6, -8, -5, 2, -3, 5, 1,
    -- layer=1 filter=219 channel=86
    2, -2, 5, 3, 0, -8, 8, 3, 6,
    -- layer=1 filter=219 channel=87
    -10, 9, 5, 3, -5, -8, -9, -3, -5,
    -- layer=1 filter=219 channel=88
    -9, -12, -5, -3, 0, 5, 0, 6, 5,
    -- layer=1 filter=219 channel=89
    -9, 1, -6, 3, 7, -3, -8, 0, -11,
    -- layer=1 filter=219 channel=90
    -2, -10, -10, 3, -9, 1, 8, 5, 1,
    -- layer=1 filter=219 channel=91
    -11, -11, -10, -5, 6, -10, -7, 0, 1,
    -- layer=1 filter=219 channel=92
    2, -11, 7, -3, 2, 6, 8, 0, 5,
    -- layer=1 filter=219 channel=93
    6, -3, 2, 0, 4, -5, 4, -2, -8,
    -- layer=1 filter=219 channel=94
    -8, 4, -7, 1, 5, -3, 0, -9, 5,
    -- layer=1 filter=219 channel=95
    -5, -10, 1, 9, -5, -2, -5, -6, 6,
    -- layer=1 filter=219 channel=96
    -10, 8, -9, -5, -7, -11, 7, -3, -3,
    -- layer=1 filter=219 channel=97
    7, -6, -3, 0, 5, -3, -2, -9, 0,
    -- layer=1 filter=219 channel=98
    7, 8, 1, -14, -4, -8, 0, -10, 7,
    -- layer=1 filter=219 channel=99
    8, 5, -8, 2, -11, -9, 2, -11, 4,
    -- layer=1 filter=219 channel=100
    -1, 4, 3, 5, -1, 4, 0, 7, 6,
    -- layer=1 filter=219 channel=101
    4, 0, -8, 1, -7, 0, 3, 7, 7,
    -- layer=1 filter=219 channel=102
    0, 4, 1, 0, 5, -10, 0, -5, 3,
    -- layer=1 filter=219 channel=103
    -6, -2, 7, 7, -1, 0, -4, 6, 4,
    -- layer=1 filter=219 channel=104
    2, 0, -6, 8, -7, -4, 6, 6, 1,
    -- layer=1 filter=219 channel=105
    -10, -2, -4, -10, 4, -2, -12, -8, -4,
    -- layer=1 filter=219 channel=106
    8, 5, 7, -5, -9, -14, 4, -8, -11,
    -- layer=1 filter=219 channel=107
    0, 3, 8, -3, 1, -8, 5, -6, -9,
    -- layer=1 filter=219 channel=108
    5, -11, -5, -1, -5, 3, 1, -7, -5,
    -- layer=1 filter=219 channel=109
    -4, 0, 0, 0, -6, 0, -6, -3, 5,
    -- layer=1 filter=219 channel=110
    -7, -3, -11, -2, -11, 0, 1, -2, 0,
    -- layer=1 filter=219 channel=111
    -1, -5, -8, 3, 0, 8, 0, 0, -5,
    -- layer=1 filter=219 channel=112
    7, -11, 0, -2, 6, 6, 4, -10, 0,
    -- layer=1 filter=219 channel=113
    -5, -2, 3, -1, 0, -7, -3, 6, -2,
    -- layer=1 filter=219 channel=114
    -1, 4, 6, -7, -12, 3, 0, 6, 1,
    -- layer=1 filter=219 channel=115
    -11, -8, -2, -4, 2, 4, 3, -1, -7,
    -- layer=1 filter=219 channel=116
    -10, -10, 3, -3, 7, 9, -3, 0, 10,
    -- layer=1 filter=219 channel=117
    -6, 2, 2, 0, -4, 2, 2, -5, -10,
    -- layer=1 filter=219 channel=118
    -6, -8, -6, -6, 0, 5, -6, 6, -10,
    -- layer=1 filter=219 channel=119
    -5, -8, -6, -9, -7, 2, 7, -6, -5,
    -- layer=1 filter=219 channel=120
    -12, 0, -16, -8, -10, -1, 0, 0, 0,
    -- layer=1 filter=219 channel=121
    -6, -4, -10, -1, 4, -9, -6, -1, -7,
    -- layer=1 filter=219 channel=122
    3, 1, 4, 9, 8, -4, 4, -1, 4,
    -- layer=1 filter=219 channel=123
    -9, -11, -7, 6, -11, -9, 0, -3, -6,
    -- layer=1 filter=219 channel=124
    11, -3, -5, -8, 0, 0, 1, 2, 6,
    -- layer=1 filter=219 channel=125
    -3, -11, 0, -7, -5, 8, -4, 5, 5,
    -- layer=1 filter=219 channel=126
    -8, -2, 6, -3, 0, -8, 0, -7, 1,
    -- layer=1 filter=219 channel=127
    -7, 8, -9, 9, -3, 0, -2, 9, 4,
    -- layer=1 filter=220 channel=0
    -5, -10, 1, 2, -2, -4, 2, -7, 2,
    -- layer=1 filter=220 channel=1
    8, -9, -4, -9, 5, -3, -9, 1, -7,
    -- layer=1 filter=220 channel=2
    -5, 0, -8, -7, 4, 0, -7, 6, 9,
    -- layer=1 filter=220 channel=3
    -3, -8, -5, -1, -2, -6, -5, 4, 3,
    -- layer=1 filter=220 channel=4
    -7, -2, 0, -7, -2, -5, 0, -9, 5,
    -- layer=1 filter=220 channel=5
    -4, -10, 6, -10, -8, -3, 2, -6, -8,
    -- layer=1 filter=220 channel=6
    1, 4, -6, 4, 5, 7, 6, -4, 10,
    -- layer=1 filter=220 channel=7
    -7, -6, 1, -9, -5, 0, -5, -2, 4,
    -- layer=1 filter=220 channel=8
    -7, -6, -8, -12, -13, -11, -5, 1, 0,
    -- layer=1 filter=220 channel=9
    2, 4, 7, -8, 0, 2, -9, 5, 3,
    -- layer=1 filter=220 channel=10
    -3, 5, -10, -5, 1, 2, -4, 0, 1,
    -- layer=1 filter=220 channel=11
    0, -9, -7, -1, -5, -8, 8, -6, 5,
    -- layer=1 filter=220 channel=12
    10, -4, 3, -10, 3, -4, -3, -8, -10,
    -- layer=1 filter=220 channel=13
    -1, 2, -5, 1, 1, -3, -5, -4, -5,
    -- layer=1 filter=220 channel=14
    1, 1, -7, 3, 0, 2, 2, 4, 3,
    -- layer=1 filter=220 channel=15
    -9, 3, 3, -2, 5, 8, 7, -1, -2,
    -- layer=1 filter=220 channel=16
    8, 1, 8, 0, 7, -10, 7, -6, 4,
    -- layer=1 filter=220 channel=17
    2, -11, 0, -6, -10, 3, 4, -10, -10,
    -- layer=1 filter=220 channel=18
    -11, -8, 5, 4, -8, 4, -7, 5, -7,
    -- layer=1 filter=220 channel=19
    -5, 7, -7, -5, -2, -10, -2, 3, -10,
    -- layer=1 filter=220 channel=20
    4, -4, 0, 0, -6, 2, 0, -9, 5,
    -- layer=1 filter=220 channel=21
    -10, 5, -7, -1, -12, -6, 4, 3, -1,
    -- layer=1 filter=220 channel=22
    -11, -7, 4, 1, -1, 1, 1, -10, 0,
    -- layer=1 filter=220 channel=23
    0, 0, -5, -9, 7, -10, 0, -8, -4,
    -- layer=1 filter=220 channel=24
    6, -8, -7, -2, -8, -6, 1, 4, -10,
    -- layer=1 filter=220 channel=25
    -8, 10, -1, 0, -13, 1, 7, -8, 3,
    -- layer=1 filter=220 channel=26
    0, -4, -4, -1, -13, 6, 0, -7, 0,
    -- layer=1 filter=220 channel=27
    -7, -1, -5, -3, -4, 5, -1, 7, 6,
    -- layer=1 filter=220 channel=28
    -6, -7, -5, 5, 6, -4, -5, -8, 0,
    -- layer=1 filter=220 channel=29
    -11, 7, 6, 2, 6, -8, -3, 5, -9,
    -- layer=1 filter=220 channel=30
    -3, -7, 7, 3, 5, -5, -11, 0, 3,
    -- layer=1 filter=220 channel=31
    4, 1, 7, -5, -2, -8, 0, -10, 5,
    -- layer=1 filter=220 channel=32
    7, 3, -4, 9, -1, 6, -4, -2, -7,
    -- layer=1 filter=220 channel=33
    -8, -2, -4, 2, -5, -7, 0, -1, -4,
    -- layer=1 filter=220 channel=34
    -5, 2, 2, 0, -3, -3, -6, -3, 1,
    -- layer=1 filter=220 channel=35
    0, 3, -1, -3, 2, 7, -9, -8, -4,
    -- layer=1 filter=220 channel=36
    0, 3, -10, 4, -8, -3, 0, 0, 8,
    -- layer=1 filter=220 channel=37
    -11, -10, -4, 9, 6, 5, -6, -9, 9,
    -- layer=1 filter=220 channel=38
    2, 1, 8, -2, -6, -9, 1, 1, 0,
    -- layer=1 filter=220 channel=39
    -10, -10, 3, 6, -2, 4, 6, 0, 1,
    -- layer=1 filter=220 channel=40
    -4, -3, -2, 1, -2, -8, 1, -3, -12,
    -- layer=1 filter=220 channel=41
    6, -1, 6, -5, -2, -3, -10, -4, -4,
    -- layer=1 filter=220 channel=42
    -5, 4, 4, -1, 5, 3, 3, -8, 8,
    -- layer=1 filter=220 channel=43
    -10, 4, -1, 5, -2, -11, 4, 0, -8,
    -- layer=1 filter=220 channel=44
    -10, -7, -5, -9, -2, -8, 7, -8, -6,
    -- layer=1 filter=220 channel=45
    -10, 9, -11, 6, -2, -6, -3, -7, -5,
    -- layer=1 filter=220 channel=46
    -2, -6, -10, -10, -4, -5, -10, -8, 5,
    -- layer=1 filter=220 channel=47
    -9, 0, 3, 0, -3, -1, 0, 1, -1,
    -- layer=1 filter=220 channel=48
    -10, -3, 8, -5, 7, 2, -9, 5, -8,
    -- layer=1 filter=220 channel=49
    -6, -10, -4, 7, 1, -7, -11, -5, -10,
    -- layer=1 filter=220 channel=50
    3, -3, -10, -9, -2, -8, 4, 1, 1,
    -- layer=1 filter=220 channel=51
    -2, -10, 6, -5, 0, -10, -1, -6, -8,
    -- layer=1 filter=220 channel=52
    -1, 5, 5, -2, 10, 0, 1, -9, 9,
    -- layer=1 filter=220 channel=53
    -7, -1, -10, -8, -5, -6, -11, -2, -8,
    -- layer=1 filter=220 channel=54
    -5, 2, -3, 7, -1, -8, 4, 4, -4,
    -- layer=1 filter=220 channel=55
    -1, 2, -13, 5, -5, 6, -4, -5, -3,
    -- layer=1 filter=220 channel=56
    -3, 0, -10, -5, 0, -1, -5, 5, -2,
    -- layer=1 filter=220 channel=57
    5, 2, 1, 0, 9, -4, -11, 1, -6,
    -- layer=1 filter=220 channel=58
    -2, 10, 8, -4, 0, 4, -8, 8, 7,
    -- layer=1 filter=220 channel=59
    0, 6, 3, -2, 0, -4, 8, 1, -3,
    -- layer=1 filter=220 channel=60
    -9, -2, 0, 7, -7, -2, 4, 4, 3,
    -- layer=1 filter=220 channel=61
    -6, -4, 6, -7, 9, 0, 1, 9, 0,
    -- layer=1 filter=220 channel=62
    0, -9, -3, 1, 7, -5, 3, 5, -6,
    -- layer=1 filter=220 channel=63
    8, 7, -1, -8, 0, -3, -3, 0, -1,
    -- layer=1 filter=220 channel=64
    -3, 5, -8, -10, -11, -3, -1, 0, -2,
    -- layer=1 filter=220 channel=65
    1, -3, -2, 7, 0, 1, 8, -7, -4,
    -- layer=1 filter=220 channel=66
    -2, -10, 6, -1, -8, -10, -3, -7, 0,
    -- layer=1 filter=220 channel=67
    0, 7, -3, -4, 8, -10, 8, 2, -4,
    -- layer=1 filter=220 channel=68
    7, -6, -11, 6, -11, 0, 5, -2, -7,
    -- layer=1 filter=220 channel=69
    8, -6, 3, -3, -14, -6, 0, -5, 8,
    -- layer=1 filter=220 channel=70
    -2, -6, 0, 7, 6, -10, -1, 3, 8,
    -- layer=1 filter=220 channel=71
    6, 0, 6, -7, -2, 3, -8, -3, -9,
    -- layer=1 filter=220 channel=72
    1, 0, -2, 1, 3, 8, 7, -3, -3,
    -- layer=1 filter=220 channel=73
    -1, -3, 1, 0, 1, 8, 7, 0, -6,
    -- layer=1 filter=220 channel=74
    -8, -12, -7, 2, -10, 8, 6, -3, 0,
    -- layer=1 filter=220 channel=75
    2, -3, -2, 5, 5, 9, -5, -9, -6,
    -- layer=1 filter=220 channel=76
    -2, 5, -5, -7, -6, 0, -8, -3, 2,
    -- layer=1 filter=220 channel=77
    -5, -11, 5, -6, 0, -3, -11, -1, -11,
    -- layer=1 filter=220 channel=78
    -7, 6, -8, -7, 2, 4, 5, 1, -5,
    -- layer=1 filter=220 channel=79
    6, 3, 4, -1, 1, 10, 6, -11, 2,
    -- layer=1 filter=220 channel=80
    -8, 7, 2, 7, -9, -5, -9, 0, 9,
    -- layer=1 filter=220 channel=81
    7, 4, 6, 1, -2, 6, 2, -9, 0,
    -- layer=1 filter=220 channel=82
    5, 5, -8, 2, -7, 4, -9, 3, -4,
    -- layer=1 filter=220 channel=83
    -11, -9, -2, -2, 7, -2, 1, -4, -2,
    -- layer=1 filter=220 channel=84
    -1, 0, 0, 4, -7, -8, -9, -9, 6,
    -- layer=1 filter=220 channel=85
    1, -6, 5, -1, -8, 8, -2, -5, 4,
    -- layer=1 filter=220 channel=86
    1, 3, 4, -10, -3, 6, -2, 5, 8,
    -- layer=1 filter=220 channel=87
    5, 0, -11, 5, -9, -5, 6, -6, 8,
    -- layer=1 filter=220 channel=88
    -3, -8, 4, 6, 7, -7, 4, 8, 9,
    -- layer=1 filter=220 channel=89
    7, -1, -3, -5, 0, -2, 5, 0, 3,
    -- layer=1 filter=220 channel=90
    6, 2, 7, -1, 7, -2, -11, -8, 1,
    -- layer=1 filter=220 channel=91
    -1, 1, -9, -2, 8, 9, 8, 2, -2,
    -- layer=1 filter=220 channel=92
    0, 3, -5, -7, 0, 5, -7, -1, -10,
    -- layer=1 filter=220 channel=93
    -9, -10, -8, 1, 0, 6, -9, -10, -8,
    -- layer=1 filter=220 channel=94
    -3, -7, 2, 8, 3, -3, -10, 7, -5,
    -- layer=1 filter=220 channel=95
    -11, -8, -11, -8, -9, -10, -6, -3, 5,
    -- layer=1 filter=220 channel=96
    -9, 7, 0, -10, -8, 0, -7, 7, -7,
    -- layer=1 filter=220 channel=97
    -6, -3, -3, -1, 0, -3, 4, 0, -11,
    -- layer=1 filter=220 channel=98
    -10, 2, 5, 1, 7, 0, 2, 9, -5,
    -- layer=1 filter=220 channel=99
    -4, 5, -7, 5, 2, -3, 0, -3, -4,
    -- layer=1 filter=220 channel=100
    2, -4, 8, 0, 0, 6, 8, -1, -7,
    -- layer=1 filter=220 channel=101
    -9, -2, 2, 5, 7, 5, 5, 7, -6,
    -- layer=1 filter=220 channel=102
    0, -10, -6, -3, 4, 4, 5, -13, -9,
    -- layer=1 filter=220 channel=103
    -8, 6, -9, -6, 0, -6, 7, -2, -7,
    -- layer=1 filter=220 channel=104
    -3, -4, -2, 0, 4, -3, 7, 0, -4,
    -- layer=1 filter=220 channel=105
    -10, 0, -6, -6, 9, -6, 0, 0, 2,
    -- layer=1 filter=220 channel=106
    4, -7, 0, -4, -2, -2, 1, -4, 3,
    -- layer=1 filter=220 channel=107
    -3, 9, -5, 9, -2, 7, 10, 0, -11,
    -- layer=1 filter=220 channel=108
    -6, -3, 3, -5, -1, 5, -2, 2, 1,
    -- layer=1 filter=220 channel=109
    4, -3, 1, 2, -8, -2, 9, 5, -1,
    -- layer=1 filter=220 channel=110
    -9, 0, 2, 0, 2, 6, 3, -13, -9,
    -- layer=1 filter=220 channel=111
    -7, -3, 2, -8, 9, -2, 5, 8, -6,
    -- layer=1 filter=220 channel=112
    1, 5, 4, -8, -1, 0, 4, 1, -12,
    -- layer=1 filter=220 channel=113
    6, -9, 5, 2, -1, 2, -11, 3, 1,
    -- layer=1 filter=220 channel=114
    -1, -1, -12, 0, -5, 3, 3, 2, -7,
    -- layer=1 filter=220 channel=115
    -8, -3, 6, -10, -4, 3, 0, -8, 6,
    -- layer=1 filter=220 channel=116
    -7, 10, 7, 2, 8, 10, 8, 9, -3,
    -- layer=1 filter=220 channel=117
    5, 4, 8, -5, -8, 5, -7, 9, 8,
    -- layer=1 filter=220 channel=118
    1, -3, 0, -3, -4, 4, 1, 5, -8,
    -- layer=1 filter=220 channel=119
    0, 5, 0, 7, -5, -1, -10, 6, 7,
    -- layer=1 filter=220 channel=120
    1, -8, 4, -7, 4, -10, 1, -3, 5,
    -- layer=1 filter=220 channel=121
    7, -7, 0, -8, 6, -9, -6, 9, 2,
    -- layer=1 filter=220 channel=122
    0, -10, -1, -6, 4, 1, 8, -1, 2,
    -- layer=1 filter=220 channel=123
    7, 2, -10, 4, 2, 7, 3, -2, 4,
    -- layer=1 filter=220 channel=124
    -4, 8, -3, 8, 2, 0, -4, -7, -2,
    -- layer=1 filter=220 channel=125
    0, 5, 5, -9, -1, 5, 5, 6, -3,
    -- layer=1 filter=220 channel=126
    -1, -11, 5, 0, -3, 0, -4, 1, 5,
    -- layer=1 filter=220 channel=127
    -7, -3, -8, -1, 10, -7, 3, 6, -6,
    -- layer=1 filter=221 channel=0
    -5, -8, 2, 3, -10, -8, 5, 1, -2,
    -- layer=1 filter=221 channel=1
    3, 8, 4, -12, -8, -2, -2, -10, -8,
    -- layer=1 filter=221 channel=2
    -9, -13, -4, -10, -1, 2, 1, -13, 0,
    -- layer=1 filter=221 channel=3
    -9, -7, 4, 4, 9, -9, -9, 0, -4,
    -- layer=1 filter=221 channel=4
    1, -11, 0, -6, 0, -8, 6, -2, 1,
    -- layer=1 filter=221 channel=5
    3, -7, 2, 6, 0, -4, 0, -18, -12,
    -- layer=1 filter=221 channel=6
    -7, 0, -12, 8, 1, -2, -8, 2, -7,
    -- layer=1 filter=221 channel=7
    -7, 4, 1, -6, 7, 7, 7, 5, 0,
    -- layer=1 filter=221 channel=8
    -6, -5, -12, 7, -5, -8, 9, -10, 0,
    -- layer=1 filter=221 channel=9
    15, 2, 6, 0, -8, 8, 9, 3, -9,
    -- layer=1 filter=221 channel=10
    6, 0, 4, 10, -6, -2, -3, -11, 7,
    -- layer=1 filter=221 channel=11
    2, -8, 1, -12, 3, 5, -12, 0, 3,
    -- layer=1 filter=221 channel=12
    -1, -6, -6, -8, -1, -7, -7, -9, 7,
    -- layer=1 filter=221 channel=13
    -7, -4, 2, -10, -2, 4, -7, 1, -9,
    -- layer=1 filter=221 channel=14
    -12, -7, 0, 6, -6, -12, -2, 6, -2,
    -- layer=1 filter=221 channel=15
    4, 2, -6, 8, 7, -2, 6, -3, 3,
    -- layer=1 filter=221 channel=16
    2, -12, -12, -5, -1, 5, 6, 2, 0,
    -- layer=1 filter=221 channel=17
    -1, 0, 1, -13, 9, -1, 7, -1, -8,
    -- layer=1 filter=221 channel=18
    0, -5, -8, -9, -3, -1, 0, -5, 4,
    -- layer=1 filter=221 channel=19
    2, -7, -2, -2, -10, 4, 0, -11, -11,
    -- layer=1 filter=221 channel=20
    -14, -5, -2, 6, -12, 3, -9, -4, 0,
    -- layer=1 filter=221 channel=21
    -4, 4, -4, -2, -3, -11, -10, 0, -14,
    -- layer=1 filter=221 channel=22
    -6, -12, -3, 8, -11, -1, -5, -3, 5,
    -- layer=1 filter=221 channel=23
    -1, -1, -8, -3, -5, -12, 3, -12, -3,
    -- layer=1 filter=221 channel=24
    -3, -2, 0, 0, -10, -1, -15, -3, 1,
    -- layer=1 filter=221 channel=25
    4, -11, -7, -6, -6, 2, -9, -7, -1,
    -- layer=1 filter=221 channel=26
    5, 8, -6, -15, -2, -1, -5, -9, 4,
    -- layer=1 filter=221 channel=27
    -14, 6, 1, -7, -9, 0, -7, -5, 3,
    -- layer=1 filter=221 channel=28
    -5, -8, 1, 9, 7, -8, -4, 0, -5,
    -- layer=1 filter=221 channel=29
    -11, -11, 0, 3, 3, -7, 7, 0, 0,
    -- layer=1 filter=221 channel=30
    1, 1, -12, 3, -6, -2, 7, 6, -11,
    -- layer=1 filter=221 channel=31
    -1, -2, 6, 6, -6, -11, 3, 4, -9,
    -- layer=1 filter=221 channel=32
    -3, -9, -5, -3, 5, 8, -11, -5, 4,
    -- layer=1 filter=221 channel=33
    1, -2, -7, 5, 0, 1, -9, 2, -3,
    -- layer=1 filter=221 channel=34
    -6, -5, -5, -9, -9, -3, -10, 1, 5,
    -- layer=1 filter=221 channel=35
    1, 0, -6, 1, -2, -8, 0, -11, -3,
    -- layer=1 filter=221 channel=36
    -9, -16, -6, -12, -1, 9, 3, -2, 5,
    -- layer=1 filter=221 channel=37
    3, 0, -7, 7, -7, -8, -5, -3, -2,
    -- layer=1 filter=221 channel=38
    -6, -11, -9, -13, -1, -5, 1, 2, -10,
    -- layer=1 filter=221 channel=39
    8, -8, 3, -3, -4, 8, 5, -12, 5,
    -- layer=1 filter=221 channel=40
    -2, 0, 0, -7, -4, 0, 0, -7, -2,
    -- layer=1 filter=221 channel=41
    6, -10, -4, -8, 7, 3, 0, 4, 8,
    -- layer=1 filter=221 channel=42
    -4, 4, -1, -3, 5, 2, -8, 7, 1,
    -- layer=1 filter=221 channel=43
    0, 8, -5, -7, -4, -7, 0, -4, -7,
    -- layer=1 filter=221 channel=44
    0, -8, 7, 3, 5, 13, -1, -12, -4,
    -- layer=1 filter=221 channel=45
    -13, -8, -4, -8, 0, 4, 5, -6, 5,
    -- layer=1 filter=221 channel=46
    1, 0, 1, 11, -12, 0, -9, 0, -6,
    -- layer=1 filter=221 channel=47
    1, 10, -10, -4, -12, 1, 0, -7, 0,
    -- layer=1 filter=221 channel=48
    -11, -7, -10, 7, -10, 0, -3, -4, -4,
    -- layer=1 filter=221 channel=49
    -8, 3, -1, 1, 2, -3, -4, -1, -10,
    -- layer=1 filter=221 channel=50
    -4, 7, -7, -7, -5, -10, 4, 6, 2,
    -- layer=1 filter=221 channel=51
    -3, 6, 4, -1, 0, 0, -2, 0, 1,
    -- layer=1 filter=221 channel=52
    -1, -4, -7, 10, 0, -5, 9, 3, 8,
    -- layer=1 filter=221 channel=53
    0, -1, 0, -9, -8, -1, -2, 4, -11,
    -- layer=1 filter=221 channel=54
    3, -15, -10, 7, 5, -5, 5, -11, -2,
    -- layer=1 filter=221 channel=55
    -11, -4, -8, -6, -2, -4, -10, 0, 1,
    -- layer=1 filter=221 channel=56
    -8, 7, -5, 11, 9, 10, 10, -4, 11,
    -- layer=1 filter=221 channel=57
    9, 1, -2, -5, -5, 1, 9, -2, 4,
    -- layer=1 filter=221 channel=58
    13, 9, -8, 8, 0, 2, -3, 6, -1,
    -- layer=1 filter=221 channel=59
    -5, -4, 8, 8, -2, -8, 2, 6, 8,
    -- layer=1 filter=221 channel=60
    -8, 0, 6, -8, -4, -11, -1, -3, 3,
    -- layer=1 filter=221 channel=61
    -11, 10, -10, -4, 0, -1, -4, 0, 8,
    -- layer=1 filter=221 channel=62
    6, 0, 3, 0, 0, 4, 0, -17, 10,
    -- layer=1 filter=221 channel=63
    -7, -12, -8, -14, 5, 2, -5, 8, -1,
    -- layer=1 filter=221 channel=64
    -6, -10, 1, 3, -9, 0, -6, 0, 3,
    -- layer=1 filter=221 channel=65
    -4, 5, -2, 4, 2, -11, 4, 2, 1,
    -- layer=1 filter=221 channel=66
    -13, 7, -12, -3, -4, -7, -4, -9, -7,
    -- layer=1 filter=221 channel=67
    -6, -1, -2, -9, -2, 11, 10, -5, 2,
    -- layer=1 filter=221 channel=68
    -1, -3, 7, -4, -1, -5, 0, -6, 8,
    -- layer=1 filter=221 channel=69
    -2, -7, -5, -8, -9, -1, -4, -11, -2,
    -- layer=1 filter=221 channel=70
    -6, 0, 3, 3, -8, -9, -6, -4, 6,
    -- layer=1 filter=221 channel=71
    1, -3, -7, 10, -1, -3, -2, -7, 3,
    -- layer=1 filter=221 channel=72
    0, -11, -6, 0, -11, 9, -6, 2, -3,
    -- layer=1 filter=221 channel=73
    -11, 3, 9, 5, -2, -7, 6, -7, 9,
    -- layer=1 filter=221 channel=74
    2, 4, -5, -10, -9, 1, 8, -11, 0,
    -- layer=1 filter=221 channel=75
    6, -9, -5, 5, -3, -8, 6, 2, 0,
    -- layer=1 filter=221 channel=76
    -4, 5, 8, -1, 1, -2, -10, 5, -9,
    -- layer=1 filter=221 channel=77
    -11, 1, 2, -5, 8, -9, -2, 3, 5,
    -- layer=1 filter=221 channel=78
    -3, 0, 7, 0, 5, -6, -4, -6, 0,
    -- layer=1 filter=221 channel=79
    5, -13, -7, -8, -3, 3, -11, -11, 1,
    -- layer=1 filter=221 channel=80
    8, 3, 0, 2, -11, 4, -6, -9, -7,
    -- layer=1 filter=221 channel=81
    7, -9, -9, -2, 1, 2, 1, -1, 0,
    -- layer=1 filter=221 channel=82
    -1, -1, -1, -1, -4, 0, 5, -5, 1,
    -- layer=1 filter=221 channel=83
    -4, -6, -9, 0, -8, -7, 6, -4, 0,
    -- layer=1 filter=221 channel=84
    -16, -5, 0, -11, 11, 6, 7, 1, -4,
    -- layer=1 filter=221 channel=85
    9, -1, -12, -4, 8, -9, -10, -4, -7,
    -- layer=1 filter=221 channel=86
    -15, -2, -3, -15, -2, 1, -5, 0, -14,
    -- layer=1 filter=221 channel=87
    7, -9, -1, 3, 8, 0, -11, 3, 5,
    -- layer=1 filter=221 channel=88
    0, 5, 2, -5, -2, 6, -4, -9, -11,
    -- layer=1 filter=221 channel=89
    5, -9, -7, -3, -3, -1, 7, -5, -6,
    -- layer=1 filter=221 channel=90
    -10, 9, -7, -2, -9, 3, -8, 6, 5,
    -- layer=1 filter=221 channel=91
    -6, 5, -6, -3, 0, -13, -13, -6, -6,
    -- layer=1 filter=221 channel=92
    -2, -4, -9, -11, -7, -6, -1, 7, 2,
    -- layer=1 filter=221 channel=93
    0, -4, -17, 0, -10, -17, -13, -6, 1,
    -- layer=1 filter=221 channel=94
    8, -4, -4, -9, 1, -7, -11, 0, -5,
    -- layer=1 filter=221 channel=95
    4, -9, -10, -15, -1, 7, 3, -11, 3,
    -- layer=1 filter=221 channel=96
    5, 2, -8, -10, -5, -5, -12, -8, 8,
    -- layer=1 filter=221 channel=97
    -6, -13, -11, 0, -13, 7, -1, -13, -2,
    -- layer=1 filter=221 channel=98
    0, -6, -10, 0, -1, -7, -2, -6, 2,
    -- layer=1 filter=221 channel=99
    -2, -7, -1, 8, -5, 7, 4, 7, 5,
    -- layer=1 filter=221 channel=100
    -11, -2, 4, 3, 3, 9, -8, 9, 4,
    -- layer=1 filter=221 channel=101
    5, -4, -1, 1, 5, 3, -1, -2, 0,
    -- layer=1 filter=221 channel=102
    -6, 7, -3, 4, 0, 6, 1, -9, 1,
    -- layer=1 filter=221 channel=103
    -4, 0, 1, 8, 4, -10, -2, 0, -5,
    -- layer=1 filter=221 channel=104
    8, -8, -9, -5, 2, -8, 4, 8, -11,
    -- layer=1 filter=221 channel=105
    7, 5, -8, -7, 0, 8, 1, 1, -7,
    -- layer=1 filter=221 channel=106
    3, -10, -2, -4, -10, -7, -1, -4, -13,
    -- layer=1 filter=221 channel=107
    -4, 0, 9, 3, 7, -5, -4, -8, 5,
    -- layer=1 filter=221 channel=108
    -3, -1, 6, -1, -8, 13, -1, -4, 11,
    -- layer=1 filter=221 channel=109
    -3, 0, 5, -7, 5, 4, -3, 0, -2,
    -- layer=1 filter=221 channel=110
    3, 0, -2, -10, 5, -6, -12, -1, -1,
    -- layer=1 filter=221 channel=111
    -2, -4, -1, -11, 0, -4, -11, -5, -13,
    -- layer=1 filter=221 channel=112
    -8, -1, -7, -11, -6, 0, -7, 4, 8,
    -- layer=1 filter=221 channel=113
    -10, -1, -10, -4, -8, 5, 4, -4, -12,
    -- layer=1 filter=221 channel=114
    1, -1, 9, -7, -1, 1, 0, 6, -5,
    -- layer=1 filter=221 channel=115
    7, 0, -5, -4, 0, 0, 8, 0, 9,
    -- layer=1 filter=221 channel=116
    3, -3, -1, 3, -9, 8, -5, 0, 0,
    -- layer=1 filter=221 channel=117
    -12, 0, -5, -10, 0, -1, -1, -7, 9,
    -- layer=1 filter=221 channel=118
    -7, 7, 4, -4, 5, 0, -6, 8, 9,
    -- layer=1 filter=221 channel=119
    -3, 5, -9, 1, -1, -5, -14, -5, -2,
    -- layer=1 filter=221 channel=120
    3, -8, 0, -6, -5, -8, -9, 1, -9,
    -- layer=1 filter=221 channel=121
    -3, -1, 0, -2, -13, -11, 7, -6, -3,
    -- layer=1 filter=221 channel=122
    10, 9, -7, 8, 6, -8, 3, 5, 3,
    -- layer=1 filter=221 channel=123
    2, -8, 11, -1, 5, 4, -2, 2, 8,
    -- layer=1 filter=221 channel=124
    -4, -1, 7, 4, 7, -1, 0, 5, 3,
    -- layer=1 filter=221 channel=125
    6, -5, -3, 8, 2, 5, -5, -10, -9,
    -- layer=1 filter=221 channel=126
    -5, 8, -11, -3, 7, 5, -4, -8, 2,
    -- layer=1 filter=221 channel=127
    -10, 1, 5, -12, -12, -3, -9, -11, 0,
    -- layer=1 filter=222 channel=0
    1, -6, 15, 17, -1, -14, -8, -8, -2,
    -- layer=1 filter=222 channel=1
    12, -3, -34, 4, 8, 23, -6, 5, 2,
    -- layer=1 filter=222 channel=2
    -5, 11, 25, 33, 11, 24, 47, 35, 16,
    -- layer=1 filter=222 channel=3
    8, -1, 3, 1, -9, 3, -2, 4, 9,
    -- layer=1 filter=222 channel=4
    -2, 6, 7, 2, -7, 5, -3, 5, -7,
    -- layer=1 filter=222 channel=5
    26, -11, -33, 19, 26, 21, 17, 7, 0,
    -- layer=1 filter=222 channel=6
    -10, 3, -13, 5, -6, 24, -17, -1, 15,
    -- layer=1 filter=222 channel=7
    -23, -41, -30, -25, -68, -21, -17, 11, 4,
    -- layer=1 filter=222 channel=8
    12, -18, -44, 11, 31, 8, 0, 6, 6,
    -- layer=1 filter=222 channel=9
    8, 11, 27, 21, -6, 10, -3, -1, 16,
    -- layer=1 filter=222 channel=10
    -8, -36, -13, -7, -20, -19, -17, 9, 22,
    -- layer=1 filter=222 channel=11
    -6, -13, 0, -8, -3, -18, 8, 16, 16,
    -- layer=1 filter=222 channel=12
    12, 9, -14, 52, -1, -45, -1, 16, 11,
    -- layer=1 filter=222 channel=13
    11, -3, 25, -4, 20, 5, -20, -27, -9,
    -- layer=1 filter=222 channel=14
    -41, -31, -23, 4, -44, -35, -1, -4, -21,
    -- layer=1 filter=222 channel=15
    -35, -10, -44, -4, -25, -2, 14, -37, -21,
    -- layer=1 filter=222 channel=16
    26, -8, -14, 0, 24, 22, 6, 14, -15,
    -- layer=1 filter=222 channel=17
    11, 2, 21, 3, 10, -4, -8, 0, 7,
    -- layer=1 filter=222 channel=18
    -6, 10, 17, 28, 6, -10, 11, 22, 37,
    -- layer=1 filter=222 channel=19
    81, 40, 31, 80, 90, 66, 70, 66, 52,
    -- layer=1 filter=222 channel=20
    10, 15, 5, -5, 7, 27, -21, -12, -19,
    -- layer=1 filter=222 channel=21
    14, 24, 1, 3, -12, 22, -11, -13, -18,
    -- layer=1 filter=222 channel=22
    7, -4, -8, -12, -1, 3, -11, -4, -10,
    -- layer=1 filter=222 channel=23
    -28, 2, -18, -40, -58, 11, -20, -7, -19,
    -- layer=1 filter=222 channel=24
    20, -10, 24, 9, 12, 14, 4, -28, -4,
    -- layer=1 filter=222 channel=25
    -8, 4, -20, -20, -13, -2, 1, 20, 8,
    -- layer=1 filter=222 channel=26
    -9, 3, 17, -12, 0, -21, 0, -57, -9,
    -- layer=1 filter=222 channel=27
    5, 5, 9, 3, 10, 26, -3, 1, 9,
    -- layer=1 filter=222 channel=28
    -10, -14, -16, -20, -47, -4, -20, 5, -17,
    -- layer=1 filter=222 channel=29
    -10, 3, 20, -2, 9, 24, -18, 5, 26,
    -- layer=1 filter=222 channel=30
    14, -17, 14, 40, 43, 22, 12, 36, 39,
    -- layer=1 filter=222 channel=31
    3, -14, 17, 12, 14, 7, -8, 21, 15,
    -- layer=1 filter=222 channel=32
    -34, -17, -31, -7, -37, -29, -3, -42, 12,
    -- layer=1 filter=222 channel=33
    1, 12, -10, -7, -3, 10, -18, -17, -23,
    -- layer=1 filter=222 channel=34
    -12, 1, -4, -22, -26, 1, -8, -8, -2,
    -- layer=1 filter=222 channel=35
    -15, -7, -13, -14, -12, -23, 0, -4, -19,
    -- layer=1 filter=222 channel=36
    -14, -15, -10, -15, -16, -8, -18, 0, -3,
    -- layer=1 filter=222 channel=37
    25, 2, -14, 25, 27, 37, 36, 5, 18,
    -- layer=1 filter=222 channel=38
    8, 6, 14, 0, 10, 18, -7, -11, -8,
    -- layer=1 filter=222 channel=39
    4, -11, 7, -21, 0, -18, -18, -21, -9,
    -- layer=1 filter=222 channel=40
    -4, 6, 10, 13, 3, 0, -15, 8, 13,
    -- layer=1 filter=222 channel=41
    -6, -35, -1, 5, -29, 2, -23, -51, -12,
    -- layer=1 filter=222 channel=42
    -34, -8, 2, 10, 21, 29, 17, 31, 18,
    -- layer=1 filter=222 channel=43
    28, -4, -36, 0, -12, 2, 0, 25, -1,
    -- layer=1 filter=222 channel=44
    -35, -21, -20, -28, -21, -27, 0, -60, 7,
    -- layer=1 filter=222 channel=45
    11, -7, -5, -14, 11, -2, 1, -27, -13,
    -- layer=1 filter=222 channel=46
    71, 57, 38, 77, 71, 67, 78, 77, 38,
    -- layer=1 filter=222 channel=47
    -27, -7, -5, -5, -20, 16, 0, 14, 5,
    -- layer=1 filter=222 channel=48
    20, -2, 16, 13, 4, 9, -14, -19, -5,
    -- layer=1 filter=222 channel=49
    18, 1, 18, 19, 0, -2, -10, -12, -4,
    -- layer=1 filter=222 channel=50
    4, -6, 0, -12, -1, -6, -13, -12, -3,
    -- layer=1 filter=222 channel=51
    9, -12, 10, 8, -4, -9, -18, 3, -11,
    -- layer=1 filter=222 channel=52
    1, -8, -4, 13, -17, -1, 15, 20, 13,
    -- layer=1 filter=222 channel=53
    3, 8, -6, 17, 15, 11, 8, 21, 14,
    -- layer=1 filter=222 channel=54
    12, 5, -11, -10, 8, 12, 18, 26, 20,
    -- layer=1 filter=222 channel=55
    -22, -19, -13, 4, -17, -17, 17, 0, 3,
    -- layer=1 filter=222 channel=56
    7, 5, -10, -3, -2, 0, 3, -3, 10,
    -- layer=1 filter=222 channel=57
    -9, -48, -5, -9, -6, -13, -23, 8, 14,
    -- layer=1 filter=222 channel=58
    -29, -30, -13, -34, -8, 0, -11, 4, 16,
    -- layer=1 filter=222 channel=59
    3, 6, -15, 1, -4, -5, -3, 0, -7,
    -- layer=1 filter=222 channel=60
    3, -21, -5, 0, -13, -3, -5, 5, 7,
    -- layer=1 filter=222 channel=61
    -8, 13, -10, 6, -8, -5, -3, 5, 0,
    -- layer=1 filter=222 channel=62
    40, 4, -13, 4, 26, 26, 24, 12, 12,
    -- layer=1 filter=222 channel=63
    -8, 4, 2, 2, -16, -26, 2, -1, 1,
    -- layer=1 filter=222 channel=64
    0, 15, -9, 10, 9, 2, -1, 3, -8,
    -- layer=1 filter=222 channel=65
    19, 17, 22, -6, -13, 14, -30, -29, -23,
    -- layer=1 filter=222 channel=66
    2, 10, -9, -9, -13, -13, -14, 10, -12,
    -- layer=1 filter=222 channel=67
    18, 25, 12, 30, 29, 38, 17, 8, 13,
    -- layer=1 filter=222 channel=68
    -32, -29, -7, -37, -8, -32, -7, -49, 7,
    -- layer=1 filter=222 channel=69
    21, -24, -40, -3, 27, 15, 23, -16, 0,
    -- layer=1 filter=222 channel=70
    22, 23, 4, 11, 19, 21, 10, 19, 26,
    -- layer=1 filter=222 channel=71
    25, 21, 13, -5, -7, 4, -9, -9, -6,
    -- layer=1 filter=222 channel=72
    -2, -2, 0, 44, 42, 47, 26, 44, 44,
    -- layer=1 filter=222 channel=73
    -3, 6, -2, 0, 3, -3, -10, 2, -5,
    -- layer=1 filter=222 channel=74
    -5, -37, 0, 11, -9, 9, -16, 15, 40,
    -- layer=1 filter=222 channel=75
    -17, -7, -18, 41, 12, 8, 28, 45, 23,
    -- layer=1 filter=222 channel=76
    -9, -5, 1, 0, -13, -9, 0, -8, 9,
    -- layer=1 filter=222 channel=77
    18, 3, 10, -15, 6, -1, -26, -25, -8,
    -- layer=1 filter=222 channel=78
    3, -6, -2, -15, 13, 0, -12, 0, 4,
    -- layer=1 filter=222 channel=79
    20, -10, -12, -8, 19, 8, 13, -1, -3,
    -- layer=1 filter=222 channel=80
    18, 10, 16, 4, 11, 11, 5, 6, 9,
    -- layer=1 filter=222 channel=81
    18, 21, 4, -13, 3, 0, -11, -25, -4,
    -- layer=1 filter=222 channel=82
    7, 22, 10, 9, -2, 4, -13, -21, 0,
    -- layer=1 filter=222 channel=83
    -11, -18, -1, 4, 6, -8, -11, -33, 13,
    -- layer=1 filter=222 channel=84
    16, 23, 38, 40, 15, 4, 17, 36, 54,
    -- layer=1 filter=222 channel=85
    -40, -2, -14, -22, -3, -1, 2, -8, 18,
    -- layer=1 filter=222 channel=86
    -13, 0, -8, 5, -3, 17, -1, 8, 3,
    -- layer=1 filter=222 channel=87
    48, 22, -5, 51, 34, 35, 9, 51, 29,
    -- layer=1 filter=222 channel=88
    -2, -5, 14, 0, 10, -1, -12, -19, -26,
    -- layer=1 filter=222 channel=89
    4, 36, 16, 15, 3, 12, -21, -9, -12,
    -- layer=1 filter=222 channel=90
    -36, -46, -19, -52, -29, -46, -5, -63, -10,
    -- layer=1 filter=222 channel=91
    4, 6, 8, 11, 0, 11, -12, 4, 3,
    -- layer=1 filter=222 channel=92
    -12, -37, 2, -1, -23, 15, 10, -61, 31,
    -- layer=1 filter=222 channel=93
    19, 7, 0, 4, 2, 14, -16, -17, -4,
    -- layer=1 filter=222 channel=94
    -12, 0, -1, 10, -10, -5, -2, 3, 3,
    -- layer=1 filter=222 channel=95
    16, 6, 9, 44, 11, 6, 22, 42, 33,
    -- layer=1 filter=222 channel=96
    -3, -10, 3, -11, -11, -1, -1, -11, -6,
    -- layer=1 filter=222 channel=97
    18, 19, 9, -5, -11, 2, -20, -8, -8,
    -- layer=1 filter=222 channel=98
    14, -16, -10, 4, 10, 2, -1, 13, 16,
    -- layer=1 filter=222 channel=99
    8, -52, 5, 2, -16, -37, -3, 4, -4,
    -- layer=1 filter=222 channel=100
    -12, -11, -8, 1, 0, -2, 0, -13, 3,
    -- layer=1 filter=222 channel=101
    2, 11, 5, 4, -3, 16, -3, -3, -3,
    -- layer=1 filter=222 channel=102
    5, 9, 4, 19, -5, 15, -7, 0, 9,
    -- layer=1 filter=222 channel=103
    1, 7, -2, 19, 15, 6, 1, 4, 14,
    -- layer=1 filter=222 channel=104
    -22, 1, -23, -2, -17, 14, -4, 11, 7,
    -- layer=1 filter=222 channel=105
    6, 13, 18, 9, -2, -11, -20, -9, 0,
    -- layer=1 filter=222 channel=106
    8, 14, 3, 12, 3, -3, -7, -11, 7,
    -- layer=1 filter=222 channel=107
    -2, -17, -3, -16, -15, -6, -20, -3, -15,
    -- layer=1 filter=222 channel=108
    -13, -39, -29, -32, -27, -35, 12, -71, -17,
    -- layer=1 filter=222 channel=109
    1, -5, -2, -1, -7, 2, -4, 3, -3,
    -- layer=1 filter=222 channel=110
    6, 3, 8, 1, 7, 2, -2, -18, -6,
    -- layer=1 filter=222 channel=111
    27, -3, 33, 53, 28, -1, 15, 44, 49,
    -- layer=1 filter=222 channel=112
    22, 32, 15, 42, 19, 0, 36, 42, 58,
    -- layer=1 filter=222 channel=113
    5, -1, 5, 1, 5, 3, -10, 6, -23,
    -- layer=1 filter=222 channel=114
    -9, -10, -29, -22, -5, 2, -8, -22, -27,
    -- layer=1 filter=222 channel=115
    1, -9, 12, 7, -1, 8, -3, -7, 0,
    -- layer=1 filter=222 channel=116
    4, 3, -7, 0, -14, -10, 6, -6, -8,
    -- layer=1 filter=222 channel=117
    62, 62, 54, 84, 60, 19, 68, 71, 83,
    -- layer=1 filter=222 channel=118
    10, 3, 0, 32, 31, 3, 16, 28, 34,
    -- layer=1 filter=222 channel=119
    -29, -31, -15, -27, -28, -40, -5, -56, -8,
    -- layer=1 filter=222 channel=120
    6, 0, 5, -4, -1, 8, -15, -9, -2,
    -- layer=1 filter=222 channel=121
    14, 20, -11, 48, 37, 37, 31, 59, 11,
    -- layer=1 filter=222 channel=122
    10, 2, -1, -9, 3, 0, -3, -3, -6,
    -- layer=1 filter=222 channel=123
    -18, -8, -20, 7, -1, 13, 3, 18, -1,
    -- layer=1 filter=222 channel=124
    -10, 7, -7, 5, -1, 0, 0, 13, 0,
    -- layer=1 filter=222 channel=125
    22, 13, -3, 9, 25, 3, -8, 16, 2,
    -- layer=1 filter=222 channel=126
    18, -9, 5, 38, 57, 18, 30, 21, 41,
    -- layer=1 filter=222 channel=127
    -1, -5, 9, 50, 26, 16, 24, 59, 45,
    -- layer=1 filter=223 channel=0
    0, -3, -7, 8, 6, -1, 6, 2, 5,
    -- layer=1 filter=223 channel=1
    0, 8, -9, 6, 0, 8, 2, -10, -1,
    -- layer=1 filter=223 channel=2
    -11, -10, 7, 8, -12, 0, -3, 7, -5,
    -- layer=1 filter=223 channel=3
    5, 6, 4, -6, -1, 8, 8, 2, 1,
    -- layer=1 filter=223 channel=4
    -5, -8, 1, -7, 7, -2, 9, 6, -6,
    -- layer=1 filter=223 channel=5
    -4, -9, 9, 4, 7, -2, 6, -11, -2,
    -- layer=1 filter=223 channel=6
    8, -3, 6, -7, -6, -7, -6, -5, -2,
    -- layer=1 filter=223 channel=7
    -4, 4, 5, -1, -7, -2, 2, -9, 1,
    -- layer=1 filter=223 channel=8
    -6, -5, 2, 2, -8, 4, 6, 6, 5,
    -- layer=1 filter=223 channel=9
    0, 0, -8, 7, -7, 4, 0, 0, 0,
    -- layer=1 filter=223 channel=10
    0, -12, 0, 7, -3, 0, 0, -11, -10,
    -- layer=1 filter=223 channel=11
    2, 2, -10, -9, 3, -4, -12, -5, -3,
    -- layer=1 filter=223 channel=12
    7, 8, 1, -1, 6, 3, 5, -8, -6,
    -- layer=1 filter=223 channel=13
    -2, -1, -6, 0, 3, 3, -11, -7, -2,
    -- layer=1 filter=223 channel=14
    0, 6, 9, -2, 3, -6, 5, -5, -1,
    -- layer=1 filter=223 channel=15
    6, 0, -9, 7, -6, 3, -10, -4, -9,
    -- layer=1 filter=223 channel=16
    -7, -5, -9, -9, 10, -10, -4, -9, -1,
    -- layer=1 filter=223 channel=17
    8, 1, -6, 5, -9, -6, 3, 0, 0,
    -- layer=1 filter=223 channel=18
    7, -9, 0, -10, -5, 2, 9, 3, -3,
    -- layer=1 filter=223 channel=19
    0, 2, 1, -10, -1, 6, -10, 3, -12,
    -- layer=1 filter=223 channel=20
    1, 2, -1, -8, -8, 0, -7, -8, 3,
    -- layer=1 filter=223 channel=21
    -11, 1, -12, 0, -7, 2, 1, 2, 4,
    -- layer=1 filter=223 channel=22
    -11, 7, 8, -3, 8, -3, -4, -7, -10,
    -- layer=1 filter=223 channel=23
    -2, -3, 10, 1, -6, -4, 4, -1, -3,
    -- layer=1 filter=223 channel=24
    2, 6, -2, 0, -13, -3, 0, -9, 1,
    -- layer=1 filter=223 channel=25
    6, 1, 0, 0, 3, -11, -2, 3, -2,
    -- layer=1 filter=223 channel=26
    2, -2, 0, -9, -4, -4, 4, 1, -4,
    -- layer=1 filter=223 channel=27
    -4, 8, 0, 8, -1, 9, 3, 8, 0,
    -- layer=1 filter=223 channel=28
    -10, -11, -5, 9, 7, 0, 2, -8, 1,
    -- layer=1 filter=223 channel=29
    -1, 0, -10, -6, 7, -3, 0, 0, 7,
    -- layer=1 filter=223 channel=30
    -10, -3, -3, 5, -7, -11, -6, -7, 1,
    -- layer=1 filter=223 channel=31
    1, -6, 1, -8, -8, 5, 4, -7, -8,
    -- layer=1 filter=223 channel=32
    -2, -9, -8, 7, 1, -4, -3, -1, 4,
    -- layer=1 filter=223 channel=33
    0, -6, 6, -4, -5, 0, 7, -5, 3,
    -- layer=1 filter=223 channel=34
    1, -8, 4, -7, -3, 9, 4, 0, 9,
    -- layer=1 filter=223 channel=35
    -11, 8, -5, 9, -6, -5, -3, -3, 0,
    -- layer=1 filter=223 channel=36
    -6, 1, 0, -11, -2, 2, 5, 6, -5,
    -- layer=1 filter=223 channel=37
    1, 5, -6, -9, 0, 4, -5, -9, 6,
    -- layer=1 filter=223 channel=38
    -4, -11, 5, 6, -7, 0, 4, 4, 7,
    -- layer=1 filter=223 channel=39
    -11, 0, -7, 3, 11, -8, -8, -8, -9,
    -- layer=1 filter=223 channel=40
    9, 4, -7, -4, 8, 5, 10, 6, -5,
    -- layer=1 filter=223 channel=41
    7, -7, -3, -10, 2, 9, -8, -5, 1,
    -- layer=1 filter=223 channel=42
    -4, 4, -2, -5, -9, 0, -9, -9, -5,
    -- layer=1 filter=223 channel=43
    -1, -8, -11, -1, -10, -6, 0, -7, -2,
    -- layer=1 filter=223 channel=44
    -6, 4, -1, -10, 3, 11, -6, -2, 0,
    -- layer=1 filter=223 channel=45
    4, 2, 4, -5, -9, 3, 5, 0, -2,
    -- layer=1 filter=223 channel=46
    1, 8, -1, -9, 3, -6, 1, -9, -4,
    -- layer=1 filter=223 channel=47
    5, -1, -10, -3, 1, 7, 6, -8, 6,
    -- layer=1 filter=223 channel=48
    -8, -6, -8, 5, -5, 8, -12, -6, -13,
    -- layer=1 filter=223 channel=49
    -10, -7, 5, 6, -3, -12, -4, 1, 3,
    -- layer=1 filter=223 channel=50
    -3, -7, -1, -6, 6, 3, -10, 3, -6,
    -- layer=1 filter=223 channel=51
    1, 0, -6, -11, -11, -12, -9, -11, -3,
    -- layer=1 filter=223 channel=52
    -5, -7, -1, -3, -8, 0, 5, -8, -1,
    -- layer=1 filter=223 channel=53
    1, -6, -6, -7, -3, 5, 3, 7, -6,
    -- layer=1 filter=223 channel=54
    3, -10, 0, 0, 8, 0, 1, 0, -5,
    -- layer=1 filter=223 channel=55
    0, 7, -9, 7, 9, -10, 3, -3, 3,
    -- layer=1 filter=223 channel=56
    9, 0, 8, 0, 0, -7, 2, 0, -6,
    -- layer=1 filter=223 channel=57
    -9, 3, 7, 8, -6, 2, -6, -13, 7,
    -- layer=1 filter=223 channel=58
    4, 7, 4, -3, -9, -11, 0, 1, -10,
    -- layer=1 filter=223 channel=59
    -3, 1, -2, -6, 0, -2, 6, -5, -9,
    -- layer=1 filter=223 channel=60
    7, 0, -3, 9, 7, 7, 9, 7, 1,
    -- layer=1 filter=223 channel=61
    8, -10, -3, 0, -9, -4, 0, 9, 3,
    -- layer=1 filter=223 channel=62
    0, 5, 0, 0, 1, -7, -1, 6, 7,
    -- layer=1 filter=223 channel=63
    -7, -11, 2, -11, 0, 9, -6, -6, 10,
    -- layer=1 filter=223 channel=64
    7, -2, 7, -10, -12, -7, -2, -11, 1,
    -- layer=1 filter=223 channel=65
    6, 6, 0, 1, -5, 5, 0, -7, -12,
    -- layer=1 filter=223 channel=66
    7, 1, -8, -3, -8, -5, 6, -5, 8,
    -- layer=1 filter=223 channel=67
    10, 0, 5, 9, -2, -4, 9, 1, -2,
    -- layer=1 filter=223 channel=68
    5, -10, -2, 0, 0, -9, 4, -8, 0,
    -- layer=1 filter=223 channel=69
    1, 8, -9, -4, 3, -10, -1, 1, -6,
    -- layer=1 filter=223 channel=70
    0, 0, 7, -11, 7, 0, 0, 0, -1,
    -- layer=1 filter=223 channel=71
    -8, 3, 0, -10, -6, -9, -5, 0, 1,
    -- layer=1 filter=223 channel=72
    -1, 1, 5, 1, -1, 5, 1, 3, 4,
    -- layer=1 filter=223 channel=73
    3, 2, -8, -8, -4, 3, -6, 6, 0,
    -- layer=1 filter=223 channel=74
    -1, 5, -11, 6, -11, -7, 3, -8, -4,
    -- layer=1 filter=223 channel=75
    6, -8, 6, -11, -2, -10, 5, -8, -1,
    -- layer=1 filter=223 channel=76
    0, 0, 2, 3, -7, 0, -7, 3, 1,
    -- layer=1 filter=223 channel=77
    -9, 3, 0, -10, -1, -7, -12, -9, -2,
    -- layer=1 filter=223 channel=78
    0, 0, 5, -7, -9, -9, 4, -5, 10,
    -- layer=1 filter=223 channel=79
    4, 2, -10, 6, -7, -2, -8, -13, -2,
    -- layer=1 filter=223 channel=80
    -6, 6, 7, 3, -6, 3, 7, -7, 5,
    -- layer=1 filter=223 channel=81
    -8, -4, -2, 8, -6, 2, 0, -3, 5,
    -- layer=1 filter=223 channel=82
    -10, -9, 2, 0, 5, 0, 4, 7, 7,
    -- layer=1 filter=223 channel=83
    -7, 2, -3, 4, -5, -1, -5, -7, -5,
    -- layer=1 filter=223 channel=84
    -9, -1, -4, 5, 3, 0, 2, -1, 4,
    -- layer=1 filter=223 channel=85
    5, 8, -1, 0, 2, -1, 5, -2, 6,
    -- layer=1 filter=223 channel=86
    5, -11, 1, -9, -5, 8, 4, -5, 4,
    -- layer=1 filter=223 channel=87
    -6, -11, 5, 0, 9, 6, 7, -2, 2,
    -- layer=1 filter=223 channel=88
    1, 7, 3, 0, -1, 4, -2, 1, 6,
    -- layer=1 filter=223 channel=89
    4, -1, 0, 5, 0, -6, -6, -2, 2,
    -- layer=1 filter=223 channel=90
    5, -8, 3, -6, 3, 3, 2, -3, 0,
    -- layer=1 filter=223 channel=91
    2, -10, 6, 1, -11, -10, 1, -5, 3,
    -- layer=1 filter=223 channel=92
    -12, -2, 2, 2, -7, 8, 4, -3, -9,
    -- layer=1 filter=223 channel=93
    -1, 3, 6, -10, -3, 0, -8, -3, -8,
    -- layer=1 filter=223 channel=94
    -11, 3, -6, 0, 0, -10, -1, -7, -9,
    -- layer=1 filter=223 channel=95
    4, 6, 3, -4, 3, 7, -1, -8, -2,
    -- layer=1 filter=223 channel=96
    -8, -11, 1, -1, -2, -11, 5, -2, -11,
    -- layer=1 filter=223 channel=97
    -8, 0, 8, -12, -10, 8, -9, 0, -9,
    -- layer=1 filter=223 channel=98
    -4, 0, 4, -9, -1, -6, 3, 2, -9,
    -- layer=1 filter=223 channel=99
    -1, 6, 5, 5, 3, 1, 7, -10, 0,
    -- layer=1 filter=223 channel=100
    4, -11, -3, 4, 7, -1, -4, -9, 9,
    -- layer=1 filter=223 channel=101
    0, -8, -10, -1, -1, 6, -1, -2, -12,
    -- layer=1 filter=223 channel=102
    7, 5, 2, 7, -8, 4, 7, 0, 4,
    -- layer=1 filter=223 channel=103
    -5, 7, -2, 7, 8, 0, 4, -5, 7,
    -- layer=1 filter=223 channel=104
    -8, 0, -10, -4, -10, -8, -4, -5, -3,
    -- layer=1 filter=223 channel=105
    -4, -5, -9, -3, -11, 0, -7, 2, 7,
    -- layer=1 filter=223 channel=106
    -12, -6, -12, -9, -2, 0, -9, -10, 6,
    -- layer=1 filter=223 channel=107
    -9, 8, -1, 9, 9, -1, 1, 4, -1,
    -- layer=1 filter=223 channel=108
    4, -2, -5, -2, 4, -9, 2, 6, -3,
    -- layer=1 filter=223 channel=109
    6, -8, 8, -2, 9, -6, -8, -5, -7,
    -- layer=1 filter=223 channel=110
    6, -5, 7, 4, 4, 0, -6, -8, -9,
    -- layer=1 filter=223 channel=111
    9, 6, 1, 0, 0, 0, -8, 6, 6,
    -- layer=1 filter=223 channel=112
    2, 7, -8, -9, 0, -11, -12, -8, 5,
    -- layer=1 filter=223 channel=113
    -10, -3, -1, -7, -1, 0, 7, -2, 4,
    -- layer=1 filter=223 channel=114
    0, 9, -6, 6, -6, 5, -6, -6, 2,
    -- layer=1 filter=223 channel=115
    -7, -1, -9, 2, -6, -10, -2, 5, -12,
    -- layer=1 filter=223 channel=116
    -2, -5, -1, 9, 6, 3, 6, -5, -2,
    -- layer=1 filter=223 channel=117
    -5, -10, -9, -6, 9, -1, 3, 9, 4,
    -- layer=1 filter=223 channel=118
    -7, -6, 2, 3, -9, 4, 0, 0, 4,
    -- layer=1 filter=223 channel=119
    -7, -9, 7, -4, 0, -7, 3, 4, -7,
    -- layer=1 filter=223 channel=120
    4, -8, -8, 2, -4, -10, 2, -3, -8,
    -- layer=1 filter=223 channel=121
    5, -2, 0, 2, -7, 3, -3, -1, 8,
    -- layer=1 filter=223 channel=122
    -10, -9, -9, 3, 8, -6, 1, -6, 4,
    -- layer=1 filter=223 channel=123
    -8, -2, 0, -1, -11, 5, 8, 0, -9,
    -- layer=1 filter=223 channel=124
    0, 4, -2, -5, -11, -6, -8, 3, -11,
    -- layer=1 filter=223 channel=125
    6, 8, -2, 4, 5, -1, -7, 1, -11,
    -- layer=1 filter=223 channel=126
    0, -6, 7, -4, -1, 0, -3, -1, 3,
    -- layer=1 filter=223 channel=127
    -1, -5, -7, -1, -2, 0, -6, -10, 4,
    -- layer=1 filter=224 channel=0
    4, 7, -4, -10, 0, -6, 4, 6, 4,
    -- layer=1 filter=224 channel=1
    4, -11, 6, 4, 6, -9, 0, -3, -2,
    -- layer=1 filter=224 channel=2
    5, 5, 0, 2, -10, -7, 3, -10, 1,
    -- layer=1 filter=224 channel=3
    -7, 0, -6, -7, 8, 8, -3, -6, 2,
    -- layer=1 filter=224 channel=4
    -8, 2, 7, -1, 8, -4, -9, -9, 3,
    -- layer=1 filter=224 channel=5
    -3, -10, -4, 3, 3, 3, -8, -1, 1,
    -- layer=1 filter=224 channel=6
    -8, -8, 6, -4, -6, -10, 1, -4, -10,
    -- layer=1 filter=224 channel=7
    0, -6, 1, 6, 1, 0, -1, 8, -5,
    -- layer=1 filter=224 channel=8
    -5, 7, -5, 11, -5, -9, 5, 3, 0,
    -- layer=1 filter=224 channel=9
    8, 3, -9, 0, -1, 2, 5, 6, 0,
    -- layer=1 filter=224 channel=10
    -8, 8, -6, 10, -11, 7, 7, -5, -6,
    -- layer=1 filter=224 channel=11
    5, 9, 10, 0, -5, 4, 0, -8, 3,
    -- layer=1 filter=224 channel=12
    0, 8, 1, -7, 11, -10, 6, -5, -6,
    -- layer=1 filter=224 channel=13
    -7, 0, 1, 7, -3, -4, 1, 5, -2,
    -- layer=1 filter=224 channel=14
    -7, 7, 1, 4, 1, 1, -1, -6, -6,
    -- layer=1 filter=224 channel=15
    -2, -8, 5, -3, -1, 1, -7, -10, 4,
    -- layer=1 filter=224 channel=16
    7, 3, 1, -5, 7, -2, 0, 8, -4,
    -- layer=1 filter=224 channel=17
    -6, -4, -6, 7, -9, -10, -7, 1, 3,
    -- layer=1 filter=224 channel=18
    5, 1, -11, 5, 4, 2, -6, 2, -9,
    -- layer=1 filter=224 channel=19
    3, -1, 4, -2, 0, -8, -8, -11, -5,
    -- layer=1 filter=224 channel=20
    5, 0, -1, -3, -4, 0, -1, -1, -9,
    -- layer=1 filter=224 channel=21
    -10, 0, 0, 3, -1, -11, 1, -7, -1,
    -- layer=1 filter=224 channel=22
    -8, -12, -11, 2, -12, -1, 2, 0, -9,
    -- layer=1 filter=224 channel=23
    7, 3, 3, -10, -5, 4, 7, -3, 0,
    -- layer=1 filter=224 channel=24
    -4, 5, 2, -3, -4, 2, 7, -10, 1,
    -- layer=1 filter=224 channel=25
    10, -10, 6, -10, 6, 2, -2, -4, 2,
    -- layer=1 filter=224 channel=26
    -1, -1, 3, -1, 9, -10, -5, 2, -3,
    -- layer=1 filter=224 channel=27
    3, -5, -4, -2, 1, 4, -2, 0, 0,
    -- layer=1 filter=224 channel=28
    -5, 1, -4, 0, -12, 2, -9, -12, -7,
    -- layer=1 filter=224 channel=29
    1, -7, -9, -8, 1, 2, -4, 3, 2,
    -- layer=1 filter=224 channel=30
    -8, 4, 4, -3, -4, 1, -5, 4, 2,
    -- layer=1 filter=224 channel=31
    6, 4, -7, 2, 11, -1, 9, -1, 1,
    -- layer=1 filter=224 channel=32
    3, 2, -1, -6, 0, -12, -1, -6, -2,
    -- layer=1 filter=224 channel=33
    -8, -3, -10, -7, -2, -11, -2, 4, 5,
    -- layer=1 filter=224 channel=34
    -3, 0, 3, -4, -7, -8, 3, 0, 1,
    -- layer=1 filter=224 channel=35
    0, 4, 4, 2, 4, 0, 3, 7, -2,
    -- layer=1 filter=224 channel=36
    0, -3, -7, -3, -7, -2, 6, 1, -6,
    -- layer=1 filter=224 channel=37
    -11, -7, -5, 2, -11, 3, 1, 5, -4,
    -- layer=1 filter=224 channel=38
    6, -5, 5, 8, -4, -4, 4, 6, 0,
    -- layer=1 filter=224 channel=39
    -7, 4, -2, -5, -2, -12, -2, -9, 0,
    -- layer=1 filter=224 channel=40
    0, 3, -8, 6, 8, 0, 1, 2, -9,
    -- layer=1 filter=224 channel=41
    -11, -1, 3, 3, 4, 4, 5, 7, 1,
    -- layer=1 filter=224 channel=42
    -1, 8, -3, -2, 2, -5, -1, 8, -9,
    -- layer=1 filter=224 channel=43
    -5, -7, 0, 3, 4, 0, -1, 1, 0,
    -- layer=1 filter=224 channel=44
    -2, 0, 6, 6, 0, -11, -5, 9, -9,
    -- layer=1 filter=224 channel=45
    6, 5, -9, 2, -8, -5, 0, 5, -2,
    -- layer=1 filter=224 channel=46
    -8, -3, -10, -7, 7, 9, 3, 7, 1,
    -- layer=1 filter=224 channel=47
    -4, 11, -8, -11, -3, 10, -3, 0, 0,
    -- layer=1 filter=224 channel=48
    7, -5, 0, 1, 3, 0, -3, -2, -7,
    -- layer=1 filter=224 channel=49
    -4, -8, -3, 6, 8, 0, 2, -6, -7,
    -- layer=1 filter=224 channel=50
    7, 0, -1, 6, -9, -8, 2, -6, -9,
    -- layer=1 filter=224 channel=51
    0, -8, 7, -8, 6, 3, -9, 6, -9,
    -- layer=1 filter=224 channel=52
    6, -6, -4, -3, 7, -6, 3, 8, 9,
    -- layer=1 filter=224 channel=53
    -10, -6, 0, -8, 0, 2, -1, 0, -7,
    -- layer=1 filter=224 channel=54
    -4, 4, 2, 5, -1, -4, -11, -3, 3,
    -- layer=1 filter=224 channel=55
    0, 4, -6, 1, 4, 8, -9, -10, 0,
    -- layer=1 filter=224 channel=56
    6, 5, 1, 7, -11, -10, -1, 4, -7,
    -- layer=1 filter=224 channel=57
    -10, 3, 2, 1, -5, 3, -6, -2, 3,
    -- layer=1 filter=224 channel=58
    5, 7, 5, -1, -11, -8, -4, -8, 3,
    -- layer=1 filter=224 channel=59
    5, -2, 0, -5, 8, 8, -3, -12, 0,
    -- layer=1 filter=224 channel=60
    5, 0, 11, -5, -8, 0, -5, 7, -9,
    -- layer=1 filter=224 channel=61
    6, 8, 3, -11, 2, 3, 1, -1, -5,
    -- layer=1 filter=224 channel=62
    12, -11, 2, -8, 1, 8, -11, 7, 4,
    -- layer=1 filter=224 channel=63
    -12, -10, 2, 2, 7, -2, -3, 2, 8,
    -- layer=1 filter=224 channel=64
    -7, -9, 5, -5, 8, -3, -2, -2, -9,
    -- layer=1 filter=224 channel=65
    -3, -1, 5, 5, 6, -9, 5, 3, -2,
    -- layer=1 filter=224 channel=66
    -1, -9, -11, -1, -5, 1, -8, -10, -1,
    -- layer=1 filter=224 channel=67
    0, -8, 0, 4, -6, -3, 4, 2, 6,
    -- layer=1 filter=224 channel=68
    -6, -8, -9, -1, -12, -8, -7, 3, 4,
    -- layer=1 filter=224 channel=69
    2, -1, -2, -4, 0, -8, -11, 0, -3,
    -- layer=1 filter=224 channel=70
    -7, -2, -9, -4, -8, -9, -2, -3, -4,
    -- layer=1 filter=224 channel=71
    -11, 6, 0, 8, -10, 0, 2, 0, -6,
    -- layer=1 filter=224 channel=72
    -4, -12, -12, 3, 7, -4, -10, 4, 2,
    -- layer=1 filter=224 channel=73
    -6, -1, 5, -5, -8, 8, -7, -10, 1,
    -- layer=1 filter=224 channel=74
    1, 5, 4, 3, -3, 3, 7, 2, 1,
    -- layer=1 filter=224 channel=75
    -3, -1, -9, -1, -6, 9, -9, 7, 1,
    -- layer=1 filter=224 channel=76
    4, 0, 1, -2, 1, -11, -4, -3, -7,
    -- layer=1 filter=224 channel=77
    -5, 6, 3, 2, 7, 7, -8, -4, -8,
    -- layer=1 filter=224 channel=78
    -10, -10, 0, 0, 2, -12, -8, 7, -2,
    -- layer=1 filter=224 channel=79
    -3, -6, -2, -8, -5, 7, -12, 2, -1,
    -- layer=1 filter=224 channel=80
    3, -1, 0, 9, 8, 0, 7, -11, 0,
    -- layer=1 filter=224 channel=81
    -11, -3, -10, 0, -7, -6, 9, -7, 4,
    -- layer=1 filter=224 channel=82
    -2, 3, -7, -7, -8, -9, -5, 8, 8,
    -- layer=1 filter=224 channel=83
    3, 3, -12, 0, -5, 0, -3, 2, -4,
    -- layer=1 filter=224 channel=84
    -11, -2, -2, -1, -4, -2, 0, 2, -10,
    -- layer=1 filter=224 channel=85
    -10, -2, -1, -5, -1, -7, -6, 1, -10,
    -- layer=1 filter=224 channel=86
    -4, 2, 7, -3, 1, 5, 3, -7, -9,
    -- layer=1 filter=224 channel=87
    -1, 5, 1, -5, -1, -6, 3, 0, 2,
    -- layer=1 filter=224 channel=88
    4, 1, 7, 4, -5, 8, -6, -3, 0,
    -- layer=1 filter=224 channel=89
    5, 8, 1, 1, 7, 6, 0, -7, -4,
    -- layer=1 filter=224 channel=90
    -9, 3, -3, -5, 9, -6, -9, 6, -10,
    -- layer=1 filter=224 channel=91
    6, 5, -5, -7, -1, 3, 1, -9, 4,
    -- layer=1 filter=224 channel=92
    1, 3, -12, -1, -1, -1, -7, 7, 2,
    -- layer=1 filter=224 channel=93
    -12, -12, 6, 4, -4, -3, 7, 1, -2,
    -- layer=1 filter=224 channel=94
    -7, -8, 0, 6, -5, 5, -6, 2, -9,
    -- layer=1 filter=224 channel=95
    2, -2, -1, -5, -3, -9, -9, 5, 6,
    -- layer=1 filter=224 channel=96
    -8, -4, -11, -8, 1, -6, -5, -5, -2,
    -- layer=1 filter=224 channel=97
    -11, -11, 0, -10, 5, -5, -9, -5, 8,
    -- layer=1 filter=224 channel=98
    4, 4, 6, 0, 6, -5, -7, 3, -2,
    -- layer=1 filter=224 channel=99
    -11, -6, 0, -11, -8, -1, 3, -4, -2,
    -- layer=1 filter=224 channel=100
    -8, -1, -9, -9, 2, -1, -3, 2, -9,
    -- layer=1 filter=224 channel=101
    -6, 3, 6, -11, 6, -12, 3, 0, 4,
    -- layer=1 filter=224 channel=102
    -3, 5, -1, -5, -4, 6, 8, -9, -5,
    -- layer=1 filter=224 channel=103
    10, 0, 4, -2, -6, 2, 8, 9, 5,
    -- layer=1 filter=224 channel=104
    -7, 8, -2, 7, -6, -4, -2, 7, -8,
    -- layer=1 filter=224 channel=105
    0, -6, -8, 8, -4, -10, 7, -7, 4,
    -- layer=1 filter=224 channel=106
    -10, -1, -10, -12, 0, -3, 6, 0, 0,
    -- layer=1 filter=224 channel=107
    1, 0, 8, 6, 1, -6, 2, -6, -4,
    -- layer=1 filter=224 channel=108
    -2, 3, -11, 4, 11, -11, -4, -3, -4,
    -- layer=1 filter=224 channel=109
    -8, 8, -9, 4, 1, 9, -10, -6, -11,
    -- layer=1 filter=224 channel=110
    4, 6, -8, -1, 3, 4, -2, -6, 6,
    -- layer=1 filter=224 channel=111
    7, -10, -1, 5, 7, -8, 3, 0, -9,
    -- layer=1 filter=224 channel=112
    -5, -7, 7, -3, -3, -6, -9, 8, 0,
    -- layer=1 filter=224 channel=113
    4, 2, -9, -8, 5, -4, -4, -12, -7,
    -- layer=1 filter=224 channel=114
    3, 11, 0, -7, -3, 6, 0, -5, -8,
    -- layer=1 filter=224 channel=115
    -1, 4, 7, 1, 7, 4, -1, -4, -8,
    -- layer=1 filter=224 channel=116
    -1, 9, -5, 3, -1, 4, -7, 9, -2,
    -- layer=1 filter=224 channel=117
    -7, 7, 7, 7, 0, -6, -6, -4, -10,
    -- layer=1 filter=224 channel=118
    -4, -2, -6, -12, 1, 8, -4, -4, 3,
    -- layer=1 filter=224 channel=119
    -9, 0, -1, -5, -11, -5, -5, -5, -5,
    -- layer=1 filter=224 channel=120
    -4, -1, -8, 3, 1, 2, 0, 6, -9,
    -- layer=1 filter=224 channel=121
    0, -6, -1, 1, -5, 4, -9, -9, 9,
    -- layer=1 filter=224 channel=122
    4, -7, -4, 4, 9, -10, 0, -6, 8,
    -- layer=1 filter=224 channel=123
    -4, 3, 5, 9, -3, -6, -3, -10, 0,
    -- layer=1 filter=224 channel=124
    -2, -6, -7, 8, 3, -9, -10, -8, 3,
    -- layer=1 filter=224 channel=125
    3, 5, -9, -7, 7, 2, 7, -8, -4,
    -- layer=1 filter=224 channel=126
    -7, -12, -1, 1, -2, -3, -9, 1, 1,
    -- layer=1 filter=224 channel=127
    -2, -12, 0, 6, -5, 8, -8, -3, -3,
    -- layer=1 filter=225 channel=0
    -12, -8, 11, 4, -6, -4, -19, -1, -10,
    -- layer=1 filter=225 channel=1
    27, 13, 13, -26, 13, 0, -6, 2, -24,
    -- layer=1 filter=225 channel=2
    -12, -14, -9, 1, 6, 8, 32, -5, 6,
    -- layer=1 filter=225 channel=3
    6, -7, -4, -10, 3, -4, 3, -6, 7,
    -- layer=1 filter=225 channel=4
    -2, -1, 14, 8, 1, -3, -8, 5, 0,
    -- layer=1 filter=225 channel=5
    -11, 3, -5, -11, 40, 9, 11, -6, -6,
    -- layer=1 filter=225 channel=6
    21, 25, 18, 15, 0, -3, -25, -36, -51,
    -- layer=1 filter=225 channel=7
    -30, -36, -1, -29, -64, -31, -13, -25, 3,
    -- layer=1 filter=225 channel=8
    19, 9, 7, -32, -17, -21, 5, 0, 0,
    -- layer=1 filter=225 channel=9
    -20, -12, 8, 6, -6, 4, -32, -9, -40,
    -- layer=1 filter=225 channel=10
    -16, -34, 5, -25, -22, -16, -12, -29, 5,
    -- layer=1 filter=225 channel=11
    -22, -20, -11, 11, 2, 15, 4, 24, 10,
    -- layer=1 filter=225 channel=12
    -31, 20, 4, 52, 14, -10, -8, 11, -16,
    -- layer=1 filter=225 channel=13
    22, 32, 19, 2, 7, -11, -17, -30, -43,
    -- layer=1 filter=225 channel=14
    -20, -27, -18, -20, -13, -27, 25, -18, 0,
    -- layer=1 filter=225 channel=15
    -11, 31, -26, -10, 9, -45, 35, -22, -8,
    -- layer=1 filter=225 channel=16
    10, 11, 13, -25, 26, 0, -2, 0, 8,
    -- layer=1 filter=225 channel=17
    23, 14, 12, -2, 3, -19, -31, -30, -16,
    -- layer=1 filter=225 channel=18
    -40, -36, -16, 35, 40, 21, 26, 26, 13,
    -- layer=1 filter=225 channel=19
    15, 36, 15, 81, 59, 47, 35, 44, 14,
    -- layer=1 filter=225 channel=20
    41, 30, 25, 6, 0, 0, -34, -30, -32,
    -- layer=1 filter=225 channel=21
    14, 9, 29, -20, -4, -11, -33, -40, -39,
    -- layer=1 filter=225 channel=22
    49, 36, 10, -6, -9, -12, -33, -42, -31,
    -- layer=1 filter=225 channel=23
    4, 29, 3, -2, -26, -11, 8, 6, 20,
    -- layer=1 filter=225 channel=24
    18, 11, 20, -19, -10, -8, -1, -4, -5,
    -- layer=1 filter=225 channel=25
    -7, 6, 36, -48, -17, -12, -11, -13, 6,
    -- layer=1 filter=225 channel=26
    11, 35, 9, -28, -23, -10, 0, -14, -26,
    -- layer=1 filter=225 channel=27
    -19, -5, 6, -7, 7, 9, -3, -18, -18,
    -- layer=1 filter=225 channel=28
    4, -9, 30, -39, -50, -41, -24, -43, -13,
    -- layer=1 filter=225 channel=29
    10, 7, 13, -10, 6, 2, -6, -6, -16,
    -- layer=1 filter=225 channel=30
    -35, -39, 7, 24, 40, 24, 24, 34, 3,
    -- layer=1 filter=225 channel=31
    20, 22, 8, 34, 22, 17, -2, -6, -8,
    -- layer=1 filter=225 channel=32
    -19, -1, 7, 18, 21, -6, 23, -7, 0,
    -- layer=1 filter=225 channel=33
    24, 9, 3, -13, 1, 0, -23, -24, -32,
    -- layer=1 filter=225 channel=34
    2, 30, 5, 4, -6, -9, -25, -26, -28,
    -- layer=1 filter=225 channel=35
    -20, 1, -20, -1, -21, -21, 4, -4, -4,
    -- layer=1 filter=225 channel=36
    -24, -29, -9, 4, 24, 14, 8, 27, 4,
    -- layer=1 filter=225 channel=37
    3, 13, 2, 19, 73, 28, 17, 15, 3,
    -- layer=1 filter=225 channel=38
    40, 29, 25, 24, 7, -3, -22, -39, -19,
    -- layer=1 filter=225 channel=39
    5, 10, 9, -13, -9, -6, -9, 2, 7,
    -- layer=1 filter=225 channel=40
    35, 12, 16, 9, 10, -1, -16, -9, -35,
    -- layer=1 filter=225 channel=41
    -56, -56, -6, 7, -11, 11, -5, -8, -35,
    -- layer=1 filter=225 channel=42
    -25, 17, -12, -13, -3, -4, 7, 22, 0,
    -- layer=1 filter=225 channel=43
    24, 0, 4, -44, -34, -24, -14, 8, 13,
    -- layer=1 filter=225 channel=44
    -21, 6, -3, -9, -8, -22, -15, -30, -15,
    -- layer=1 filter=225 channel=45
    31, 19, -9, -14, 1, -14, -6, -15, -15,
    -- layer=1 filter=225 channel=46
    20, 41, 15, 67, 60, 37, 15, 9, 26,
    -- layer=1 filter=225 channel=47
    3, 25, 19, 38, 22, 13, 22, -13, 0,
    -- layer=1 filter=225 channel=48
    22, 25, 16, 1, -13, 0, -15, -27, -37,
    -- layer=1 filter=225 channel=49
    9, 16, 19, 17, 6, 7, -9, -28, -23,
    -- layer=1 filter=225 channel=50
    8, 0, -3, -3, -11, 2, -18, -11, -20,
    -- layer=1 filter=225 channel=51
    27, 20, 19, 11, -6, -5, -12, -41, -22,
    -- layer=1 filter=225 channel=52
    -15, 2, 3, -6, 0, 2, 6, 11, 2,
    -- layer=1 filter=225 channel=53
    -1, 16, 10, -3, -1, 9, -1, 4, 20,
    -- layer=1 filter=225 channel=54
    -12, -9, 1, -13, 32, 5, -5, 4, -1,
    -- layer=1 filter=225 channel=55
    -13, -18, -16, -2, -3, -2, 15, 26, 12,
    -- layer=1 filter=225 channel=56
    0, 8, 5, -5, -7, 6, -2, -7, -4,
    -- layer=1 filter=225 channel=57
    8, -6, 8, 1, -8, -10, -22, -19, -6,
    -- layer=1 filter=225 channel=58
    -1, 17, 4, 10, -17, 9, 24, -10, 19,
    -- layer=1 filter=225 channel=59
    -6, -8, -20, -17, -12, -11, -8, 9, -5,
    -- layer=1 filter=225 channel=60
    10, -4, 4, -6, -1, -12, 8, -8, -2,
    -- layer=1 filter=225 channel=61
    -7, 2, -7, 8, -12, 0, 7, 8, 0,
    -- layer=1 filter=225 channel=62
    21, 10, 11, -40, 0, -10, -9, 3, -8,
    -- layer=1 filter=225 channel=63
    -37, -22, -17, 7, 20, 14, 2, 1, -11,
    -- layer=1 filter=225 channel=64
    13, 3, 5, -2, 8, 5, -22, -28, -32,
    -- layer=1 filter=225 channel=65
    28, 20, 7, -12, -11, -6, -41, -35, -26,
    -- layer=1 filter=225 channel=66
    1, -5, -3, 1, 6, 10, -11, -2, 4,
    -- layer=1 filter=225 channel=67
    22, 19, 16, 18, 18, 16, -21, -19, -23,
    -- layer=1 filter=225 channel=68
    -19, 4, 6, -24, -18, -9, -18, -14, -12,
    -- layer=1 filter=225 channel=69
    2, 10, -28, -36, -6, -36, 21, -2, 14,
    -- layer=1 filter=225 channel=70
    23, 14, -1, 25, 29, 25, -6, -17, -7,
    -- layer=1 filter=225 channel=71
    21, 5, 18, -17, -9, -4, -16, -13, -8,
    -- layer=1 filter=225 channel=72
    -42, -4, 22, 48, 29, 28, 11, 26, 5,
    -- layer=1 filter=225 channel=73
    -7, -1, -9, 8, -6, 14, -4, -8, -12,
    -- layer=1 filter=225 channel=74
    14, -6, 17, 11, 11, 34, -6, -8, -12,
    -- layer=1 filter=225 channel=75
    -74, -32, -8, 40, 28, 4, 31, 26, 21,
    -- layer=1 filter=225 channel=76
    -33, -17, 12, 11, 10, 10, 13, -21, -3,
    -- layer=1 filter=225 channel=77
    25, 22, 19, -13, -7, -5, -22, -20, -34,
    -- layer=1 filter=225 channel=78
    -10, 9, -4, 7, 4, -8, -3, -1, 8,
    -- layer=1 filter=225 channel=79
    29, 9, 3, -34, -6, -5, -18, 3, 6,
    -- layer=1 filter=225 channel=80
    -9, -8, 2, 5, -3, -1, 7, 15, 22,
    -- layer=1 filter=225 channel=81
    31, 28, 14, -47, -47, -34, -4, 1, 7,
    -- layer=1 filter=225 channel=82
    23, 33, 24, 8, 0, 1, -33, -45, -25,
    -- layer=1 filter=225 channel=83
    23, 29, -7, -2, -25, -14, 7, -24, -18,
    -- layer=1 filter=225 channel=84
    -28, -21, 7, 35, 47, 33, 16, 10, -17,
    -- layer=1 filter=225 channel=85
    7, 19, 6, 32, -12, 9, 10, 0, -7,
    -- layer=1 filter=225 channel=86
    6, -1, -2, 9, 14, 18, 6, -2, -4,
    -- layer=1 filter=225 channel=87
    9, 44, 0, 56, 36, 11, -1, 24, 1,
    -- layer=1 filter=225 channel=88
    7, 11, -1, -13, 2, -3, -20, -34, -28,
    -- layer=1 filter=225 channel=89
    15, 24, 11, 2, -12, -6, -23, -26, -43,
    -- layer=1 filter=225 channel=90
    -8, 24, -5, -52, -36, -45, -5, -9, -19,
    -- layer=1 filter=225 channel=91
    26, 25, 10, 19, 24, -2, -18, -30, -27,
    -- layer=1 filter=225 channel=92
    -47, -16, -25, -29, -8, -30, 15, 8, -4,
    -- layer=1 filter=225 channel=93
    10, 23, 20, 0, -19, -17, -18, -30, -10,
    -- layer=1 filter=225 channel=94
    2, -16, 0, 3, -3, 8, 0, -17, 2,
    -- layer=1 filter=225 channel=95
    -24, -32, 18, 38, 39, 24, 28, 13, 3,
    -- layer=1 filter=225 channel=96
    -7, 13, 0, 4, -10, 0, 5, -6, -6,
    -- layer=1 filter=225 channel=97
    7, 17, -2, -16, 1, -14, -23, -19, -12,
    -- layer=1 filter=225 channel=98
    10, 0, 8, -45, -29, -23, -29, -3, 9,
    -- layer=1 filter=225 channel=99
    24, -18, 21, -8, -30, -5, -14, -27, 13,
    -- layer=1 filter=225 channel=100
    -40, -25, -16, 22, 29, 5, 13, -3, -1,
    -- layer=1 filter=225 channel=101
    35, 29, 10, 18, 19, 6, -22, -34, -37,
    -- layer=1 filter=225 channel=102
    -2, 6, -11, 0, 13, 6, -12, -26, -14,
    -- layer=1 filter=225 channel=103
    -10, -3, -6, 26, 29, 34, 2, 23, 8,
    -- layer=1 filter=225 channel=104
    -3, 8, -6, 29, 0, 6, 39, 2, 0,
    -- layer=1 filter=225 channel=105
    5, 5, 9, 0, -9, -5, -1, -16, 0,
    -- layer=1 filter=225 channel=106
    22, 38, 5, 25, 15, 7, -18, -29, -25,
    -- layer=1 filter=225 channel=107
    -20, -21, -22, -6, -1, 6, 11, 5, -5,
    -- layer=1 filter=225 channel=108
    -9, 6, -8, -26, -42, -53, 11, -10, 0,
    -- layer=1 filter=225 channel=109
    0, 2, -2, 7, -4, 9, -5, -10, -8,
    -- layer=1 filter=225 channel=110
    -3, -3, 5, 9, -1, 2, -17, -16, -9,
    -- layer=1 filter=225 channel=111
    -26, -46, -11, 21, 30, 31, 15, -3, -3,
    -- layer=1 filter=225 channel=112
    8, 0, 11, 36, 47, 36, 19, -12, 12,
    -- layer=1 filter=225 channel=113
    44, 30, 32, 8, 23, -5, -19, -21, -32,
    -- layer=1 filter=225 channel=114
    -8, -7, -29, -45, -29, -38, 18, 10, 11,
    -- layer=1 filter=225 channel=115
    14, 5, 9, 6, 0, 0, -10, -16, 0,
    -- layer=1 filter=225 channel=116
    5, 3, 2, 3, -12, 6, -1, -6, -1,
    -- layer=1 filter=225 channel=117
    28, -5, 13, 65, 61, 58, 42, 5, 26,
    -- layer=1 filter=225 channel=118
    -26, -32, 1, 30, 29, 39, 16, 11, -11,
    -- layer=1 filter=225 channel=119
    -30, -7, 4, -3, -4, -18, 7, -24, -15,
    -- layer=1 filter=225 channel=120
    19, 11, 18, -25, -3, -15, -16, -28, -28,
    -- layer=1 filter=225 channel=121
    -25, -16, -12, 23, 55, 29, 19, 23, 14,
    -- layer=1 filter=225 channel=122
    3, 6, 9, 4, -5, 0, 8, -2, 8,
    -- layer=1 filter=225 channel=123
    -46, -21, -39, 11, 22, 19, 15, 22, 1,
    -- layer=1 filter=225 channel=124
    11, 10, -1, -4, -10, 8, -4, -2, 4,
    -- layer=1 filter=225 channel=125
    29, 18, -1, 21, 32, 22, -9, -18, -31,
    -- layer=1 filter=225 channel=126
    39, 19, 8, 8, 9, 18, -11, 18, -1,
    -- layer=1 filter=225 channel=127
    -28, -42, 8, 31, 48, 36, 12, 29, 1,
    -- layer=1 filter=226 channel=0
    -20, -22, -8, -12, 1, -12, -2, -3, 0,
    -- layer=1 filter=226 channel=1
    -23, -13, -27, -3, -12, -1, 7, 15, 25,
    -- layer=1 filter=226 channel=2
    0, 27, -6, 10, 33, 29, 9, 15, 8,
    -- layer=1 filter=226 channel=3
    -3, -4, -3, 5, -12, -10, 5, -15, 2,
    -- layer=1 filter=226 channel=4
    0, -3, 3, 10, 0, -8, 1, 7, -1,
    -- layer=1 filter=226 channel=5
    -44, -3, -12, -8, -21, 11, 1, 5, 34,
    -- layer=1 filter=226 channel=6
    -16, -8, -6, -12, -23, -22, -32, -33, 3,
    -- layer=1 filter=226 channel=7
    -23, -3, 17, 9, -13, 19, -31, -30, -28,
    -- layer=1 filter=226 channel=8
    -22, -20, -26, -16, -28, -10, -1, 32, 28,
    -- layer=1 filter=226 channel=9
    -24, 20, -24, 0, -31, 12, -25, -10, -86,
    -- layer=1 filter=226 channel=10
    1, 10, 16, 13, -13, 24, -48, -35, -38,
    -- layer=1 filter=226 channel=11
    5, 16, 17, -6, 5, 15, 4, 5, 10,
    -- layer=1 filter=226 channel=12
    -71, -66, 7, -81, -22, 11, -37, -36, -25,
    -- layer=1 filter=226 channel=13
    22, 24, -5, 20, 0, 12, 8, 3, 19,
    -- layer=1 filter=226 channel=14
    -18, -4, 34, 7, -44, 27, -14, -33, -9,
    -- layer=1 filter=226 channel=15
    -29, -6, -28, -21, -15, -32, -5, -36, 12,
    -- layer=1 filter=226 channel=16
    -37, -14, -19, -8, -7, -3, 2, 11, 21,
    -- layer=1 filter=226 channel=17
    0, 0, 1, 12, 4, 26, 17, 33, 8,
    -- layer=1 filter=226 channel=18
    8, -3, -7, 10, 11, 18, -9, -13, 34,
    -- layer=1 filter=226 channel=19
    -34, -31, -65, -40, -71, -44, -26, -40, -85,
    -- layer=1 filter=226 channel=20
    26, 18, 2, 14, 12, 25, 24, 23, 14,
    -- layer=1 filter=226 channel=21
    10, -5, 1, 23, 6, -11, 2, 12, -12,
    -- layer=1 filter=226 channel=22
    27, 25, 15, 21, 16, 21, 16, 24, 34,
    -- layer=1 filter=226 channel=23
    0, -8, 0, -6, 24, 10, 0, -14, 17,
    -- layer=1 filter=226 channel=24
    0, -2, -25, 5, -9, 15, 18, 26, 1,
    -- layer=1 filter=226 channel=25
    7, 3, 5, 14, -11, 6, -27, -15, -39,
    -- layer=1 filter=226 channel=26
    34, 25, 18, 32, 27, 39, 35, 19, 10,
    -- layer=1 filter=226 channel=27
    -62, -55, -65, -33, -30, -34, -47, -23, -51,
    -- layer=1 filter=226 channel=28
    -19, 5, 6, 11, -9, 23, -14, -5, -36,
    -- layer=1 filter=226 channel=29
    -19, -39, -41, -23, -22, -11, -17, -13, -22,
    -- layer=1 filter=226 channel=30
    -60, -62, -64, -59, -88, -58, -57, -64, -64,
    -- layer=1 filter=226 channel=31
    -6, -7, 14, 2, -6, 4, -12, -7, 10,
    -- layer=1 filter=226 channel=32
    21, 25, 16, -4, 6, -3, 6, -36, -2,
    -- layer=1 filter=226 channel=33
    -35, -28, -40, -5, -27, -38, 3, -11, -13,
    -- layer=1 filter=226 channel=34
    -37, -63, -33, -39, -40, -36, -38, -50, -20,
    -- layer=1 filter=226 channel=35
    -5, -14, 4, -12, 4, 0, 2, -12, -9,
    -- layer=1 filter=226 channel=36
    6, -2, 22, 7, 5, 4, -5, 21, 13,
    -- layer=1 filter=226 channel=37
    -54, -22, -34, -14, -28, 1, 5, 1, 7,
    -- layer=1 filter=226 channel=38
    5, 9, -2, 25, 6, -4, 13, 2, -6,
    -- layer=1 filter=226 channel=39
    -19, -15, -25, -15, -23, -4, 5, -15, -2,
    -- layer=1 filter=226 channel=40
    -19, -18, 10, -19, -32, -3, -33, -40, 0,
    -- layer=1 filter=226 channel=41
    -7, 33, 21, 26, -34, -25, -7, -30, -71,
    -- layer=1 filter=226 channel=42
    -2, 15, 4, 18, 8, 31, 6, 5, 13,
    -- layer=1 filter=226 channel=43
    -43, -20, -45, -14, -30, -15, -15, 0, -6,
    -- layer=1 filter=226 channel=44
    13, 30, 14, 26, -2, 7, 21, -22, 17,
    -- layer=1 filter=226 channel=45
    0, 9, -10, 9, -5, -10, 14, 7, 11,
    -- layer=1 filter=226 channel=46
    -44, -45, -26, -54, -49, -32, -41, -48, -20,
    -- layer=1 filter=226 channel=47
    12, 15, -6, 1, -14, 14, -21, -36, -26,
    -- layer=1 filter=226 channel=48
    -1, -3, -18, 5, -5, -6, 14, 1, -24,
    -- layer=1 filter=226 channel=49
    19, 11, -17, 6, 7, 2, 4, -4, -10,
    -- layer=1 filter=226 channel=50
    2, 14, 6, 7, -1, -7, 4, 8, 18,
    -- layer=1 filter=226 channel=51
    0, -4, -8, -1, -8, 4, -12, -20, -36,
    -- layer=1 filter=226 channel=52
    1, 10, 3, 3, 5, 0, -6, -5, -9,
    -- layer=1 filter=226 channel=53
    4, -2, -8, 0, 4, 9, -7, 1, 0,
    -- layer=1 filter=226 channel=54
    7, -30, -23, 11, -25, 6, -20, -45, -60,
    -- layer=1 filter=226 channel=55
    16, 10, 35, 9, 18, 19, 15, 21, 1,
    -- layer=1 filter=226 channel=56
    -3, 11, -3, 8, 5, 1, -1, 0, -5,
    -- layer=1 filter=226 channel=57
    4, 18, 26, 19, -16, 38, -23, -24, -21,
    -- layer=1 filter=226 channel=58
    -5, 10, 14, 6, -22, 39, -40, -24, -38,
    -- layer=1 filter=226 channel=59
    9, 7, 16, 9, 6, -2, 8, 1, 0,
    -- layer=1 filter=226 channel=60
    -11, -16, -8, -6, -5, -24, -9, -6, -18,
    -- layer=1 filter=226 channel=61
    2, 3, -1, -4, 7, -9, -9, 0, 1,
    -- layer=1 filter=226 channel=62
    -24, -28, -39, -10, -32, 21, -9, 29, 1,
    -- layer=1 filter=226 channel=63
    -13, -13, 13, -13, -9, -8, -11, -2, 0,
    -- layer=1 filter=226 channel=64
    0, -10, -14, 13, 7, 4, -6, 15, -1,
    -- layer=1 filter=226 channel=65
    0, -18, -28, 9, -1, -23, 14, -9, -18,
    -- layer=1 filter=226 channel=66
    0, -12, -13, -8, -6, -7, 13, 8, -3,
    -- layer=1 filter=226 channel=67
    29, 12, 9, -2, -12, -20, -21, -21, -33,
    -- layer=1 filter=226 channel=68
    4, 18, -2, 7, 13, 8, 14, -1, 10,
    -- layer=1 filter=226 channel=69
    -19, 2, 8, 12, -8, 27, 18, -1, 8,
    -- layer=1 filter=226 channel=70
    -55, -55, -38, -26, -40, -53, -48, -23, -26,
    -- layer=1 filter=226 channel=71
    -18, -25, -14, 18, -5, -1, 2, 2, -10,
    -- layer=1 filter=226 channel=72
    -45, -36, -30, -49, -57, -28, -28, -53, -44,
    -- layer=1 filter=226 channel=73
    -4, 4, 5, 2, 10, -13, 2, 1, -3,
    -- layer=1 filter=226 channel=74
    -45, -34, -12, -26, -7, -51, -32, -32, 18,
    -- layer=1 filter=226 channel=75
    -77, -66, 0, -40, -60, -2, -19, -66, -3,
    -- layer=1 filter=226 channel=76
    -11, -6, -16, -12, -25, -19, -7, -25, -13,
    -- layer=1 filter=226 channel=77
    4, -11, -23, 19, 1, -13, 27, 5, -9,
    -- layer=1 filter=226 channel=78
    24, -14, 6, 14, -3, 12, 15, -5, 11,
    -- layer=1 filter=226 channel=79
    -9, -13, -15, 13, -2, 26, 20, 30, 7,
    -- layer=1 filter=226 channel=80
    0, -7, 0, -2, 0, -5, -10, -4, -7,
    -- layer=1 filter=226 channel=81
    -19, -23, -14, 9, -1, -1, 19, 19, 4,
    -- layer=1 filter=226 channel=82
    3, -15, -28, 7, -6, -18, 7, -12, -10,
    -- layer=1 filter=226 channel=83
    -3, -1, -2, -4, -39, 12, 25, -5, 4,
    -- layer=1 filter=226 channel=84
    -38, -38, -45, -46, -32, -29, -29, -42, 15,
    -- layer=1 filter=226 channel=85
    17, -2, 13, 15, -11, 45, -12, -25, -10,
    -- layer=1 filter=226 channel=86
    16, 22, 27, 12, 17, 25, 15, 32, 36,
    -- layer=1 filter=226 channel=87
    -28, -23, -50, -3, -62, -17, -28, -34, -78,
    -- layer=1 filter=226 channel=88
    15, 1, 5, 0, 17, -13, 15, 0, 0,
    -- layer=1 filter=226 channel=89
    3, -25, -15, -3, 9, -31, 23, -11, 3,
    -- layer=1 filter=226 channel=90
    12, 29, 26, 21, 0, 37, 0, 6, -5,
    -- layer=1 filter=226 channel=91
    29, 14, 7, 9, 1, 1, 14, 1, 11,
    -- layer=1 filter=226 channel=92
    35, -18, 23, 18, -33, -16, -20, -86, -55,
    -- layer=1 filter=226 channel=93
    0, -10, -13, 15, 0, -4, 7, 3, 8,
    -- layer=1 filter=226 channel=94
    -9, -14, -7, -12, 3, 0, 2, 12, 15,
    -- layer=1 filter=226 channel=95
    -50, -97, -40, -58, -40, -56, -49, -63, -1,
    -- layer=1 filter=226 channel=96
    0, 10, 7, 8, 0, -2, -7, 10, -6,
    -- layer=1 filter=226 channel=97
    -2, -15, -19, 2, -2, 5, 11, 17, 11,
    -- layer=1 filter=226 channel=98
    2, 3, -20, 7, -31, 12, 10, 18, -3,
    -- layer=1 filter=226 channel=99
    -14, -8, -14, 3, 1, -4, -45, -9, -64,
    -- layer=1 filter=226 channel=100
    -14, -7, 3, -10, -1, -9, 10, -10, 8,
    -- layer=1 filter=226 channel=101
    12, 1, 0, -1, 11, -14, -2, 0, 14,
    -- layer=1 filter=226 channel=102
    -31, -27, -33, -2, -19, -16, -10, 5, 0,
    -- layer=1 filter=226 channel=103
    2, 0, -13, -13, -22, -13, -17, -10, -6,
    -- layer=1 filter=226 channel=104
    12, 0, 5, 34, 12, -5, 0, -20, -31,
    -- layer=1 filter=226 channel=105
    -6, -6, -11, -6, 6, -6, 1, 2, -7,
    -- layer=1 filter=226 channel=106
    39, 8, 4, 27, 2, 8, 17, 7, 25,
    -- layer=1 filter=226 channel=107
    3, 2, 1, 8, -7, 2, 0, -11, -7,
    -- layer=1 filter=226 channel=108
    0, 14, 11, 15, 8, 17, 0, -26, 1,
    -- layer=1 filter=226 channel=109
    6, 2, 5, 0, 0, -1, 9, -1, 1,
    -- layer=1 filter=226 channel=110
    -10, -12, 3, -6, -8, 6, 1, -4, -5,
    -- layer=1 filter=226 channel=111
    -73, -72, -39, -65, -56, -37, -53, -59, -22,
    -- layer=1 filter=226 channel=112
    -17, -44, -21, -66, -30, -35, -42, -20, -15,
    -- layer=1 filter=226 channel=113
    -20, -30, -5, -22, -22, -4, -41, -34, -15,
    -- layer=1 filter=226 channel=114
    -82, -71, -63, -65, -78, -54, -60, -55, -17,
    -- layer=1 filter=226 channel=115
    17, 19, 10, 18, 20, 19, 16, 15, 22,
    -- layer=1 filter=226 channel=116
    3, 0, 8, 9, -4, -8, 0, 7, 5,
    -- layer=1 filter=226 channel=117
    -47, -63, -17, -58, -21, 3, -69, -52, -29,
    -- layer=1 filter=226 channel=118
    -32, -43, -50, -27, -35, -33, -30, -47, -11,
    -- layer=1 filter=226 channel=119
    12, 34, 3, 15, 11, 24, 2, -12, -7,
    -- layer=1 filter=226 channel=120
    4, 11, -10, -1, 6, 1, 8, 14, -21,
    -- layer=1 filter=226 channel=121
    -21, -13, 12, -7, -35, -29, -29, -40, -29,
    -- layer=1 filter=226 channel=122
    -5, 6, -3, 8, 7, -1, 9, 8, -8,
    -- layer=1 filter=226 channel=123
    -13, -22, 16, -12, -21, -18, -1, -21, 0,
    -- layer=1 filter=226 channel=124
    -14, -2, -17, -3, -7, -16, -16, -15, -8,
    -- layer=1 filter=226 channel=125
    -13, -35, -18, -31, -33, -27, -31, -41, -32,
    -- layer=1 filter=226 channel=126
    -5, -34, -36, -28, -75, -15, -9, -2, -9,
    -- layer=1 filter=226 channel=127
    -45, -69, -45, -45, -39, -58, -33, -68, -3,
    -- layer=1 filter=227 channel=0
    -2, -3, 8, -10, 5, -4, 0, 7, 1,
    -- layer=1 filter=227 channel=1
    5, -11, -12, -1, 5, 2, -5, -2, 7,
    -- layer=1 filter=227 channel=2
    -4, 0, -4, 2, -2, 0, -10, -9, 0,
    -- layer=1 filter=227 channel=3
    3, -5, 4, 8, 2, -2, 0, -4, 2,
    -- layer=1 filter=227 channel=4
    -10, 9, 1, -10, 7, -1, -3, 3, -7,
    -- layer=1 filter=227 channel=5
    -2, 6, -8, -3, -1, 0, -5, -4, 5,
    -- layer=1 filter=227 channel=6
    5, -5, 7, 5, -1, 1, -11, 0, -2,
    -- layer=1 filter=227 channel=7
    5, 0, -2, -7, -2, -1, -3, -10, -15,
    -- layer=1 filter=227 channel=8
    8, 4, 1, 0, -13, 0, 8, -3, 5,
    -- layer=1 filter=227 channel=9
    9, -7, -4, -17, -5, 1, 4, -11, 0,
    -- layer=1 filter=227 channel=10
    0, 5, 1, -11, 0, -15, -7, -12, -17,
    -- layer=1 filter=227 channel=11
    1, 4, -10, -12, 3, 1, 3, 3, -8,
    -- layer=1 filter=227 channel=12
    -6, 3, 6, -1, 6, -6, 3, -5, 15,
    -- layer=1 filter=227 channel=13
    6, 0, 1, 5, 4, -9, -8, -6, -3,
    -- layer=1 filter=227 channel=14
    -1, 1, 7, 0, -8, 2, -10, 1, -7,
    -- layer=1 filter=227 channel=15
    6, 2, 3, -5, 0, -13, -1, -8, 6,
    -- layer=1 filter=227 channel=16
    2, 3, 0, -8, 5, -10, 5, -6, -12,
    -- layer=1 filter=227 channel=17
    7, -2, 0, -9, 0, 4, 7, -4, -9,
    -- layer=1 filter=227 channel=18
    0, 7, 0, -8, -9, 0, 7, -12, 4,
    -- layer=1 filter=227 channel=19
    1, 1, -6, -11, 8, -7, 6, 6, -1,
    -- layer=1 filter=227 channel=20
    -1, -3, -10, -12, 0, -2, -12, -3, 1,
    -- layer=1 filter=227 channel=21
    -6, -6, 3, 0, 2, 7, 0, -4, 1,
    -- layer=1 filter=227 channel=22
    4, 4, -6, 7, -3, 0, -9, -5, -2,
    -- layer=1 filter=227 channel=23
    -10, -4, -9, -3, 1, 4, 5, -5, 7,
    -- layer=1 filter=227 channel=24
    -13, -4, 0, 3, -5, 0, -9, -2, -3,
    -- layer=1 filter=227 channel=25
    0, -7, 0, -9, -2, -4, 8, -9, -10,
    -- layer=1 filter=227 channel=26
    1, -3, -13, 6, 3, -5, 4, -1, 7,
    -- layer=1 filter=227 channel=27
    -9, 7, 3, -13, -4, -8, 3, 6, -9,
    -- layer=1 filter=227 channel=28
    0, -10, -7, 0, -1, -1, -5, 1, 1,
    -- layer=1 filter=227 channel=29
    4, -7, -9, 7, -5, -10, -4, 0, -12,
    -- layer=1 filter=227 channel=30
    -11, 4, -9, 0, 1, -3, -3, 0, 0,
    -- layer=1 filter=227 channel=31
    -6, 2, 7, -1, 3, -2, 7, -9, -1,
    -- layer=1 filter=227 channel=32
    1, -12, 0, -1, -10, -11, -11, 6, 4,
    -- layer=1 filter=227 channel=33
    7, -5, 2, -6, 1, -7, 10, -2, 11,
    -- layer=1 filter=227 channel=34
    5, 0, 0, 2, 0, 8, -6, 5, 1,
    -- layer=1 filter=227 channel=35
    -3, 8, 6, 5, -2, 0, -9, 6, -3,
    -- layer=1 filter=227 channel=36
    -11, -10, -9, -9, 4, 6, -7, -4, 6,
    -- layer=1 filter=227 channel=37
    -2, -11, 1, -1, -9, -2, -4, -7, -4,
    -- layer=1 filter=227 channel=38
    -5, 6, -10, -5, 1, -3, 1, 6, -3,
    -- layer=1 filter=227 channel=39
    -3, 3, 4, 1, -9, -3, 7, -4, 4,
    -- layer=1 filter=227 channel=40
    0, 0, 5, 6, 11, 4, -3, -9, 9,
    -- layer=1 filter=227 channel=41
    5, -6, 7, -2, -11, -9, -7, 0, -5,
    -- layer=1 filter=227 channel=42
    -10, 0, -8, -1, 7, 0, 1, 7, 0,
    -- layer=1 filter=227 channel=43
    4, -7, -2, -6, -10, -4, -5, -1, 3,
    -- layer=1 filter=227 channel=44
    2, 4, -4, 0, -7, 5, -4, -5, 7,
    -- layer=1 filter=227 channel=45
    -4, -1, 2, 5, -10, -1, -4, -10, -10,
    -- layer=1 filter=227 channel=46
    -13, 2, -8, -3, 0, -9, 11, 1, 5,
    -- layer=1 filter=227 channel=47
    1, 0, -2, 4, 0, 3, -8, 4, 1,
    -- layer=1 filter=227 channel=48
    2, 0, 8, 0, 0, -5, 7, 6, 3,
    -- layer=1 filter=227 channel=49
    1, -12, -6, -2, -4, -1, -9, -4, 1,
    -- layer=1 filter=227 channel=50
    -1, 1, 0, 3, 5, 7, -10, -2, -10,
    -- layer=1 filter=227 channel=51
    7, 7, -8, 6, -8, -10, 5, -7, 1,
    -- layer=1 filter=227 channel=52
    -2, -9, 0, -9, 10, 0, -2, 2, -3,
    -- layer=1 filter=227 channel=53
    2, 3, 4, -1, -3, -7, 2, -7, 1,
    -- layer=1 filter=227 channel=54
    6, 4, -3, 7, 4, -1, -1, 10, -2,
    -- layer=1 filter=227 channel=55
    -13, -9, -14, -16, -15, -12, -5, -13, -7,
    -- layer=1 filter=227 channel=56
    0, 5, -1, 8, 0, -8, -5, -1, 0,
    -- layer=1 filter=227 channel=57
    0, -2, 6, -2, -1, -6, -10, 9, -6,
    -- layer=1 filter=227 channel=58
    -8, 1, 3, -15, -11, 2, -7, 3, -4,
    -- layer=1 filter=227 channel=59
    5, -6, -9, 1, -11, -11, 1, -7, -5,
    -- layer=1 filter=227 channel=60
    -5, -4, 8, 2, 1, -12, 5, -9, 8,
    -- layer=1 filter=227 channel=61
    -1, -4, 1, 7, -3, -5, 9, 2, -7,
    -- layer=1 filter=227 channel=62
    -3, -15, -5, -9, 1, 0, 11, 7, 0,
    -- layer=1 filter=227 channel=63
    2, -10, -2, -9, 7, -7, -11, 5, 0,
    -- layer=1 filter=227 channel=64
    4, 7, 2, -6, 6, 2, -1, 7, 2,
    -- layer=1 filter=227 channel=65
    6, -3, 5, -7, 7, -11, -9, -6, -7,
    -- layer=1 filter=227 channel=66
    -2, -11, -5, 7, 8, -5, 2, -5, -3,
    -- layer=1 filter=227 channel=67
    -10, 3, -11, -1, 7, -4, -8, 4, -1,
    -- layer=1 filter=227 channel=68
    6, -6, 3, -7, -12, 3, 7, -4, 3,
    -- layer=1 filter=227 channel=69
    3, -15, 1, -16, -6, 3, 3, -12, -1,
    -- layer=1 filter=227 channel=70
    10, 12, -2, -8, 11, 4, 13, -6, 5,
    -- layer=1 filter=227 channel=71
    -7, 0, -2, 5, 7, 5, -7, 1, -7,
    -- layer=1 filter=227 channel=72
    -4, 6, -1, 3, -4, 1, 5, -9, -2,
    -- layer=1 filter=227 channel=73
    -7, -1, -5, -6, 6, -13, 1, 5, 8,
    -- layer=1 filter=227 channel=74
    3, 0, 3, -10, 7, 3, -2, -4, -3,
    -- layer=1 filter=227 channel=75
    -7, -16, 0, 3, 7, 5, 9, 3, 3,
    -- layer=1 filter=227 channel=76
    4, 1, -11, -7, -6, 6, 0, -6, -4,
    -- layer=1 filter=227 channel=77
    -10, 3, -6, 2, -1, -10, 6, 0, 7,
    -- layer=1 filter=227 channel=78
    3, 5, -10, -7, -5, 2, -7, 2, -7,
    -- layer=1 filter=227 channel=79
    1, -7, 4, -9, -1, -3, -2, -7, -8,
    -- layer=1 filter=227 channel=80
    2, 0, 6, 6, 2, 2, 3, -2, 9,
    -- layer=1 filter=227 channel=81
    -4, 4, -8, -8, 1, 8, 4, 0, -3,
    -- layer=1 filter=227 channel=82
    -11, -11, 4, 0, 0, -10, 4, -5, 8,
    -- layer=1 filter=227 channel=83
    -1, -6, -2, 1, 0, 7, -12, -1, -7,
    -- layer=1 filter=227 channel=84
    -9, 4, -10, -6, 2, 5, -5, 0, -3,
    -- layer=1 filter=227 channel=85
    0, -2, 0, 2, 1, 4, -3, 0, 5,
    -- layer=1 filter=227 channel=86
    2, 1, 8, -10, -3, -11, -2, -1, -7,
    -- layer=1 filter=227 channel=87
    2, 8, -11, 0, 6, 7, 1, -5, 0,
    -- layer=1 filter=227 channel=88
    -5, -12, -12, 9, 4, -7, 10, 4, 1,
    -- layer=1 filter=227 channel=89
    -11, 0, -4, -8, 0, -8, 0, 0, -5,
    -- layer=1 filter=227 channel=90
    3, -8, 7, -3, 1, 3, 4, -12, -3,
    -- layer=1 filter=227 channel=91
    -2, 4, 2, 1, -10, 5, 4, 3, -7,
    -- layer=1 filter=227 channel=92
    3, 3, 4, -7, -11, 7, -11, 2, -9,
    -- layer=1 filter=227 channel=93
    -8, 0, -9, -12, -4, -10, 2, -10, -11,
    -- layer=1 filter=227 channel=94
    -11, 1, 7, 4, -8, 3, -1, -4, -10,
    -- layer=1 filter=227 channel=95
    -11, 4, 3, 2, -1, -9, 3, 0, -9,
    -- layer=1 filter=227 channel=96
    5, -11, 0, 3, 7, 6, -2, -4, 6,
    -- layer=1 filter=227 channel=97
    -10, -2, 4, 8, -1, -11, -7, 1, -2,
    -- layer=1 filter=227 channel=98
    3, -12, -12, 4, -2, 0, -3, -3, 4,
    -- layer=1 filter=227 channel=99
    0, 1, 0, 3, 3, 2, -11, 7, 0,
    -- layer=1 filter=227 channel=100
    -1, 1, -11, 7, 0, -9, 2, 0, 2,
    -- layer=1 filter=227 channel=101
    -4, 1, -9, -8, -7, -6, -11, -4, -2,
    -- layer=1 filter=227 channel=102
    -10, 1, 6, -12, -8, -2, -5, -3, 2,
    -- layer=1 filter=227 channel=103
    -9, -7, -2, -5, 7, 0, 4, 0, 1,
    -- layer=1 filter=227 channel=104
    1, -11, 9, 8, -10, -4, 6, 4, 1,
    -- layer=1 filter=227 channel=105
    7, 0, 1, -8, 2, -5, -9, -5, -10,
    -- layer=1 filter=227 channel=106
    0, 1, -1, -9, -6, -2, -6, 1, -3,
    -- layer=1 filter=227 channel=107
    1, -2, -6, -10, 6, -3, 10, 5, 1,
    -- layer=1 filter=227 channel=108
    -7, -6, -20, -14, 0, -1, -17, -17, -11,
    -- layer=1 filter=227 channel=109
    6, -5, 4, -10, -6, 0, -1, 6, -3,
    -- layer=1 filter=227 channel=110
    5, -2, 0, 0, -1, -2, 2, 5, 0,
    -- layer=1 filter=227 channel=111
    0, -5, -10, 1, 2, 9, -4, -2, -5,
    -- layer=1 filter=227 channel=112
    -11, -3, 1, 6, 5, -1, 6, -8, -4,
    -- layer=1 filter=227 channel=113
    1, 0, -12, 8, -8, 6, 8, 2, -4,
    -- layer=1 filter=227 channel=114
    -9, -3, 1, -15, -14, 2, 3, 1, -1,
    -- layer=1 filter=227 channel=115
    8, 0, -6, -4, -9, 0, 7, 7, 2,
    -- layer=1 filter=227 channel=116
    10, -9, 1, 3, -5, -5, -2, -3, -2,
    -- layer=1 filter=227 channel=117
    -5, 3, -6, 6, 0, 5, -1, 4, -6,
    -- layer=1 filter=227 channel=118
    6, 4, 3, 4, -12, 4, -9, 6, 2,
    -- layer=1 filter=227 channel=119
    -1, -3, 3, -5, 3, 3, -10, -1, -5,
    -- layer=1 filter=227 channel=120
    -1, -7, -10, 5, -2, 4, -5, -5, -11,
    -- layer=1 filter=227 channel=121
    -4, -5, -6, 7, -5, -4, -7, -8, 6,
    -- layer=1 filter=227 channel=122
    -9, 5, -7, -6, -5, 4, -5, 8, -9,
    -- layer=1 filter=227 channel=123
    -11, 6, 1, -9, -5, -1, 7, -2, -9,
    -- layer=1 filter=227 channel=124
    6, -4, -8, -8, -1, -9, -7, -3, -4,
    -- layer=1 filter=227 channel=125
    11, 8, 7, -4, -11, 0, 12, 4, -2,
    -- layer=1 filter=227 channel=126
    7, -2, -3, -10, 8, -6, -12, 2, 6,
    -- layer=1 filter=227 channel=127
    -5, -8, 8, -7, 5, -3, -4, 4, -13,
    -- layer=1 filter=228 channel=0
    6, 8, 3, 4, 2, 5, -1, 2, 0,
    -- layer=1 filter=228 channel=1
    -10, 1, -12, 5, -10, -2, 0, -8, -6,
    -- layer=1 filter=228 channel=2
    6, -13, -9, -6, -9, -11, -11, 0, -1,
    -- layer=1 filter=228 channel=3
    9, 0, -5, 2, -7, 8, -10, -1, -4,
    -- layer=1 filter=228 channel=4
    2, 0, -8, 6, -7, -6, -11, -7, -8,
    -- layer=1 filter=228 channel=5
    -2, -9, 4, 6, -4, -5, -6, -11, -3,
    -- layer=1 filter=228 channel=6
    -9, 6, -5, 7, 2, 4, 7, 6, 1,
    -- layer=1 filter=228 channel=7
    -5, 7, -2, -3, 1, -5, -5, 0, -2,
    -- layer=1 filter=228 channel=8
    8, 0, -12, -2, -9, -4, -2, -2, -4,
    -- layer=1 filter=228 channel=9
    0, 8, 0, -3, 0, -10, 3, -7, -9,
    -- layer=1 filter=228 channel=10
    -7, -5, -3, 8, -9, -6, 5, -8, -9,
    -- layer=1 filter=228 channel=11
    -5, -1, -1, -2, 2, 10, -8, -3, -8,
    -- layer=1 filter=228 channel=12
    7, 4, 6, -2, 0, 3, 10, -7, -1,
    -- layer=1 filter=228 channel=13
    -3, -1, -10, -7, -2, -8, -2, -3, -11,
    -- layer=1 filter=228 channel=14
    -1, 2, -8, -7, -3, -4, -8, -4, 3,
    -- layer=1 filter=228 channel=15
    2, 0, 0, 0, -4, -8, 0, 9, 0,
    -- layer=1 filter=228 channel=16
    11, -4, 0, 6, 11, 3, 0, 9, -8,
    -- layer=1 filter=228 channel=17
    -3, -12, -1, -12, 2, 7, 8, 3, 0,
    -- layer=1 filter=228 channel=18
    0, -3, -6, -6, 1, 2, -7, 9, -9,
    -- layer=1 filter=228 channel=19
    2, 1, 3, -2, 0, 2, -10, -10, -2,
    -- layer=1 filter=228 channel=20
    -5, -1, 8, 2, -12, 2, -4, -8, -6,
    -- layer=1 filter=228 channel=21
    -4, 4, 5, 6, 8, -12, 6, -6, 4,
    -- layer=1 filter=228 channel=22
    4, 2, -8, -10, 2, 7, 3, 4, -10,
    -- layer=1 filter=228 channel=23
    4, -1, 3, 3, -9, 0, -10, 0, -6,
    -- layer=1 filter=228 channel=24
    -9, -5, 6, 10, -6, -12, 7, 6, -13,
    -- layer=1 filter=228 channel=25
    3, 1, 0, -1, 6, -1, 8, 0, -9,
    -- layer=1 filter=228 channel=26
    -1, -13, 7, -2, -9, 0, 3, 0, 1,
    -- layer=1 filter=228 channel=27
    7, 9, 0, -5, 7, -9, 0, -7, 0,
    -- layer=1 filter=228 channel=28
    0, -5, -12, 7, 0, 1, 3, 3, 8,
    -- layer=1 filter=228 channel=29
    2, 0, -3, 1, -1, 1, -5, -2, 3,
    -- layer=1 filter=228 channel=30
    3, -7, 11, -3, -5, -7, 7, 7, 3,
    -- layer=1 filter=228 channel=31
    -4, -6, 9, -2, -10, 1, 4, -3, -7,
    -- layer=1 filter=228 channel=32
    -11, 1, 4, -9, 0, -8, 1, -13, -8,
    -- layer=1 filter=228 channel=33
    3, -6, -11, -4, 10, -2, 6, -7, -5,
    -- layer=1 filter=228 channel=34
    2, -7, -11, -4, 0, -5, 7, -9, 1,
    -- layer=1 filter=228 channel=35
    -3, 9, -2, 7, -5, 0, -7, -3, 7,
    -- layer=1 filter=228 channel=36
    -11, 1, -9, -5, -10, -2, 4, -2, 0,
    -- layer=1 filter=228 channel=37
    8, 3, 7, 10, 1, -4, 5, -8, -3,
    -- layer=1 filter=228 channel=38
    -13, 3, -5, -4, -6, -6, -15, -5, 1,
    -- layer=1 filter=228 channel=39
    -7, -1, -8, 7, -1, -8, -8, -7, 2,
    -- layer=1 filter=228 channel=40
    4, 4, -8, -6, 3, -5, -3, 0, 6,
    -- layer=1 filter=228 channel=41
    0, -3, -3, -8, -13, -12, 2, -7, -10,
    -- layer=1 filter=228 channel=42
    -8, 0, 3, -1, -7, -10, -8, -10, 4,
    -- layer=1 filter=228 channel=43
    -5, -1, -10, 0, -6, 9, -7, 7, -5,
    -- layer=1 filter=228 channel=44
    -1, -2, 7, -8, -3, 7, 1, -1, -4,
    -- layer=1 filter=228 channel=45
    4, -9, 0, -1, -3, 6, 0, 0, -5,
    -- layer=1 filter=228 channel=46
    0, 4, 0, 8, -9, 6, 0, -9, 4,
    -- layer=1 filter=228 channel=47
    -11, -8, 7, -10, 1, -1, 2, -2, -9,
    -- layer=1 filter=228 channel=48
    5, -5, -12, 0, -9, -6, 4, -12, 3,
    -- layer=1 filter=228 channel=49
    1, 1, 7, 5, 5, -4, -7, -12, -4,
    -- layer=1 filter=228 channel=50
    3, 8, 2, -11, 0, 6, -11, -11, -11,
    -- layer=1 filter=228 channel=51
    6, -7, -4, -7, 1, -8, -8, -3, 6,
    -- layer=1 filter=228 channel=52
    8, -9, 0, 4, 2, 6, -2, -2, 8,
    -- layer=1 filter=228 channel=53
    -11, 4, 5, 3, 8, -11, 2, -6, 4,
    -- layer=1 filter=228 channel=54
    -5, -1, 0, -5, -2, -3, -3, 5, 10,
    -- layer=1 filter=228 channel=55
    -4, 2, 0, 1, -8, 9, 1, 3, 11,
    -- layer=1 filter=228 channel=56
    0, 0, -5, -1, 3, -4, -9, 3, 2,
    -- layer=1 filter=228 channel=57
    -9, 2, 0, 8, -5, 9, -3, 6, -4,
    -- layer=1 filter=228 channel=58
    -13, 10, -7, 3, 0, 0, -6, -6, 5,
    -- layer=1 filter=228 channel=59
    -9, -9, 7, -5, 7, 3, 1, 3, -7,
    -- layer=1 filter=228 channel=60
    4, 9, 8, -3, 1, -7, 0, 7, -10,
    -- layer=1 filter=228 channel=61
    -6, 0, -5, 9, 1, 0, -5, 4, 0,
    -- layer=1 filter=228 channel=62
    0, 0, 8, 8, -5, -5, 9, 2, -10,
    -- layer=1 filter=228 channel=63
    -8, 5, -8, -4, -8, 6, -11, -10, 0,
    -- layer=1 filter=228 channel=64
    5, 6, -11, 7, -2, -9, -9, -9, -7,
    -- layer=1 filter=228 channel=65
    -2, 6, -4, -4, 8, -4, -9, 0, -5,
    -- layer=1 filter=228 channel=66
    -9, -4, -1, 0, 0, -8, -4, -3, -9,
    -- layer=1 filter=228 channel=67
    -10, -9, -8, -10, 9, -8, -10, -3, 2,
    -- layer=1 filter=228 channel=68
    1, -3, -11, -7, -3, 0, -3, -13, -10,
    -- layer=1 filter=228 channel=69
    -9, -11, -7, -9, 2, 2, -2, -8, 0,
    -- layer=1 filter=228 channel=70
    -1, -5, -8, -9, 8, -1, 10, 3, -4,
    -- layer=1 filter=228 channel=71
    3, 7, 0, -11, -11, 1, -7, 0, 2,
    -- layer=1 filter=228 channel=72
    0, 0, -11, 7, 6, -8, -9, -11, 4,
    -- layer=1 filter=228 channel=73
    -2, 5, 0, 1, -6, -11, 2, 6, -3,
    -- layer=1 filter=228 channel=74
    -12, -2, 7, 2, -4, 4, 7, -11, 2,
    -- layer=1 filter=228 channel=75
    11, 5, -1, -8, -16, 0, -10, 7, 2,
    -- layer=1 filter=228 channel=76
    7, 6, 8, 0, -3, -11, 5, -9, 1,
    -- layer=1 filter=228 channel=77
    -2, -2, -8, -7, -11, -6, -3, -6, 3,
    -- layer=1 filter=228 channel=78
    5, 7, -2, 0, -3, -9, 0, -11, -4,
    -- layer=1 filter=228 channel=79
    0, 3, 3, -12, 3, 8, 4, -3, -5,
    -- layer=1 filter=228 channel=80
    1, 7, -7, -4, 6, 10, 9, -5, 1,
    -- layer=1 filter=228 channel=81
    -11, 3, 4, 7, -4, -7, -9, -8, -11,
    -- layer=1 filter=228 channel=82
    5, -8, -8, -4, 3, 0, -1, -9, 3,
    -- layer=1 filter=228 channel=83
    2, -4, -2, -3, 6, -3, -5, 7, -2,
    -- layer=1 filter=228 channel=84
    -8, 7, -4, -1, 2, -7, 6, 9, 5,
    -- layer=1 filter=228 channel=85
    -11, 4, 3, 0, -8, -3, -12, -2, 0,
    -- layer=1 filter=228 channel=86
    1, -2, -9, -4, 4, 7, 9, 1, 3,
    -- layer=1 filter=228 channel=87
    5, -7, 5, -3, 8, -3, -3, -2, -8,
    -- layer=1 filter=228 channel=88
    -10, 5, -11, -1, -5, -7, 0, 0, 5,
    -- layer=1 filter=228 channel=89
    -2, 0, 0, 3, 7, 2, -3, -10, -4,
    -- layer=1 filter=228 channel=90
    -12, 6, -9, -11, -1, -8, -3, -6, -9,
    -- layer=1 filter=228 channel=91
    7, -6, -3, 1, 4, 5, -4, 0, 3,
    -- layer=1 filter=228 channel=92
    -1, -3, -2, -10, -1, -5, -7, 6, 0,
    -- layer=1 filter=228 channel=93
    -9, 3, -6, -3, -8, 1, -11, -10, 2,
    -- layer=1 filter=228 channel=94
    3, -10, -9, 0, 0, 3, -10, -10, 7,
    -- layer=1 filter=228 channel=95
    0, -8, -8, 6, 2, -2, 0, 4, 0,
    -- layer=1 filter=228 channel=96
    7, -4, -1, -5, -8, 8, 3, -8, -7,
    -- layer=1 filter=228 channel=97
    5, 2, -9, -9, -7, 2, -1, -10, 0,
    -- layer=1 filter=228 channel=98
    -14, 7, 6, 10, 9, 4, 7, -4, -11,
    -- layer=1 filter=228 channel=99
    -6, -2, 5, 7, -1, -4, 1, 1, -9,
    -- layer=1 filter=228 channel=100
    -10, -3, -1, 7, -5, -1, -8, 5, 4,
    -- layer=1 filter=228 channel=101
    0, 0, -6, -2, -2, -8, -11, 5, 0,
    -- layer=1 filter=228 channel=102
    0, -5, 6, -1, -8, -9, 4, 4, -1,
    -- layer=1 filter=228 channel=103
    -6, -7, -6, 1, -4, 0, -4, 0, 7,
    -- layer=1 filter=228 channel=104
    3, 1, -10, -4, -4, 0, -11, 2, -7,
    -- layer=1 filter=228 channel=105
    6, -1, 3, -1, 2, 5, -1, -2, -5,
    -- layer=1 filter=228 channel=106
    -9, -3, -2, -7, -3, -10, -7, 4, -11,
    -- layer=1 filter=228 channel=107
    -6, 5, 8, -10, 4, -2, -3, 10, -7,
    -- layer=1 filter=228 channel=108
    -5, -7, 5, -9, 8, 0, 5, 2, 2,
    -- layer=1 filter=228 channel=109
    5, -11, 4, 9, 6, 11, 2, 9, 6,
    -- layer=1 filter=228 channel=110
    -6, 5, 0, -7, -4, 6, 1, 1, -11,
    -- layer=1 filter=228 channel=111
    -9, 2, 9, -7, -7, -6, 3, -9, 5,
    -- layer=1 filter=228 channel=112
    5, -3, -11, 7, 0, -7, 6, 0, 2,
    -- layer=1 filter=228 channel=113
    -3, 5, -4, -4, -10, 6, 3, -1, 5,
    -- layer=1 filter=228 channel=114
    -1, -9, -2, -11, 7, -6, 4, -4, -8,
    -- layer=1 filter=228 channel=115
    1, -6, 7, -1, 7, -10, -7, 7, 4,
    -- layer=1 filter=228 channel=116
    -2, -8, 7, -7, 0, 0, 5, 5, 7,
    -- layer=1 filter=228 channel=117
    -10, -6, 2, -9, 2, -3, -4, 8, 7,
    -- layer=1 filter=228 channel=118
    5, -8, -9, 6, -2, 3, 1, 5, 1,
    -- layer=1 filter=228 channel=119
    4, 7, 9, 1, 9, 3, -1, 7, -2,
    -- layer=1 filter=228 channel=120
    -15, -2, 6, -8, 0, 11, -3, 3, 3,
    -- layer=1 filter=228 channel=121
    0, -4, 8, 5, -3, 5, 2, 1, -10,
    -- layer=1 filter=228 channel=122
    -9, 2, -6, 3, -2, 3, 5, -8, 2,
    -- layer=1 filter=228 channel=123
    -5, 6, 7, -2, 2, 0, -13, -5, 3,
    -- layer=1 filter=228 channel=124
    9, 7, 1, 0, -6, -8, 3, -5, -7,
    -- layer=1 filter=228 channel=125
    6, 5, 9, 0, -9, -3, 0, 3, -9,
    -- layer=1 filter=228 channel=126
    3, 0, 7, -7, -1, 0, -7, 6, 4,
    -- layer=1 filter=228 channel=127
    0, -9, -8, -10, -14, -4, 0, -4, -7,
    -- layer=1 filter=229 channel=0
    5, 4, 5, 5, 7, 2, 4, -11, -8,
    -- layer=1 filter=229 channel=1
    -7, 7, -2, -13, 2, -1, -7, -11, 4,
    -- layer=1 filter=229 channel=2
    6, -5, 1, 1, 1, 3, -10, 0, -8,
    -- layer=1 filter=229 channel=3
    6, -4, -3, 5, -3, 8, 2, -9, 9,
    -- layer=1 filter=229 channel=4
    -2, 8, -2, -12, 6, -3, -10, -8, 4,
    -- layer=1 filter=229 channel=5
    -7, 2, 5, -2, -3, 0, -10, -9, 0,
    -- layer=1 filter=229 channel=6
    0, -1, -8, -1, -7, 6, -8, 5, -3,
    -- layer=1 filter=229 channel=7
    2, -18, 3, 2, 0, 3, -1, -2, -7,
    -- layer=1 filter=229 channel=8
    -10, 2, -6, -2, 7, 5, -8, 3, 3,
    -- layer=1 filter=229 channel=9
    4, -14, -12, -10, 0, -11, -8, -4, -6,
    -- layer=1 filter=229 channel=10
    -13, 0, -2, -4, -4, 0, 0, 0, -8,
    -- layer=1 filter=229 channel=11
    -4, -10, -4, -3, -8, 2, 9, 0, -8,
    -- layer=1 filter=229 channel=12
    2, -5, 9, -13, -13, 0, -2, 1, -7,
    -- layer=1 filter=229 channel=13
    -9, -3, 0, -5, 5, -6, -14, -14, -1,
    -- layer=1 filter=229 channel=14
    -9, 0, 8, -2, 6, -9, -5, -5, -12,
    -- layer=1 filter=229 channel=15
    -6, 8, -1, -1, 0, 1, 1, 5, 5,
    -- layer=1 filter=229 channel=16
    3, -4, 1, -14, 2, 2, 4, -6, 0,
    -- layer=1 filter=229 channel=17
    -2, -4, -12, -3, 3, 3, -3, -8, 4,
    -- layer=1 filter=229 channel=18
    -8, -8, -5, -14, -9, -16, -12, -12, 4,
    -- layer=1 filter=229 channel=19
    7, -11, 7, -3, -8, 5, -6, -4, 6,
    -- layer=1 filter=229 channel=20
    -5, 5, -4, -8, 6, 4, -9, -3, -13,
    -- layer=1 filter=229 channel=21
    -10, 3, -8, 2, -12, -10, -2, 1, -12,
    -- layer=1 filter=229 channel=22
    4, -11, -10, -3, -9, -11, -11, 5, -7,
    -- layer=1 filter=229 channel=23
    7, -5, -8, 3, -10, 6, -9, 7, 7,
    -- layer=1 filter=229 channel=24
    3, -5, -14, -16, 6, 2, -1, 5, -14,
    -- layer=1 filter=229 channel=25
    -3, 0, 0, 0, -9, -2, -2, 5, -2,
    -- layer=1 filter=229 channel=26
    -14, 3, -2, -8, -10, -11, -16, -6, 2,
    -- layer=1 filter=229 channel=27
    -4, 3, -6, 7, 0, 6, -11, 8, 1,
    -- layer=1 filter=229 channel=28
    4, -10, 9, 4, -8, -3, 1, -6, -9,
    -- layer=1 filter=229 channel=29
    8, -9, 7, -6, -4, 1, -5, -2, 1,
    -- layer=1 filter=229 channel=30
    -13, 0, -14, -9, -5, -14, 4, -2, -5,
    -- layer=1 filter=229 channel=31
    0, -9, -17, 3, -2, 2, -9, -3, 1,
    -- layer=1 filter=229 channel=32
    -1, -6, -3, -12, -7, -8, 4, -1, -2,
    -- layer=1 filter=229 channel=33
    -11, -10, -11, 4, 9, 1, 4, 6, -7,
    -- layer=1 filter=229 channel=34
    -3, 8, 10, -12, 0, -4, -4, -5, 2,
    -- layer=1 filter=229 channel=35
    2, -10, 4, 5, 7, 3, -7, -9, -6,
    -- layer=1 filter=229 channel=36
    -10, -9, 7, -4, 6, 0, 6, -6, -9,
    -- layer=1 filter=229 channel=37
    6, -11, -15, -12, 0, -11, -12, -6, -1,
    -- layer=1 filter=229 channel=38
    -1, -7, 0, -3, 3, 1, 1, -1, -4,
    -- layer=1 filter=229 channel=39
    3, 6, -10, -8, -2, 9, 0, 4, 2,
    -- layer=1 filter=229 channel=40
    6, -11, -2, -1, -1, -3, 0, -9, -12,
    -- layer=1 filter=229 channel=41
    -8, -6, 2, 8, 9, -10, -9, 6, 9,
    -- layer=1 filter=229 channel=42
    0, -2, -2, -7, -8, -3, -8, -18, -15,
    -- layer=1 filter=229 channel=43
    -9, 6, 10, 3, -3, 8, -7, 2, -2,
    -- layer=1 filter=229 channel=44
    0, -10, 1, -14, -8, -8, 1, -11, -3,
    -- layer=1 filter=229 channel=45
    -10, -4, 2, 1, -10, 0, 5, 1, 3,
    -- layer=1 filter=229 channel=46
    -13, -9, -13, -18, -14, -1, -6, -13, -1,
    -- layer=1 filter=229 channel=47
    -12, 5, -13, -8, -7, -3, -13, -4, 8,
    -- layer=1 filter=229 channel=48
    8, 0, 0, 7, -7, -7, 1, -9, 1,
    -- layer=1 filter=229 channel=49
    -3, 6, -8, -3, -1, -5, 6, -2, -11,
    -- layer=1 filter=229 channel=50
    9, -3, -10, 7, 1, 1, -12, -1, 7,
    -- layer=1 filter=229 channel=51
    -7, -4, -5, 3, -3, -4, 6, -12, -2,
    -- layer=1 filter=229 channel=52
    -3, -2, 4, -3, 2, 8, -1, -12, 8,
    -- layer=1 filter=229 channel=53
    -2, 1, -7, 7, 4, -1, 0, -9, -8,
    -- layer=1 filter=229 channel=54
    8, -17, 6, -5, 0, -5, -1, 3, -6,
    -- layer=1 filter=229 channel=55
    3, 2, -2, 1, -5, -2, -1, -12, -6,
    -- layer=1 filter=229 channel=56
    -5, 0, -5, 4, 6, 0, -7, -6, -6,
    -- layer=1 filter=229 channel=57
    -10, -19, -6, 5, -9, 5, 0, 0, -12,
    -- layer=1 filter=229 channel=58
    4, -10, 6, -6, 2, -11, -10, 10, -1,
    -- layer=1 filter=229 channel=59
    -9, -7, -4, 8, 2, -5, 7, 3, 4,
    -- layer=1 filter=229 channel=60
    3, -10, -10, 2, -3, 1, 0, 4, 6,
    -- layer=1 filter=229 channel=61
    -9, 3, -10, 7, 0, -11, 6, -6, 7,
    -- layer=1 filter=229 channel=62
    10, -3, -9, -15, -9, 3, 3, 10, 3,
    -- layer=1 filter=229 channel=63
    -6, 1, -2, 5, 0, 5, -12, 6, -6,
    -- layer=1 filter=229 channel=64
    4, -1, 0, -2, 0, 4, -11, -8, 6,
    -- layer=1 filter=229 channel=65
    0, -4, 5, -12, 1, 2, -5, -2, 7,
    -- layer=1 filter=229 channel=66
    6, -9, 2, 1, -7, -5, -3, -11, -5,
    -- layer=1 filter=229 channel=67
    1, 4, 1, -7, -6, -4, -3, 4, -2,
    -- layer=1 filter=229 channel=68
    -1, -12, -10, -13, -4, -1, 1, 4, -7,
    -- layer=1 filter=229 channel=69
    -6, 0, 1, -3, -3, 1, -9, -5, -10,
    -- layer=1 filter=229 channel=70
    -2, -10, -13, 3, -5, 0, 2, -7, -15,
    -- layer=1 filter=229 channel=71
    1, -8, -1, -9, -3, -11, 2, 0, 0,
    -- layer=1 filter=229 channel=72
    1, -8, 7, -9, 6, -5, -6, -7, 8,
    -- layer=1 filter=229 channel=73
    0, -7, 7, -7, 2, -8, 4, 0, -9,
    -- layer=1 filter=229 channel=74
    4, -2, 5, -11, 1, 6, 6, -1, 6,
    -- layer=1 filter=229 channel=75
    -5, -11, -3, -1, -2, -8, 3, -2, 5,
    -- layer=1 filter=229 channel=76
    -4, 2, -11, -11, -5, 1, -6, -6, 6,
    -- layer=1 filter=229 channel=77
    4, -11, 7, -5, -1, 0, 1, 6, 5,
    -- layer=1 filter=229 channel=78
    4, -10, 0, -6, 0, 6, -8, 0, -10,
    -- layer=1 filter=229 channel=79
    7, -5, -13, -13, -9, -9, -8, 8, -6,
    -- layer=1 filter=229 channel=80
    0, 3, -2, 7, -1, 0, -7, -13, -9,
    -- layer=1 filter=229 channel=81
    -7, 0, 3, -4, -8, 2, 0, 0, 1,
    -- layer=1 filter=229 channel=82
    8, 7, 0, 0, -1, -2, -12, -7, 5,
    -- layer=1 filter=229 channel=83
    -2, 0, 0, 5, 7, 3, 7, -3, -6,
    -- layer=1 filter=229 channel=84
    0, -1, 0, -18, -10, -13, -5, -11, 3,
    -- layer=1 filter=229 channel=85
    10, -6, 0, -3, 4, -3, -10, 0, 4,
    -- layer=1 filter=229 channel=86
    4, 0, -10, 0, -11, 7, -10, 7, 4,
    -- layer=1 filter=229 channel=87
    -7, -9, 9, -10, 5, -3, 7, 2, 2,
    -- layer=1 filter=229 channel=88
    1, -9, 0, -8, -10, -12, 4, -3, -8,
    -- layer=1 filter=229 channel=89
    0, -12, -9, -4, -12, -2, -12, -4, -2,
    -- layer=1 filter=229 channel=90
    -4, 0, 0, -11, -4, 0, -11, -3, 0,
    -- layer=1 filter=229 channel=91
    7, -9, 0, -1, -5, -8, -13, 0, -10,
    -- layer=1 filter=229 channel=92
    4, 0, 3, -10, 5, -3, 3, 3, -8,
    -- layer=1 filter=229 channel=93
    -5, -7, -5, -12, -8, 4, -4, -10, 5,
    -- layer=1 filter=229 channel=94
    -4, 5, -9, -4, -9, 2, -8, -5, 5,
    -- layer=1 filter=229 channel=95
    0, -8, -12, -6, -6, 2, 0, 2, -6,
    -- layer=1 filter=229 channel=96
    6, 4, 4, 6, 4, -6, 7, 7, 9,
    -- layer=1 filter=229 channel=97
    4, -5, 4, -8, 0, -11, -5, 0, 1,
    -- layer=1 filter=229 channel=98
    -5, -1, -5, -15, -2, -1, -4, 5, 3,
    -- layer=1 filter=229 channel=99
    -6, 0, -8, -11, -1, -4, 5, 2, -10,
    -- layer=1 filter=229 channel=100
    7, 0, -6, 9, 1, -2, 1, 0, 1,
    -- layer=1 filter=229 channel=101
    1, 5, 6, -11, -11, 1, 6, 0, 0,
    -- layer=1 filter=229 channel=102
    3, -3, -9, -11, 0, -10, 0, -11, -5,
    -- layer=1 filter=229 channel=103
    -1, 2, 8, 9, -5, 1, -9, -2, 1,
    -- layer=1 filter=229 channel=104
    -2, -4, 6, -8, -8, 7, 2, -10, -6,
    -- layer=1 filter=229 channel=105
    -11, -9, 8, -9, -5, -2, -3, 5, -8,
    -- layer=1 filter=229 channel=106
    -2, -13, 2, -2, -1, 0, 7, -2, 4,
    -- layer=1 filter=229 channel=107
    6, -5, -7, 3, -2, 1, 0, -9, -1,
    -- layer=1 filter=229 channel=108
    -18, 3, 0, -6, 3, -10, -10, -11, 10,
    -- layer=1 filter=229 channel=109
    1, -10, 0, -6, -8, -4, 1, -5, -6,
    -- layer=1 filter=229 channel=110
    -2, -1, -8, -4, 0, -2, 5, -8, 4,
    -- layer=1 filter=229 channel=111
    -2, -9, -13, -4, 2, 0, -7, 4, 4,
    -- layer=1 filter=229 channel=112
    3, 5, 2, -11, 8, 2, -7, 4, 2,
    -- layer=1 filter=229 channel=113
    2, -9, -5, -11, 4, 2, -8, -7, -1,
    -- layer=1 filter=229 channel=114
    -4, 10, -6, -11, -10, -5, -6, 0, 8,
    -- layer=1 filter=229 channel=115
    -10, -7, 3, 2, -1, -11, 2, 7, -7,
    -- layer=1 filter=229 channel=116
    7, 8, 10, 0, -1, -5, 3, 8, -8,
    -- layer=1 filter=229 channel=117
    0, 5, -9, 3, 1, 4, -9, -2, 4,
    -- layer=1 filter=229 channel=118
    -5, -11, -13, 2, 2, 3, 8, 6, 0,
    -- layer=1 filter=229 channel=119
    0, 7, 2, 1, -2, -9, -5, 0, 0,
    -- layer=1 filter=229 channel=120
    -1, -2, -5, -15, 5, -6, -11, -1, -8,
    -- layer=1 filter=229 channel=121
    1, -12, -6, -18, -8, 0, -3, -8, 1,
    -- layer=1 filter=229 channel=122
    7, 6, 9, -4, -9, -8, 7, -9, -4,
    -- layer=1 filter=229 channel=123
    -8, -6, 7, -13, 2, 6, -1, -10, -10,
    -- layer=1 filter=229 channel=124
    6, -11, 2, 3, -10, -4, 0, -12, -5,
    -- layer=1 filter=229 channel=125
    3, -2, -17, 4, 11, -12, 0, -3, -9,
    -- layer=1 filter=229 channel=126
    1, -10, 0, 6, -6, -6, -2, -12, -9,
    -- layer=1 filter=229 channel=127
    -5, -10, 1, -15, -15, -8, -8, 7, 9,
    -- layer=1 filter=230 channel=0
    -5, 3, -29, -5, -8, -28, -23, 6, -13,
    -- layer=1 filter=230 channel=1
    -29, -21, 6, -46, -39, 22, -1, -85, -11,
    -- layer=1 filter=230 channel=2
    62, 61, 65, 61, 53, 49, 77, 75, 49,
    -- layer=1 filter=230 channel=3
    15, 1, -8, -6, 5, -4, 1, -3, 10,
    -- layer=1 filter=230 channel=4
    -17, -5, -18, -8, -8, 0, -4, -2, -9,
    -- layer=1 filter=230 channel=5
    -25, -20, -11, -47, -48, 6, -2, -45, 17,
    -- layer=1 filter=230 channel=6
    -4, -31, 2, -60, -21, -35, -73, -17, -1,
    -- layer=1 filter=230 channel=7
    61, -21, -41, 8, -51, -35, -49, -20, 15,
    -- layer=1 filter=230 channel=8
    -34, -34, -8, -83, -38, 38, -40, -66, 2,
    -- layer=1 filter=230 channel=9
    59, 83, 85, 36, 72, 30, 74, 53, 62,
    -- layer=1 filter=230 channel=10
    68, -43, -37, -15, -28, -31, -39, 6, 20,
    -- layer=1 filter=230 channel=11
    -79, -39, -42, -35, -19, -20, -11, -16, -25,
    -- layer=1 filter=230 channel=12
    57, 56, 70, 86, 29, 61, 64, 76, 73,
    -- layer=1 filter=230 channel=13
    -65, 14, -20, -43, -32, -25, -46, -40, -23,
    -- layer=1 filter=230 channel=14
    72, 21, 22, 50, 11, -24, 35, 36, 38,
    -- layer=1 filter=230 channel=15
    16, 70, 31, 58, 38, 56, 68, 26, 72,
    -- layer=1 filter=230 channel=16
    -34, -30, -5, -57, -34, 8, -22, -48, 37,
    -- layer=1 filter=230 channel=17
    -41, 32, -14, -29, -10, 3, -30, 6, -28,
    -- layer=1 filter=230 channel=18
    -30, -34, 1, -19, -17, -45, -49, -42, -32,
    -- layer=1 filter=230 channel=19
    49, 28, 20, -32, 36, -12, -26, -25, 81,
    -- layer=1 filter=230 channel=20
    -59, -22, -37, -76, -29, -23, -59, -68, -14,
    -- layer=1 filter=230 channel=21
    -9, -9, 5, -13, -6, 8, -9, -14, -6,
    -- layer=1 filter=230 channel=22
    -81, -37, -51, -50, -36, 6, -43, -73, -48,
    -- layer=1 filter=230 channel=23
    61, 21, -1, 23, -33, 7, -1, 0, 52,
    -- layer=1 filter=230 channel=24
    0, 10, 19, -6, 0, 2, -3, -5, 24,
    -- layer=1 filter=230 channel=25
    53, -27, -20, -18, -20, -7, -46, -13, 15,
    -- layer=1 filter=230 channel=26
    -67, 33, 19, -32, -11, -7, -29, -65, -14,
    -- layer=1 filter=230 channel=27
    43, 46, 45, 59, 65, 54, 70, 69, 44,
    -- layer=1 filter=230 channel=28
    45, -51, -39, -20, -39, -36, -69, -5, 0,
    -- layer=1 filter=230 channel=29
    27, 6, 25, 26, 9, 12, 13, 11, 21,
    -- layer=1 filter=230 channel=30
    1, -16, 15, -79, -9, -53, -33, -52, 11,
    -- layer=1 filter=230 channel=31
    30, 9, 43, 43, 39, 15, 37, 48, 27,
    -- layer=1 filter=230 channel=32
    -55, 39, 7, -28, -18, -25, -22, -37, -17,
    -- layer=1 filter=230 channel=33
    -18, -15, -14, 3, 19, 1, -3, 26, 36,
    -- layer=1 filter=230 channel=34
    9, -8, -15, 33, -11, -13, -25, -13, 9,
    -- layer=1 filter=230 channel=35
    13, 8, 17, 0, -1, 10, 17, 12, 4,
    -- layer=1 filter=230 channel=36
    -56, -27, -33, -37, -10, -26, -13, -17, -18,
    -- layer=1 filter=230 channel=37
    5, -5, 15, -33, -13, 13, -21, -22, 43,
    -- layer=1 filter=230 channel=38
    -9, -14, -13, -37, -12, -27, -20, -18, -3,
    -- layer=1 filter=230 channel=39
    -44, -9, 2, -36, -35, -21, -12, -43, 6,
    -- layer=1 filter=230 channel=40
    -2, -38, -10, -15, -10, -51, -29, -11, -6,
    -- layer=1 filter=230 channel=41
    0, 63, 52, -12, 25, 28, 13, 16, 0,
    -- layer=1 filter=230 channel=42
    51, 41, 56, 52, 57, 51, 69, 65, 41,
    -- layer=1 filter=230 channel=43
    -36, -28, -36, -65, -44, 6, -49, -40, 24,
    -- layer=1 filter=230 channel=44
    -82, 47, -13, -52, -35, -32, -38, -71, -3,
    -- layer=1 filter=230 channel=45
    -38, 26, -4, -24, -1, -12, -17, -35, 9,
    -- layer=1 filter=230 channel=46
    71, 49, 61, 47, 48, 29, 24, 29, 76,
    -- layer=1 filter=230 channel=47
    54, 30, 50, 43, -2, 49, 39, 43, 28,
    -- layer=1 filter=230 channel=48
    27, -13, -17, -4, -1, -14, -14, 2, 11,
    -- layer=1 filter=230 channel=49
    28, 35, 39, 34, 13, 35, 38, 36, 20,
    -- layer=1 filter=230 channel=50
    10, -6, -13, 16, -3, 6, 6, -20, 3,
    -- layer=1 filter=230 channel=51
    34, -26, -23, -13, -26, -25, -13, -15, -4,
    -- layer=1 filter=230 channel=52
    -6, -4, -12, -20, 38, 2, -9, -2, -19,
    -- layer=1 filter=230 channel=53
    1, 10, -8, 6, 0, -6, -8, -7, -9,
    -- layer=1 filter=230 channel=54
    51, 7, -4, 0, 14, 5, -9, 15, 46,
    -- layer=1 filter=230 channel=55
    2, 0, 19, -8, 8, 5, 12, 5, 7,
    -- layer=1 filter=230 channel=56
    0, -10, -5, -2, -4, 1, -7, -6, 7,
    -- layer=1 filter=230 channel=57
    45, -31, -17, -11, 0, -19, -28, 9, 20,
    -- layer=1 filter=230 channel=58
    89, -19, -4, 20, -19, 6, 6, -2, 45,
    -- layer=1 filter=230 channel=59
    6, -5, 1, -11, -12, -7, -12, 0, 4,
    -- layer=1 filter=230 channel=60
    -7, -29, 9, -2, 20, 19, -12, 40, -5,
    -- layer=1 filter=230 channel=61
    4, -9, 8, 9, -3, 0, 4, -5, -4,
    -- layer=1 filter=230 channel=62
    -53, -51, -27, -92, -41, 21, -38, -30, 34,
    -- layer=1 filter=230 channel=63
    -54, -41, -19, -32, -18, -32, -32, -20, -12,
    -- layer=1 filter=230 channel=64
    14, -6, 0, -9, -19, -1, -6, 3, -42,
    -- layer=1 filter=230 channel=65
    -1, -7, -12, -13, -6, 2, 5, -5, 2,
    -- layer=1 filter=230 channel=66
    0, -16, -37, 4, -6, -8, -13, 0, -7,
    -- layer=1 filter=230 channel=67
    16, 4, 13, -9, 0, 13, -7, 0, 7,
    -- layer=1 filter=230 channel=68
    -82, 31, 5, -60, -19, -23, -62, -52, -8,
    -- layer=1 filter=230 channel=69
    -9, 15, 7, -11, -9, 3, -1, -24, 27,
    -- layer=1 filter=230 channel=70
    35, 24, 37, -5, 3, -19, -56, -4, 54,
    -- layer=1 filter=230 channel=71
    18, 4, 0, 4, -13, -9, -5, -9, 10,
    -- layer=1 filter=230 channel=72
    13, 11, 29, -28, 10, -19, -29, -33, 51,
    -- layer=1 filter=230 channel=73
    -2, 0, -4, -2, -4, -3, 11, 0, -5,
    -- layer=1 filter=230 channel=74
    -17, 1, 30, -80, 10, -59, -67, 36, -18,
    -- layer=1 filter=230 channel=75
    71, 25, 38, 52, 17, 22, 18, 49, 48,
    -- layer=1 filter=230 channel=76
    -60, 24, -3, -26, -20, -3, -43, -13, -25,
    -- layer=1 filter=230 channel=77
    -4, 7, -9, -33, 2, 1, -25, -15, 0,
    -- layer=1 filter=230 channel=78
    21, 0, -17, -7, -7, -37, -14, -4, -4,
    -- layer=1 filter=230 channel=79
    -31, -42, -13, -66, -30, 29, -44, -32, 47,
    -- layer=1 filter=230 channel=80
    51, 3, 37, 32, 9, 46, 39, 10, 37,
    -- layer=1 filter=230 channel=81
    -12, -16, 3, -7, 1, 8, -25, -20, 13,
    -- layer=1 filter=230 channel=82
    -9, -3, -15, -6, -17, -5, -28, -19, -9,
    -- layer=1 filter=230 channel=83
    -26, 30, -5, -49, -15, -14, -20, -71, 19,
    -- layer=1 filter=230 channel=84
    -64, -32, 0, -67, -27, -50, -78, -42, -68,
    -- layer=1 filter=230 channel=85
    56, 28, 0, 27, -8, 42, 11, 34, 57,
    -- layer=1 filter=230 channel=86
    -18, -22, -23, -29, -36, -44, -13, -23, -27,
    -- layer=1 filter=230 channel=87
    84, 54, 64, 26, 67, 49, 52, 48, 103,
    -- layer=1 filter=230 channel=88
    25, 27, 19, 32, 22, 25, 37, 26, 37,
    -- layer=1 filter=230 channel=89
    -23, -9, -16, -17, -30, -24, -22, -24, -11,
    -- layer=1 filter=230 channel=90
    -83, 49, -11, -91, -32, -30, -41, -85, -4,
    -- layer=1 filter=230 channel=91
    -4, -51, -32, -34, -47, -53, -56, -54, -30,
    -- layer=1 filter=230 channel=92
    17, 77, 47, 27, 43, 69, 51, 20, 66,
    -- layer=1 filter=230 channel=93
    -30, -25, -36, -33, -45, -29, -44, -31, -7,
    -- layer=1 filter=230 channel=94
    1, -30, -22, 5, -3, -43, 5, 4, -30,
    -- layer=1 filter=230 channel=95
    -18, -39, 12, -51, -16, -65, -62, -36, -6,
    -- layer=1 filter=230 channel=96
    53, 48, 57, 77, 48, 61, 71, 61, 50,
    -- layer=1 filter=230 channel=97
    -26, -13, -28, -11, -14, -15, -26, -16, -21,
    -- layer=1 filter=230 channel=98
    -49, -35, -27, -78, -23, 25, -64, -34, 0,
    -- layer=1 filter=230 channel=99
    -2, -44, -38, -90, 0, -53, -39, 27, -31,
    -- layer=1 filter=230 channel=100
    -49, -31, 11, -13, -8, -14, -8, -4, -18,
    -- layer=1 filter=230 channel=101
    -46, -48, -44, -45, -54, -40, -64, -38, -47,
    -- layer=1 filter=230 channel=102
    -6, -15, 0, -4, 12, -23, -7, 0, -24,
    -- layer=1 filter=230 channel=103
    -43, -9, -14, -7, 4, 9, 14, -19, -25,
    -- layer=1 filter=230 channel=104
    61, 45, 25, 13, -12, 29, 14, -29, 18,
    -- layer=1 filter=230 channel=105
    -10, -23, -50, -19, -8, -39, -12, -8, -20,
    -- layer=1 filter=230 channel=106
    -68, 7, -14, -49, -30, -36, -45, -44, -49,
    -- layer=1 filter=230 channel=107
    -19, -16, -11, -3, -6, 0, -17, -1, 0,
    -- layer=1 filter=230 channel=108
    -41, 46, 10, -27, -35, -11, -12, -42, 7,
    -- layer=1 filter=230 channel=109
    -7, -2, -6, -6, -10, 8, 5, -3, -7,
    -- layer=1 filter=230 channel=110
    3, 11, 24, -11, -8, -18, -3, -14, -2,
    -- layer=1 filter=230 channel=111
    -31, -25, -4, -61, -11, -65, -41, -30, -4,
    -- layer=1 filter=230 channel=112
    -35, -26, 2, -13, -22, -12, -80, -52, -33,
    -- layer=1 filter=230 channel=113
    42, 31, 42, 55, 59, 51, 42, 57, 49,
    -- layer=1 filter=230 channel=114
    1, 6, 31, -28, -15, 12, 7, -29, 45,
    -- layer=1 filter=230 channel=115
    18, -47, -42, -11, -50, -49, -30, -12, 7,
    -- layer=1 filter=230 channel=116
    2, -3, 3, 9, 6, 6, 7, 1, 0,
    -- layer=1 filter=230 channel=117
    11, 13, -9, 0, 26, -31, -16, -52, 11,
    -- layer=1 filter=230 channel=118
    -28, -18, 2, -68, -4, -54, -55, -37, -14,
    -- layer=1 filter=230 channel=119
    -58, 49, 8, -62, -33, -30, -37, -47, -22,
    -- layer=1 filter=230 channel=120
    28, -8, -8, -16, -23, -6, -17, -10, 17,
    -- layer=1 filter=230 channel=121
    45, 0, 44, 30, 33, 18, 27, 38, 17,
    -- layer=1 filter=230 channel=122
    6, -8, -3, 9, -6, -3, -2, -1, -10,
    -- layer=1 filter=230 channel=123
    23, -5, 20, 20, 3, -1, 8, 13, 15,
    -- layer=1 filter=230 channel=124
    23, 34, 35, 23, 38, 24, 30, 15, 40,
    -- layer=1 filter=230 channel=125
    52, -2, 44, -19, 1, 4, 4, 0, 35,
    -- layer=1 filter=230 channel=126
    -46, 42, 0, -43, -10, 30, -87, -63, -33,
    -- layer=1 filter=230 channel=127
    -30, -36, -2, -54, -14, -49, -63, -27, -5,
    -- layer=1 filter=231 channel=0
    -1, 27, 26, -47, -1, 37, -58, -29, 15,
    -- layer=1 filter=231 channel=1
    -15, -24, 19, -12, -53, -26, 13, -13, -73,
    -- layer=1 filter=231 channel=2
    -22, -19, -10, -14, -15, -49, -6, 9, 31,
    -- layer=1 filter=231 channel=3
    -3, 6, 3, -9, -1, -1, 4, -2, 7,
    -- layer=1 filter=231 channel=4
    8, 19, 8, -4, -15, -3, 4, 1, 0,
    -- layer=1 filter=231 channel=5
    -50, -28, -1, 15, -61, -81, 49, -35, -104,
    -- layer=1 filter=231 channel=6
    -17, -38, -69, 19, -6, -32, 0, -11, 19,
    -- layer=1 filter=231 channel=7
    81, 81, 27, 56, 93, 100, -37, 64, 100,
    -- layer=1 filter=231 channel=8
    -73, -35, -6, -31, -76, -43, 6, -80, -118,
    -- layer=1 filter=231 channel=9
    -15, -45, -11, -7, -59, 37, 31, -47, -37,
    -- layer=1 filter=231 channel=10
    69, 69, 38, 28, 70, 100, -42, 37, 100,
    -- layer=1 filter=231 channel=11
    -7, 12, 20, -1, 0, 14, -5, -15, -6,
    -- layer=1 filter=231 channel=12
    16, 10, -43, -2, 23, -20, 6, -3, 26,
    -- layer=1 filter=231 channel=13
    -12, -11, 11, -4, -45, -9, 14, -41, -26,
    -- layer=1 filter=231 channel=14
    59, 72, 19, 73, 67, 97, -28, 66, 108,
    -- layer=1 filter=231 channel=15
    31, 14, 67, 52, 71, 6, 103, 72, 8,
    -- layer=1 filter=231 channel=16
    -97, -52, -25, -60, -93, -86, -10, -109, -130,
    -- layer=1 filter=231 channel=17
    -4, 16, 44, -69, -16, 33, -33, -70, -8,
    -- layer=1 filter=231 channel=18
    67, 45, -6, 31, 41, 51, -14, 4, 74,
    -- layer=1 filter=231 channel=19
    -44, -68, -9, -32, -31, -78, -28, -53, -37,
    -- layer=1 filter=231 channel=20
    -22, -1, 24, 3, 2, -7, 3, -12, -22,
    -- layer=1 filter=231 channel=21
    19, -15, 0, 23, 2, 7, 36, 27, 13,
    -- layer=1 filter=231 channel=22
    -5, -13, 35, 0, -17, -11, 29, 5, -51,
    -- layer=1 filter=231 channel=23
    -9, -1, -55, -43, -15, -10, -31, -18, 24,
    -- layer=1 filter=231 channel=24
    -13, 4, 19, 10, -21, 0, 49, 3, -49,
    -- layer=1 filter=231 channel=25
    -32, -1, 6, -41, -5, 27, -60, -35, 17,
    -- layer=1 filter=231 channel=26
    -37, -28, 34, -23, -52, -4, 48, -23, -94,
    -- layer=1 filter=231 channel=27
    -29, -17, -4, -15, -21, -41, 16, 1, -27,
    -- layer=1 filter=231 channel=28
    27, 30, 23, -2, 37, 92, -42, 18, 60,
    -- layer=1 filter=231 channel=29
    -11, 10, -13, 7, 12, -8, 3, 4, -3,
    -- layer=1 filter=231 channel=30
    64, 27, -11, 16, 77, 48, -2, 23, 78,
    -- layer=1 filter=231 channel=31
    37, 18, -57, 43, 62, 22, 9, 40, 92,
    -- layer=1 filter=231 channel=32
    -32, -73, -5, -19, -90, -49, 41, -21, -94,
    -- layer=1 filter=231 channel=33
    -31, -6, -14, 31, 32, 1, 52, 51, -11,
    -- layer=1 filter=231 channel=34
    15, 23, 14, 13, 16, 32, 39, 23, 30,
    -- layer=1 filter=231 channel=35
    -2, 0, -11, -6, -3, -8, 1, -12, 1,
    -- layer=1 filter=231 channel=36
    -7, 7, 28, -43, -8, 12, -21, -30, -18,
    -- layer=1 filter=231 channel=37
    -96, -63, -15, -40, -82, -102, 3, -74, -91,
    -- layer=1 filter=231 channel=38
    3, -1, 12, 19, 6, 7, -4, 15, 1,
    -- layer=1 filter=231 channel=39
    -23, -2, 14, -29, -31, 8, -44, -46, -27,
    -- layer=1 filter=231 channel=40
    71, 28, -52, 35, 60, 56, -32, 20, 97,
    -- layer=1 filter=231 channel=41
    -34, -106, -48, -41, -99, -30, 18, -82, -107,
    -- layer=1 filter=231 channel=42
    -14, -23, -45, -10, -18, -49, -7, 1, 30,
    -- layer=1 filter=231 channel=43
    -89, -46, 0, -79, -73, -59, -28, -61, -85,
    -- layer=1 filter=231 channel=44
    -48, -25, 54, -2, -69, 5, 43, 10, -74,
    -- layer=1 filter=231 channel=45
    1, 6, 52, 1, -26, -10, 58, 8, -48,
    -- layer=1 filter=231 channel=46
    12, -31, -13, 57, 14, -56, 40, 45, 50,
    -- layer=1 filter=231 channel=47
    -39, -33, -60, -18, -51, -60, 10, -45, -6,
    -- layer=1 filter=231 channel=48
    21, 20, 3, -9, 20, 26, -12, -13, 35,
    -- layer=1 filter=231 channel=49
    -13, -23, -56, 8, -22, -35, 20, -1, 6,
    -- layer=1 filter=231 channel=50
    -1, 41, 0, 13, -4, 1, 20, 33, 12,
    -- layer=1 filter=231 channel=51
    28, 28, 5, 16, 55, 28, -28, 38, 44,
    -- layer=1 filter=231 channel=52
    -73, -67, -45, -38, 14, -9, -62, -54, -19,
    -- layer=1 filter=231 channel=53
    20, 6, 16, 13, 9, 16, 8, 13, -1,
    -- layer=1 filter=231 channel=54
    -88, -67, -4, -82, -22, -32, -88, -58, -4,
    -- layer=1 filter=231 channel=55
    -19, -24, 7, 7, -28, -3, 35, 5, -59,
    -- layer=1 filter=231 channel=56
    1, -5, 8, -6, -10, 6, 0, 1, 6,
    -- layer=1 filter=231 channel=57
    61, 66, 28, 18, 69, 80, -29, 39, 90,
    -- layer=1 filter=231 channel=58
    -10, 9, -16, -43, 3, 3, -40, -54, 56,
    -- layer=1 filter=231 channel=59
    1, -4, 6, -13, -4, -5, -10, 8, 10,
    -- layer=1 filter=231 channel=60
    0, 70, 20, 5, -23, -23, 0, 35, 3,
    -- layer=1 filter=231 channel=61
    -5, -2, -8, 2, 5, -5, 6, 7, 1,
    -- layer=1 filter=231 channel=62
    -100, -46, -12, -64, -85, -86, -14, -109, -138,
    -- layer=1 filter=231 channel=63
    13, 10, 11, -6, -20, -7, -33, -20, 11,
    -- layer=1 filter=231 channel=64
    -8, 0, 6, -5, 1, 0, -10, 0, 0,
    -- layer=1 filter=231 channel=65
    -10, 0, 1, 0, 19, 13, -10, 10, 11,
    -- layer=1 filter=231 channel=66
    -11, 3, 28, -18, -14, 32, -51, -16, -5,
    -- layer=1 filter=231 channel=67
    -43, -48, -52, -3, -24, -37, -4, -8, -7,
    -- layer=1 filter=231 channel=68
    -63, -60, 60, -49, -109, -24, 7, -46, -113,
    -- layer=1 filter=231 channel=69
    -3, 4, 74, 35, -35, -30, 81, 28, -76,
    -- layer=1 filter=231 channel=70
    14, 10, -65, 52, 4, -21, -5, 32, 37,
    -- layer=1 filter=231 channel=71
    19, 8, 3, 34, 6, -17, 34, 35, 14,
    -- layer=1 filter=231 channel=72
    32, -6, 5, -15, -9, -15, 32, 3, 5,
    -- layer=1 filter=231 channel=73
    7, 4, -11, 7, -4, 3, -25, 4, 5,
    -- layer=1 filter=231 channel=74
    -26, -52, -12, -36, -67, -30, -60, -58, -3,
    -- layer=1 filter=231 channel=75
    105, 56, -1, 76, 84, 40, 29, 85, 117,
    -- layer=1 filter=231 channel=76
    -30, -8, 41, -35, -56, -7, -7, -54, -21,
    -- layer=1 filter=231 channel=77
    8, 11, 12, -2, 1, 32, 20, -13, 29,
    -- layer=1 filter=231 channel=78
    1, -11, 23, -24, -4, 37, -40, 0, 40,
    -- layer=1 filter=231 channel=79
    -73, -34, -19, -49, -76, -84, 5, -79, -119,
    -- layer=1 filter=231 channel=80
    11, -7, -2, 2, 10, 5, -49, 20, -5,
    -- layer=1 filter=231 channel=81
    15, 0, 24, 2, -12, 11, 32, -14, -1,
    -- layer=1 filter=231 channel=82
    14, -5, -3, 22, 14, -7, 17, 19, -9,
    -- layer=1 filter=231 channel=83
    3, 11, 54, 0, -13, 48, 53, 6, -38,
    -- layer=1 filter=231 channel=84
    -14, -10, -59, -19, -20, -9, -52, -79, 14,
    -- layer=1 filter=231 channel=85
    -49, -21, -34, -97, -65, -34, 4, -101, -9,
    -- layer=1 filter=231 channel=86
    -16, 5, 17, -15, -10, 29, -35, -20, -12,
    -- layer=1 filter=231 channel=87
    -32, -94, -39, -12, -21, -39, 17, -8, -57,
    -- layer=1 filter=231 channel=88
    20, 8, -25, 18, -5, -36, 31, 13, -27,
    -- layer=1 filter=231 channel=89
    6, -9, -5, 19, 22, -10, 21, 22, 7,
    -- layer=1 filter=231 channel=90
    -25, -3, 76, -6, -42, 48, 56, 0, -57,
    -- layer=1 filter=231 channel=91
    25, 25, 9, 1, 30, 44, -11, 4, 40,
    -- layer=1 filter=231 channel=92
    -13, -11, 40, -8, 16, 13, 44, 28, -66,
    -- layer=1 filter=231 channel=93
    -7, 2, 23, -8, -6, 12, 2, -11, -17,
    -- layer=1 filter=231 channel=94
    13, 35, 19, -29, 13, 48, -85, -20, 17,
    -- layer=1 filter=231 channel=95
    35, 26, -33, 12, 12, 21, -28, -4, 52,
    -- layer=1 filter=231 channel=96
    10, 2, 7, 2, 9, 0, 1, -5, 3,
    -- layer=1 filter=231 channel=97
    -16, 23, 47, -45, -19, 26, -24, -38, -13,
    -- layer=1 filter=231 channel=98
    -34, 5, 29, -85, -46, -29, -4, -79, -86,
    -- layer=1 filter=231 channel=99
    37, 42, 66, -18, 41, 112, -57, 29, 56,
    -- layer=1 filter=231 channel=100
    -37, -26, -4, 8, -15, -13, 7, 5, -7,
    -- layer=1 filter=231 channel=101
    1, 6, -8, 15, 4, 12, -4, 17, 9,
    -- layer=1 filter=231 channel=102
    -4, 24, 12, -38, 2, 35, -85, -31, 28,
    -- layer=1 filter=231 channel=103
    -24, -20, 1, -8, 5, 7, 5, -33, -28,
    -- layer=1 filter=231 channel=104
    -24, 8, -26, -26, -17, -27, 20, -40, -10,
    -- layer=1 filter=231 channel=105
    0, 42, 41, -36, 10, 57, -62, -22, 28,
    -- layer=1 filter=231 channel=106
    -24, -35, -10, -20, -61, -37, 12, -13, -39,
    -- layer=1 filter=231 channel=107
    6, 10, 17, 4, -2, -9, 12, 1, 14,
    -- layer=1 filter=231 channel=108
    -28, -44, 10, 16, -78, 1, 69, 0, -136,
    -- layer=1 filter=231 channel=109
    10, 3, 11, 9, 0, -3, -5, -7, 11,
    -- layer=1 filter=231 channel=110
    20, 22, 9, -14, 7, 5, -34, -3, 17,
    -- layer=1 filter=231 channel=111
    70, 72, -20, 0, 49, 61, -31, 3, 104,
    -- layer=1 filter=231 channel=112
    1, 2, -18, 0, 0, 27, -72, -50, 7,
    -- layer=1 filter=231 channel=113
    -14, -2, -59, 15, 24, -43, 18, 47, -14,
    -- layer=1 filter=231 channel=114
    -23, -8, 29, 46, -44, -74, 25, 5, -85,
    -- layer=1 filter=231 channel=115
    22, 44, 16, -19, 37, 55, -73, -2, 34,
    -- layer=1 filter=231 channel=116
    0, 6, -4, 4, 10, 6, 0, -9, 3,
    -- layer=1 filter=231 channel=117
    74, 110, 10, 56, 75, 93, -87, 2, 99,
    -- layer=1 filter=231 channel=118
    11, -6, -32, -13, 5, 8, -21, -26, 38,
    -- layer=1 filter=231 channel=119
    -33, -38, 25, -19, -73, -23, 40, -32, -130,
    -- layer=1 filter=231 channel=120
    13, 23, 3, 4, 21, 34, -11, -9, 36,
    -- layer=1 filter=231 channel=121
    50, 34, 8, 61, 58, 36, 35, 67, 62,
    -- layer=1 filter=231 channel=122
    8, -6, -8, -3, -9, -7, -8, -9, 7,
    -- layer=1 filter=231 channel=123
    17, 23, 9, 37, 34, 25, 29, 44, 73,
    -- layer=1 filter=231 channel=124
    3, -12, -12, 4, -12, -6, 12, -7, -11,
    -- layer=1 filter=231 channel=125
    7, 20, -58, 25, 3, -38, -21, 9, 5,
    -- layer=1 filter=231 channel=126
    16, 11, 78, -35, -62, 45, 19, -82, -48,
    -- layer=1 filter=231 channel=127
    24, 12, -28, 13, 34, 23, -24, -17, 73,
    -- layer=1 filter=232 channel=0
    -4, 0, -5, -11, 3, 4, -9, -1, -5,
    -- layer=1 filter=232 channel=1
    1, -11, 5, -4, 6, 2, -6, 7, -1,
    -- layer=1 filter=232 channel=2
    5, -11, -3, -13, 4, 2, -12, 4, 2,
    -- layer=1 filter=232 channel=3
    10, 0, -6, 5, 2, -8, 10, -10, 1,
    -- layer=1 filter=232 channel=4
    -1, 3, -7, -10, 0, 0, 7, -4, 1,
    -- layer=1 filter=232 channel=5
    -14, -3, -8, 3, -1, -6, 7, -7, -10,
    -- layer=1 filter=232 channel=6
    -12, 5, 0, 3, -12, -4, -1, -11, 8,
    -- layer=1 filter=232 channel=7
    -6, -6, -7, 0, 2, -8, -12, 4, -1,
    -- layer=1 filter=232 channel=8
    -8, 0, 0, 7, -4, 3, -3, -5, -6,
    -- layer=1 filter=232 channel=9
    2, -1, -6, 0, 2, 4, 2, 2, 7,
    -- layer=1 filter=232 channel=10
    -2, 3, 3, -3, -11, -3, 2, 0, 0,
    -- layer=1 filter=232 channel=11
    -2, 3, -12, 7, -5, -6, -12, -4, 5,
    -- layer=1 filter=232 channel=12
    2, 7, -7, -8, 4, 4, 10, 8, 5,
    -- layer=1 filter=232 channel=13
    -2, 1, 7, -2, 7, -13, 6, -2, 0,
    -- layer=1 filter=232 channel=14
    -3, 3, -1, 0, 2, 2, 5, -6, -1,
    -- layer=1 filter=232 channel=15
    -2, -18, -9, 8, 4, 0, -2, -9, 2,
    -- layer=1 filter=232 channel=16
    -4, -7, -2, -1, -10, -10, 2, 3, -8,
    -- layer=1 filter=232 channel=17
    5, 0, -11, 2, -1, 6, -2, 1, 0,
    -- layer=1 filter=232 channel=18
    -6, -7, 4, 0, -12, -4, -2, -10, 1,
    -- layer=1 filter=232 channel=19
    3, 2, 3, -8, -8, 1, -9, 2, 1,
    -- layer=1 filter=232 channel=20
    6, -1, -4, 6, -7, 3, -12, 6, -10,
    -- layer=1 filter=232 channel=21
    -7, 1, 3, 2, -12, -9, 6, -4, 0,
    -- layer=1 filter=232 channel=22
    -1, 6, -7, -4, 0, -9, -6, -2, -6,
    -- layer=1 filter=232 channel=23
    -8, -3, 7, 8, -11, 8, -7, -11, 2,
    -- layer=1 filter=232 channel=24
    0, -8, -2, -2, -3, -1, 0, -12, 7,
    -- layer=1 filter=232 channel=25
    0, -4, -2, -8, -5, -2, -15, 0, 5,
    -- layer=1 filter=232 channel=26
    -3, -5, -13, 2, -10, -14, 0, 2, -11,
    -- layer=1 filter=232 channel=27
    10, 8, -11, 0, -2, 2, 7, 4, -3,
    -- layer=1 filter=232 channel=28
    -1, 7, 7, 0, 7, -6, 0, -10, -6,
    -- layer=1 filter=232 channel=29
    1, -9, 1, -1, 1, -4, -8, -4, -5,
    -- layer=1 filter=232 channel=30
    0, 0, -10, 4, -7, -3, 5, -9, -12,
    -- layer=1 filter=232 channel=31
    -6, 1, -14, -10, 3, 3, 5, 3, 0,
    -- layer=1 filter=232 channel=32
    -8, -7, -11, -6, -3, -5, 4, -3, 4,
    -- layer=1 filter=232 channel=33
    -6, 0, 1, 4, 3, 4, -3, 5, 9,
    -- layer=1 filter=232 channel=34
    1, -9, -2, -10, -10, 5, 1, 1, -8,
    -- layer=1 filter=232 channel=35
    -1, -5, -1, 0, 4, 2, -9, 0, 6,
    -- layer=1 filter=232 channel=36
    4, 3, -1, -9, -5, -7, 0, -9, 8,
    -- layer=1 filter=232 channel=37
    -6, -4, -3, 6, 6, 6, -9, -8, 3,
    -- layer=1 filter=232 channel=38
    -12, -1, -5, -3, -12, -7, -4, -8, 0,
    -- layer=1 filter=232 channel=39
    4, -2, 6, 5, 4, -6, -4, 1, -8,
    -- layer=1 filter=232 channel=40
    -4, -8, 4, 1, -1, -10, 0, 6, 4,
    -- layer=1 filter=232 channel=41
    -10, -8, 0, 0, -2, 5, -6, -1, 7,
    -- layer=1 filter=232 channel=42
    -5, 6, 1, -1, 0, -8, 0, 7, 0,
    -- layer=1 filter=232 channel=43
    8, -13, -8, -1, 6, -3, -4, 5, 6,
    -- layer=1 filter=232 channel=44
    -3, -6, 6, 4, -4, 0, -11, 5, -4,
    -- layer=1 filter=232 channel=45
    5, -5, 6, -4, 5, -4, -5, -9, 2,
    -- layer=1 filter=232 channel=46
    -17, 2, 0, -4, 7, 3, -1, 1, -5,
    -- layer=1 filter=232 channel=47
    -17, 0, -1, 0, -7, -8, 0, -3, -9,
    -- layer=1 filter=232 channel=48
    4, 6, -6, 2, -8, -6, 6, -9, -9,
    -- layer=1 filter=232 channel=49
    -9, 7, -3, 7, 0, 2, -8, 0, -5,
    -- layer=1 filter=232 channel=50
    -2, 7, 0, 2, -11, 0, -9, -1, 0,
    -- layer=1 filter=232 channel=51
    -4, 5, 5, -7, -6, 0, -9, -8, -3,
    -- layer=1 filter=232 channel=52
    11, -2, 10, -5, -9, -2, -1, -9, -5,
    -- layer=1 filter=232 channel=53
    -3, -1, -11, -5, -5, 7, 1, 0, -9,
    -- layer=1 filter=232 channel=54
    -11, 0, 1, -9, -7, -5, -8, -19, 8,
    -- layer=1 filter=232 channel=55
    -2, -8, -3, 4, -2, -14, -7, 6, -1,
    -- layer=1 filter=232 channel=56
    3, -8, 0, 7, 2, -6, 0, 7, 1,
    -- layer=1 filter=232 channel=57
    5, -14, 4, 1, 0, -7, -7, -11, 8,
    -- layer=1 filter=232 channel=58
    -2, -10, -10, 8, -12, 2, 6, -2, -5,
    -- layer=1 filter=232 channel=59
    0, -11, 8, -10, -5, -9, -11, 6, 6,
    -- layer=1 filter=232 channel=60
    -5, 0, -6, -5, -12, 9, 1, -2, -4,
    -- layer=1 filter=232 channel=61
    -8, -11, -7, 5, 4, -8, 1, -5, 4,
    -- layer=1 filter=232 channel=62
    0, -14, -6, -7, -10, -4, 4, -14, 3,
    -- layer=1 filter=232 channel=63
    6, -7, 7, -7, 5, 0, -10, 5, 0,
    -- layer=1 filter=232 channel=64
    6, -7, -4, 1, 8, -9, -7, -11, -11,
    -- layer=1 filter=232 channel=65
    -5, 4, 3, 0, -5, 4, -5, 3, 6,
    -- layer=1 filter=232 channel=66
    1, -11, -6, 3, 7, 1, -11, 3, 2,
    -- layer=1 filter=232 channel=67
    0, -5, 4, 0, 1, 10, 5, -1, -6,
    -- layer=1 filter=232 channel=68
    -16, -8, 4, -11, -9, -4, -6, -1, -1,
    -- layer=1 filter=232 channel=69
    -5, -1, 8, -9, 3, -5, -7, -12, -5,
    -- layer=1 filter=232 channel=70
    7, -7, 6, -2, -7, -6, -8, -12, -2,
    -- layer=1 filter=232 channel=71
    -5, 0, -4, 6, -4, 2, 4, -6, -2,
    -- layer=1 filter=232 channel=72
    -10, -5, 0, -3, 2, -6, 0, -9, 5,
    -- layer=1 filter=232 channel=73
    -10, 0, -2, -10, 1, -5, 4, 1, 5,
    -- layer=1 filter=232 channel=74
    6, 0, 7, 7, 1, -5, 5, 5, -1,
    -- layer=1 filter=232 channel=75
    1, 4, -1, -6, 0, -4, -4, -2, -4,
    -- layer=1 filter=232 channel=76
    -6, -4, -9, -9, 0, -8, -1, -7, -3,
    -- layer=1 filter=232 channel=77
    -11, -2, 4, -2, 7, -2, -4, 0, 5,
    -- layer=1 filter=232 channel=78
    4, 5, 6, -9, 1, 5, 7, 5, -6,
    -- layer=1 filter=232 channel=79
    4, 2, -7, -9, -1, 2, -14, -1, 0,
    -- layer=1 filter=232 channel=80
    -7, -4, 6, 7, -8, 2, 0, 10, 10,
    -- layer=1 filter=232 channel=81
    5, -5, -6, 7, 4, 3, -12, -1, -4,
    -- layer=1 filter=232 channel=82
    2, 0, 8, 0, -9, -10, -2, -10, 2,
    -- layer=1 filter=232 channel=83
    4, -2, -6, -7, 7, -4, 6, -8, 1,
    -- layer=1 filter=232 channel=84
    6, 4, -5, -6, -2, -3, 6, -7, -9,
    -- layer=1 filter=232 channel=85
    0, 1, 0, -12, 1, -11, 6, 6, -8,
    -- layer=1 filter=232 channel=86
    -8, -14, -13, -5, 0, -9, 4, -9, -3,
    -- layer=1 filter=232 channel=87
    -11, -2, 1, -2, -2, 4, -4, 2, 6,
    -- layer=1 filter=232 channel=88
    -4, -4, -7, -4, -5, 4, -6, -9, -4,
    -- layer=1 filter=232 channel=89
    -3, 2, -3, 4, -10, -4, -11, -11, -10,
    -- layer=1 filter=232 channel=90
    -7, -9, 1, -5, 7, 4, 3, -1, -5,
    -- layer=1 filter=232 channel=91
    4, -8, -1, 0, 1, -2, 3, 5, -12,
    -- layer=1 filter=232 channel=92
    3, 2, -10, -4, 8, -2, 5, 6, 6,
    -- layer=1 filter=232 channel=93
    7, -8, 7, 5, -7, -4, 7, 4, -10,
    -- layer=1 filter=232 channel=94
    -1, 8, 2, -11, 6, 5, 2, -10, -9,
    -- layer=1 filter=232 channel=95
    9, -2, -4, -5, -5, -10, 6, -11, 1,
    -- layer=1 filter=232 channel=96
    -4, -1, 2, 2, -11, -2, -9, -2, 2,
    -- layer=1 filter=232 channel=97
    1, 6, -9, 0, -2, -3, -2, -10, -8,
    -- layer=1 filter=232 channel=98
    -7, -6, 4, 3, 6, 1, 4, -13, 1,
    -- layer=1 filter=232 channel=99
    3, -9, 0, -4, -7, 6, 8, -9, 2,
    -- layer=1 filter=232 channel=100
    -1, -8, 4, 2, 3, 5, -11, -4, 0,
    -- layer=1 filter=232 channel=101
    4, -5, -6, 0, -6, 7, 4, -4, -8,
    -- layer=1 filter=232 channel=102
    7, -4, -11, 7, -11, 2, 1, -10, 6,
    -- layer=1 filter=232 channel=103
    7, -1, 0, -9, -11, -2, -5, -7, -12,
    -- layer=1 filter=232 channel=104
    3, 5, -6, 3, -11, 5, -7, 6, -5,
    -- layer=1 filter=232 channel=105
    3, -1, -5, 3, 8, 2, -12, 4, -11,
    -- layer=1 filter=232 channel=106
    -3, 5, -13, 0, -5, -9, 4, 3, -13,
    -- layer=1 filter=232 channel=107
    -3, -10, 3, -2, -5, -10, -9, 4, -6,
    -- layer=1 filter=232 channel=108
    -12, -8, -14, -10, -3, -14, -8, -4, -1,
    -- layer=1 filter=232 channel=109
    -7, -5, 6, 7, 1, 7, -8, 3, 0,
    -- layer=1 filter=232 channel=110
    0, -11, -8, -9, -8, -2, -3, 5, -7,
    -- layer=1 filter=232 channel=111
    6, 0, 0, -2, -5, -6, 1, -6, 0,
    -- layer=1 filter=232 channel=112
    -7, 0, 8, 7, -5, -6, -9, 5, -9,
    -- layer=1 filter=232 channel=113
    -13, -11, 0, -5, 4, 5, -4, 5, -5,
    -- layer=1 filter=232 channel=114
    -11, 1, -10, -8, -7, -8, 4, -1, 1,
    -- layer=1 filter=232 channel=115
    -2, -2, 1, -7, 3, -10, -7, -5, -7,
    -- layer=1 filter=232 channel=116
    -2, -2, -3, -5, 9, 2, 2, -7, 6,
    -- layer=1 filter=232 channel=117
    -2, 0, 4, 0, -7, 1, -1, -6, 3,
    -- layer=1 filter=232 channel=118
    -2, 8, -3, -1, -10, 7, -5, -6, -1,
    -- layer=1 filter=232 channel=119
    -1, -8, 0, -1, -4, -7, -7, 0, 5,
    -- layer=1 filter=232 channel=120
    -6, -16, -4, -12, 5, -14, 1, -9, -4,
    -- layer=1 filter=232 channel=121
    8, -2, -11, 0, -10, -5, -13, 0, -4,
    -- layer=1 filter=232 channel=122
    2, -3, -4, -6, 5, -2, 3, -10, -5,
    -- layer=1 filter=232 channel=123
    -7, -11, -5, 3, 2, -1, -7, -4, -9,
    -- layer=1 filter=232 channel=124
    6, 0, 1, 4, -10, 6, -7, -5, 11,
    -- layer=1 filter=232 channel=125
    0, -8, -12, 7, -10, 0, -8, -8, -7,
    -- layer=1 filter=232 channel=126
    -3, 7, -9, 0, -2, -2, 7, 5, -11,
    -- layer=1 filter=232 channel=127
    -11, -10, 0, -2, -19, 7, 5, -10, -5,
    -- layer=1 filter=233 channel=0
    1, 5, 8, 8, -6, 8, -8, 1, -6,
    -- layer=1 filter=233 channel=1
    6, 7, 1, -11, -4, 2, 0, -4, 1,
    -- layer=1 filter=233 channel=2
    1, 7, -5, -2, -4, -10, 1, -10, 7,
    -- layer=1 filter=233 channel=3
    -10, 3, -1, -9, 3, 11, -4, -3, 2,
    -- layer=1 filter=233 channel=4
    -6, 4, 7, -1, 4, -7, -8, 4, 4,
    -- layer=1 filter=233 channel=5
    5, 5, 2, -7, -4, -7, 3, -7, -4,
    -- layer=1 filter=233 channel=6
    -5, -6, 4, 1, 0, -1, 6, -9, -10,
    -- layer=1 filter=233 channel=7
    3, -2, 5, -5, -7, 5, -8, -5, -5,
    -- layer=1 filter=233 channel=8
    2, 0, -8, -11, -9, -5, -4, -2, -7,
    -- layer=1 filter=233 channel=9
    -2, -7, -1, 5, -10, 0, -5, 1, -10,
    -- layer=1 filter=233 channel=10
    -3, 5, 2, -5, 9, -9, 0, 9, 4,
    -- layer=1 filter=233 channel=11
    -5, 8, -7, 7, 8, 0, 3, -3, -1,
    -- layer=1 filter=233 channel=12
    -2, 1, 3, -7, -10, -8, -10, -2, 0,
    -- layer=1 filter=233 channel=13
    -9, -4, -7, 2, 7, 7, 0, 3, 6,
    -- layer=1 filter=233 channel=14
    -1, 9, 2, -5, -10, -4, 2, 7, 5,
    -- layer=1 filter=233 channel=15
    -3, -4, 0, -8, -11, -6, 0, 1, 0,
    -- layer=1 filter=233 channel=16
    -5, 4, -2, 10, 0, 11, -9, -9, 6,
    -- layer=1 filter=233 channel=17
    0, -6, 7, -2, -3, 6, -8, -5, -8,
    -- layer=1 filter=233 channel=18
    -4, 6, -11, 7, 4, -2, 4, 0, -7,
    -- layer=1 filter=233 channel=19
    -10, -3, -5, 0, -5, -6, 3, 7, 2,
    -- layer=1 filter=233 channel=20
    -1, -9, -3, 6, 4, -11, 3, -11, 1,
    -- layer=1 filter=233 channel=21
    -9, -11, 4, -11, -1, -12, -3, 0, -9,
    -- layer=1 filter=233 channel=22
    -9, -3, 11, -1, -8, -10, 0, 7, -11,
    -- layer=1 filter=233 channel=23
    3, -5, 5, 1, 0, 0, 7, -3, -9,
    -- layer=1 filter=233 channel=24
    5, -8, -2, -5, 4, -1, -7, 1, -6,
    -- layer=1 filter=233 channel=25
    -5, 0, -5, 2, 7, -1, -5, 9, 0,
    -- layer=1 filter=233 channel=26
    -6, -8, 0, 1, -1, -8, -6, 7, 5,
    -- layer=1 filter=233 channel=27
    10, 11, 0, 0, -3, -6, -6, 3, -4,
    -- layer=1 filter=233 channel=28
    -4, -5, 7, -9, -8, 0, -8, 6, 1,
    -- layer=1 filter=233 channel=29
    -1, -2, -8, 0, 3, 0, -6, -3, 0,
    -- layer=1 filter=233 channel=30
    2, 3, 9, -11, 3, -5, -4, -3, 1,
    -- layer=1 filter=233 channel=31
    -4, -7, 0, -5, -7, 5, 6, 0, -6,
    -- layer=1 filter=233 channel=32
    4, -4, -1, -1, 0, 5, 0, -3, -7,
    -- layer=1 filter=233 channel=33
    -8, -5, -4, -4, 7, -6, 0, 1, 5,
    -- layer=1 filter=233 channel=34
    1, -3, 2, -3, 0, -1, -3, -3, 3,
    -- layer=1 filter=233 channel=35
    4, -4, 0, -3, -5, 7, -10, 8, 1,
    -- layer=1 filter=233 channel=36
    -7, -9, 7, 0, -1, -10, -11, 4, 5,
    -- layer=1 filter=233 channel=37
    -3, -9, -8, -4, 5, -9, 0, 5, -1,
    -- layer=1 filter=233 channel=38
    -7, -2, -10, -2, 6, 6, -10, 3, -1,
    -- layer=1 filter=233 channel=39
    -5, -10, 8, -12, 2, 8, -9, -11, -11,
    -- layer=1 filter=233 channel=40
    9, -2, -8, -3, -9, 5, -3, 9, 0,
    -- layer=1 filter=233 channel=41
    0, 7, -3, -1, -6, -7, 1, 1, 6,
    -- layer=1 filter=233 channel=42
    1, -12, 4, 7, 6, -13, -3, 0, -7,
    -- layer=1 filter=233 channel=43
    0, -3, 8, -5, -5, -6, -3, -2, -9,
    -- layer=1 filter=233 channel=44
    0, -5, -1, 2, 2, 8, 1, 6, 3,
    -- layer=1 filter=233 channel=45
    -1, 0, -10, -2, -9, 7, -3, -11, -2,
    -- layer=1 filter=233 channel=46
    10, -2, 9, 5, -2, 9, 3, -3, 1,
    -- layer=1 filter=233 channel=47
    -7, 0, -5, 0, 4, -10, -7, -9, -4,
    -- layer=1 filter=233 channel=48
    5, -7, 3, 5, 6, -6, 0, -6, -5,
    -- layer=1 filter=233 channel=49
    4, -4, -6, -2, 5, 5, 2, 5, 3,
    -- layer=1 filter=233 channel=50
    -9, 0, 0, -8, -7, 2, -1, 2, -9,
    -- layer=1 filter=233 channel=51
    -7, -10, -12, 6, -8, -5, -8, 7, 2,
    -- layer=1 filter=233 channel=52
    4, -9, -8, -7, -3, 0, 2, 7, 0,
    -- layer=1 filter=233 channel=53
    5, -11, -11, 0, 7, 1, -10, -7, 5,
    -- layer=1 filter=233 channel=54
    -7, 4, 8, 10, -8, 4, -6, -7, -2,
    -- layer=1 filter=233 channel=55
    0, 5, 0, 2, 4, -11, 3, -4, -4,
    -- layer=1 filter=233 channel=56
    -1, 8, -1, 5, -4, -11, -5, 5, 1,
    -- layer=1 filter=233 channel=57
    -5, 6, -3, -4, -9, -3, 0, -6, 2,
    -- layer=1 filter=233 channel=58
    0, -8, -10, 5, -6, -3, 7, 7, 0,
    -- layer=1 filter=233 channel=59
    -11, 2, -5, 7, -9, 4, -10, -10, -1,
    -- layer=1 filter=233 channel=60
    -3, -9, -2, 5, 3, 1, 1, 6, 0,
    -- layer=1 filter=233 channel=61
    5, 5, -6, -6, 0, -6, 9, 10, 2,
    -- layer=1 filter=233 channel=62
    -10, -5, -1, -3, 0, 3, 5, -10, 0,
    -- layer=1 filter=233 channel=63
    -1, 6, -4, 8, -3, -11, 7, -6, -7,
    -- layer=1 filter=233 channel=64
    -2, -12, 2, 6, 0, -10, -8, -3, -1,
    -- layer=1 filter=233 channel=65
    -1, -7, -7, 7, 5, -3, 1, 5, -5,
    -- layer=1 filter=233 channel=66
    0, 8, 4, -9, -10, -11, 8, -8, -3,
    -- layer=1 filter=233 channel=67
    10, -8, -3, 2, 4, 8, 0, 2, 0,
    -- layer=1 filter=233 channel=68
    -8, 0, -4, -2, 0, 0, 5, 0, 0,
    -- layer=1 filter=233 channel=69
    3, 5, 1, 6, 5, 8, -6, -6, 1,
    -- layer=1 filter=233 channel=70
    -11, 1, -4, -2, 2, -5, 1, 0, -4,
    -- layer=1 filter=233 channel=71
    -8, -6, -2, 1, -4, -3, -8, 1, -8,
    -- layer=1 filter=233 channel=72
    -1, 7, 5, -4, 2, -11, -10, 2, -10,
    -- layer=1 filter=233 channel=73
    2, -5, 6, 2, 0, -6, 2, 3, -6,
    -- layer=1 filter=233 channel=74
    -2, 8, -11, 6, -11, -11, 8, 0, 1,
    -- layer=1 filter=233 channel=75
    -7, -6, -2, 8, -8, 10, -10, 1, 7,
    -- layer=1 filter=233 channel=76
    -8, -3, 7, 2, 5, 1, -10, 7, -7,
    -- layer=1 filter=233 channel=77
    -4, -5, 3, 7, 4, 0, 3, -10, -1,
    -- layer=1 filter=233 channel=78
    -11, -4, -9, -6, 0, -3, 1, 4, 6,
    -- layer=1 filter=233 channel=79
    -9, -4, 11, -11, -7, -7, 3, -1, 6,
    -- layer=1 filter=233 channel=80
    -5, 0, 2, 6, 5, 5, -2, 5, -8,
    -- layer=1 filter=233 channel=81
    3, 4, -3, -2, 3, -2, -11, -7, -2,
    -- layer=1 filter=233 channel=82
    -9, -3, 5, -6, 3, -1, -8, -4, -3,
    -- layer=1 filter=233 channel=83
    5, 5, -3, -7, 2, -11, 8, -3, -11,
    -- layer=1 filter=233 channel=84
    0, -7, -3, 0, -10, -11, -3, -8, -2,
    -- layer=1 filter=233 channel=85
    3, 0, 7, -3, -8, 4, 4, -9, 1,
    -- layer=1 filter=233 channel=86
    -6, -2, 9, 8, -7, 4, -4, -7, -5,
    -- layer=1 filter=233 channel=87
    -6, -5, 0, -6, -3, -2, 2, -1, -11,
    -- layer=1 filter=233 channel=88
    -9, -2, 0, -11, 8, 1, 6, -5, -10,
    -- layer=1 filter=233 channel=89
    1, 8, 5, 0, 2, 0, -7, -10, -9,
    -- layer=1 filter=233 channel=90
    -12, -10, -4, -3, -5, 3, -8, -3, 5,
    -- layer=1 filter=233 channel=91
    0, 0, -4, -5, 7, 5, 4, 2, 5,
    -- layer=1 filter=233 channel=92
    3, 0, -3, 7, 8, 8, 8, -1, 0,
    -- layer=1 filter=233 channel=93
    4, -11, 0, 7, 6, 0, 0, 0, -11,
    -- layer=1 filter=233 channel=94
    -6, 7, -1, 6, -11, -11, 3, 1, -8,
    -- layer=1 filter=233 channel=95
    3, 0, -8, 1, 7, 6, -4, -3, -2,
    -- layer=1 filter=233 channel=96
    7, 0, -3, -5, 8, 1, 8, -7, 8,
    -- layer=1 filter=233 channel=97
    2, 0, -10, 0, -7, -8, -8, -10, -9,
    -- layer=1 filter=233 channel=98
    -3, -9, -7, -4, -1, 10, 6, -3, -2,
    -- layer=1 filter=233 channel=99
    -10, -1, 7, 8, -2, 3, -10, 3, -8,
    -- layer=1 filter=233 channel=100
    -8, -7, -5, -2, 4, -6, -9, 5, -7,
    -- layer=1 filter=233 channel=101
    -5, 7, -3, 1, -6, -7, -9, 6, 6,
    -- layer=1 filter=233 channel=102
    1, -8, 1, 1, -9, -5, -3, -10, -8,
    -- layer=1 filter=233 channel=103
    -1, -5, -9, 0, 8, 2, 7, 0, 0,
    -- layer=1 filter=233 channel=104
    0, 3, -4, -12, 3, -11, -2, 5, -10,
    -- layer=1 filter=233 channel=105
    1, -7, 2, 2, -9, -1, 4, -1, 4,
    -- layer=1 filter=233 channel=106
    -6, -8, -10, -11, 3, -3, 1, -3, -4,
    -- layer=1 filter=233 channel=107
    0, -5, 8, -11, 0, -7, 1, 7, 7,
    -- layer=1 filter=233 channel=108
    -11, -7, 2, 0, 4, -6, -6, -7, -2,
    -- layer=1 filter=233 channel=109
    -9, -7, 0, -9, -6, -5, 0, 6, -7,
    -- layer=1 filter=233 channel=110
    -7, -4, 8, -6, 2, 0, -11, -9, 5,
    -- layer=1 filter=233 channel=111
    0, -8, -3, -9, -5, 0, 4, 6, -9,
    -- layer=1 filter=233 channel=112
    3, -3, 5, 3, 0, 4, 1, -2, -10,
    -- layer=1 filter=233 channel=113
    9, -3, -4, -7, -1, 2, 2, -7, -2,
    -- layer=1 filter=233 channel=114
    0, 4, -7, 4, -8, 5, -1, 8, -10,
    -- layer=1 filter=233 channel=115
    -11, -3, 0, 3, 7, -8, 3, 4, -2,
    -- layer=1 filter=233 channel=116
    -4, -5, 6, 0, 7, 4, 6, -7, 9,
    -- layer=1 filter=233 channel=117
    6, -8, -10, 1, 5, -1, 0, 2, 8,
    -- layer=1 filter=233 channel=118
    1, -2, 8, -8, -3, -2, 5, 1, 7,
    -- layer=1 filter=233 channel=119
    -7, -4, -2, 0, -6, 5, 1, -9, 5,
    -- layer=1 filter=233 channel=120
    0, -9, -6, 2, -11, -6, -4, -10, 7,
    -- layer=1 filter=233 channel=121
    -8, 3, 6, 7, 3, -10, -3, -11, -7,
    -- layer=1 filter=233 channel=122
    10, -5, -4, 6, 6, -6, 7, 3, -2,
    -- layer=1 filter=233 channel=123
    -10, -8, -9, 0, -12, 3, -10, 3, -7,
    -- layer=1 filter=233 channel=124
    3, 4, 11, 9, -9, 0, -4, -4, 1,
    -- layer=1 filter=233 channel=125
    -10, -1, -1, 2, 6, 0, 8, 9, -7,
    -- layer=1 filter=233 channel=126
    -8, 7, -4, -7, 1, -7, -6, 4, -3,
    -- layer=1 filter=233 channel=127
    7, 9, 6, 4, -4, -6, -6, 8, -6,
    -- layer=1 filter=234 channel=0
    -9, 3, -4, -8, 5, 0, -5, -2, 0,
    -- layer=1 filter=234 channel=1
    -4, -1, -6, 0, 0, -7, -9, -1, -4,
    -- layer=1 filter=234 channel=2
    -10, -2, -13, -11, -3, -2, 6, 6, -1,
    -- layer=1 filter=234 channel=3
    -1, 9, -8, -3, 6, -9, 0, 2, 7,
    -- layer=1 filter=234 channel=4
    -7, -2, 2, -1, 3, -8, 6, -9, -5,
    -- layer=1 filter=234 channel=5
    -9, 1, -3, 0, 1, 6, -4, 12, -4,
    -- layer=1 filter=234 channel=6
    0, -9, -2, 5, -6, -11, 0, 4, -1,
    -- layer=1 filter=234 channel=7
    -4, -10, -1, -6, 6, 6, -5, -2, -6,
    -- layer=1 filter=234 channel=8
    -11, -12, 5, 0, 2, 6, -5, 2, -2,
    -- layer=1 filter=234 channel=9
    2, 10, 6, -8, -3, 3, 6, -6, -5,
    -- layer=1 filter=234 channel=10
    3, -3, -4, -2, -9, -1, -11, -3, -3,
    -- layer=1 filter=234 channel=11
    -2, 10, 10, 8, 5, -7, 1, 10, 8,
    -- layer=1 filter=234 channel=12
    8, 7, 0, -1, 6, -4, -5, -9, 6,
    -- layer=1 filter=234 channel=13
    -8, -6, -2, 0, -3, -4, 7, 1, 5,
    -- layer=1 filter=234 channel=14
    -2, 13, -8, -2, -10, 7, -7, -2, 5,
    -- layer=1 filter=234 channel=15
    -7, -4, 9, 10, -1, -5, -6, -10, 3,
    -- layer=1 filter=234 channel=16
    -9, 8, -12, 3, -8, 2, -5, -7, -9,
    -- layer=1 filter=234 channel=17
    -4, -8, -6, -6, 0, -5, -2, -2, 4,
    -- layer=1 filter=234 channel=18
    9, -3, -5, 0, -7, -3, -7, -12, 0,
    -- layer=1 filter=234 channel=19
    -3, 1, 4, 0, -1, -3, -7, 6, -3,
    -- layer=1 filter=234 channel=20
    -10, 4, 4, -7, -8, 0, 1, -9, 8,
    -- layer=1 filter=234 channel=21
    -10, 4, -7, -2, -9, -2, 2, 3, -12,
    -- layer=1 filter=234 channel=22
    -2, -5, -7, -7, 7, -1, -5, -9, 0,
    -- layer=1 filter=234 channel=23
    -10, -3, -2, -4, 5, 3, -7, -4, 0,
    -- layer=1 filter=234 channel=24
    -14, -4, -9, 1, -12, 5, -8, -7, 2,
    -- layer=1 filter=234 channel=25
    -5, 4, -13, 6, 0, -5, 1, -10, -8,
    -- layer=1 filter=234 channel=26
    3, -7, 2, -4, -3, 0, 1, -5, -1,
    -- layer=1 filter=234 channel=27
    8, -1, -2, 0, 7, -2, -10, -9, -6,
    -- layer=1 filter=234 channel=28
    -5, -3, -8, -7, 7, 6, 1, -2, 2,
    -- layer=1 filter=234 channel=29
    -4, -5, 5, 8, -9, 7, 1, 1, -5,
    -- layer=1 filter=234 channel=30
    0, -4, -6, 4, 0, -8, -1, -1, -3,
    -- layer=1 filter=234 channel=31
    -1, -3, -3, -8, 5, 4, 0, 4, -12,
    -- layer=1 filter=234 channel=32
    0, 8, 6, -3, -9, -3, -6, 3, -7,
    -- layer=1 filter=234 channel=33
    -3, 1, -1, -6, 11, -4, -9, 0, 7,
    -- layer=1 filter=234 channel=34
    0, 0, 0, -10, 4, 0, -6, 5, -3,
    -- layer=1 filter=234 channel=35
    0, -4, 0, -6, 6, -1, 7, 0, 8,
    -- layer=1 filter=234 channel=36
    0, 1, -7, -1, -2, -5, 3, 4, 3,
    -- layer=1 filter=234 channel=37
    3, -1, 0, 3, -3, 0, -5, -7, -1,
    -- layer=1 filter=234 channel=38
    5, -2, 4, -7, -8, 5, 4, -12, -2,
    -- layer=1 filter=234 channel=39
    -11, -3, 0, -9, 3, -3, -6, 3, -11,
    -- layer=1 filter=234 channel=40
    -7, -6, -6, 3, -7, -2, 7, -4, -8,
    -- layer=1 filter=234 channel=41
    -9, 2, 7, 0, -4, -11, -7, -3, -10,
    -- layer=1 filter=234 channel=42
    5, 2, -7, -12, 7, 0, -10, -10, -7,
    -- layer=1 filter=234 channel=43
    -8, -3, -2, 3, -1, -11, 0, 6, 2,
    -- layer=1 filter=234 channel=44
    -3, -6, -11, 1, 7, 6, -12, 0, 6,
    -- layer=1 filter=234 channel=45
    5, -3, 2, 2, 4, -5, -2, 6, 6,
    -- layer=1 filter=234 channel=46
    -3, 0, -8, 10, 5, 1, 4, -9, 5,
    -- layer=1 filter=234 channel=47
    -8, -3, -9, -1, 4, 0, -3, 5, -3,
    -- layer=1 filter=234 channel=48
    -5, 3, 6, -8, -11, -7, -7, 2, -9,
    -- layer=1 filter=234 channel=49
    0, -10, -8, -10, -12, 1, -10, 3, -3,
    -- layer=1 filter=234 channel=50
    -2, -11, 5, 7, -1, 6, -2, 4, -4,
    -- layer=1 filter=234 channel=51
    -8, 0, -3, -8, -2, 5, 0, -9, 8,
    -- layer=1 filter=234 channel=52
    -8, -3, 2, 1, -3, 10, -8, 2, -4,
    -- layer=1 filter=234 channel=53
    -5, -3, 6, 7, 4, -4, -8, -11, 0,
    -- layer=1 filter=234 channel=54
    6, 7, 7, -1, -9, -2, -12, 1, 5,
    -- layer=1 filter=234 channel=55
    3, -2, -8, -8, 4, 0, 1, -6, 0,
    -- layer=1 filter=234 channel=56
    2, 0, -7, 8, 5, 7, 1, -9, 7,
    -- layer=1 filter=234 channel=57
    3, -10, 6, -8, -4, -11, 5, 9, -1,
    -- layer=1 filter=234 channel=58
    8, 5, 5, -12, 2, 1, 7, 2, 0,
    -- layer=1 filter=234 channel=59
    7, 7, 8, 6, -4, 4, -6, -9, -7,
    -- layer=1 filter=234 channel=60
    5, -3, 1, -10, 6, 4, 0, 7, -6,
    -- layer=1 filter=234 channel=61
    0, -7, -7, 1, -1, -6, 6, -1, 9,
    -- layer=1 filter=234 channel=62
    -5, -9, -7, 9, -8, -8, 6, -8, 0,
    -- layer=1 filter=234 channel=63
    7, -9, -7, -9, -1, -3, 8, 8, 5,
    -- layer=1 filter=234 channel=64
    -10, -10, -6, 8, -10, 3, 3, -7, 4,
    -- layer=1 filter=234 channel=65
    1, 1, -6, -5, 8, -11, 0, 2, -11,
    -- layer=1 filter=234 channel=66
    0, 0, -4, 6, -8, -5, -7, 8, -4,
    -- layer=1 filter=234 channel=67
    -8, -1, 4, -1, 0, 0, -5, -9, -5,
    -- layer=1 filter=234 channel=68
    -11, -4, -2, 6, -6, 0, -2, 4, 0,
    -- layer=1 filter=234 channel=69
    -3, 7, -11, 0, -5, 5, -6, 3, 6,
    -- layer=1 filter=234 channel=70
    3, 6, 2, -8, -5, 8, -1, -1, -8,
    -- layer=1 filter=234 channel=71
    2, -5, -11, -11, 6, 3, -12, 6, 0,
    -- layer=1 filter=234 channel=72
    -10, -7, 4, -1, 6, 5, -6, -6, -9,
    -- layer=1 filter=234 channel=73
    -2, 8, 3, 11, 0, -10, 5, -8, -5,
    -- layer=1 filter=234 channel=74
    6, -5, 4, -10, -6, -6, 2, 0, 2,
    -- layer=1 filter=234 channel=75
    2, -14, 1, 3, 3, 5, -2, -6, -3,
    -- layer=1 filter=234 channel=76
    4, -11, 6, 7, 5, -8, 0, -9, 2,
    -- layer=1 filter=234 channel=77
    -10, 3, -3, 4, -7, 6, 6, 0, -10,
    -- layer=1 filter=234 channel=78
    -10, -10, 1, -8, 2, -3, -6, -2, -1,
    -- layer=1 filter=234 channel=79
    0, -11, -6, -2, 5, 7, 7, -5, -9,
    -- layer=1 filter=234 channel=80
    1, -2, 7, -2, -5, -7, -2, 3, 3,
    -- layer=1 filter=234 channel=81
    0, -9, 1, -5, -2, 8, 0, 6, -8,
    -- layer=1 filter=234 channel=82
    1, 1, -5, -4, -11, 2, 2, -12, -2,
    -- layer=1 filter=234 channel=83
    -5, 5, -6, -2, 0, -10, 7, 8, 2,
    -- layer=1 filter=234 channel=84
    2, -9, -5, 0, -10, 11, 1, -2, 8,
    -- layer=1 filter=234 channel=85
    -3, -2, -8, 2, -12, 0, 1, -2, 2,
    -- layer=1 filter=234 channel=86
    5, -6, 7, -6, 8, -8, 3, 0, -8,
    -- layer=1 filter=234 channel=87
    -9, 8, -1, -9, 9, 2, -3, -8, 3,
    -- layer=1 filter=234 channel=88
    10, 2, -2, 3, -4, -14, -10, 6, 8,
    -- layer=1 filter=234 channel=89
    1, 6, -1, -6, 4, -8, 6, -9, -4,
    -- layer=1 filter=234 channel=90
    5, -10, 6, 4, -3, 4, 8, -2, 2,
    -- layer=1 filter=234 channel=91
    -5, 7, -2, 6, -8, 4, 7, -4, 1,
    -- layer=1 filter=234 channel=92
    0, 7, 1, 3, -2, 0, -8, -2, -4,
    -- layer=1 filter=234 channel=93
    -4, 7, -10, -11, 1, -3, 0, 2, -4,
    -- layer=1 filter=234 channel=94
    6, -2, -3, -10, -3, -2, -7, 0, 3,
    -- layer=1 filter=234 channel=95
    0, -11, 0, 7, 11, -3, -4, -10, -1,
    -- layer=1 filter=234 channel=96
    1, -11, -2, 4, 8, -4, -8, -4, 0,
    -- layer=1 filter=234 channel=97
    -2, -10, 3, -4, 3, 4, 6, 7, -3,
    -- layer=1 filter=234 channel=98
    -8, 2, -3, -8, 0, -10, -9, -5, 5,
    -- layer=1 filter=234 channel=99
    4, -4, -9, 3, 6, -9, 6, 3, 0,
    -- layer=1 filter=234 channel=100
    0, 7, 4, 1, 4, -4, -9, -1, -11,
    -- layer=1 filter=234 channel=101
    -2, 6, -11, -2, 7, -10, 8, -1, 1,
    -- layer=1 filter=234 channel=102
    0, -3, 5, -5, 3, 5, 3, 4, 8,
    -- layer=1 filter=234 channel=103
    3, -5, 2, -1, 0, -5, 0, 0, 8,
    -- layer=1 filter=234 channel=104
    0, 6, 2, -10, -9, -11, -12, -6, 0,
    -- layer=1 filter=234 channel=105
    -3, -3, -8, -6, 5, -12, 7, 2, -1,
    -- layer=1 filter=234 channel=106
    -1, -2, -7, -12, -4, -7, -6, 4, 7,
    -- layer=1 filter=234 channel=107
    2, -6, -4, 2, 8, 4, 6, 0, 4,
    -- layer=1 filter=234 channel=108
    3, -4, -13, 2, 0, -10, -2, -9, -5,
    -- layer=1 filter=234 channel=109
    6, -11, -8, -5, -8, -4, 9, -4, 6,
    -- layer=1 filter=234 channel=110
    -9, 0, -4, 7, -5, -2, -7, 1, -8,
    -- layer=1 filter=234 channel=111
    4, -3, -5, 1, 7, -6, -10, -6, -6,
    -- layer=1 filter=234 channel=112
    3, 6, 7, -5, 0, -3, 1, -9, -1,
    -- layer=1 filter=234 channel=113
    5, -9, -4, 0, 10, -1, -6, -10, 4,
    -- layer=1 filter=234 channel=114
    3, -1, -1, 0, -13, -2, 2, 9, -3,
    -- layer=1 filter=234 channel=115
    -1, 7, 0, -4, -6, -3, -3, -5, 4,
    -- layer=1 filter=234 channel=116
    -3, 0, -8, -6, -9, 0, 7, 6, -2,
    -- layer=1 filter=234 channel=117
    -9, -9, 7, 1, -2, -6, 9, -11, 0,
    -- layer=1 filter=234 channel=118
    -4, 8, 0, 6, -1, 2, 2, -4, 0,
    -- layer=1 filter=234 channel=119
    -4, 0, -12, 8, 0, -7, -1, -9, 0,
    -- layer=1 filter=234 channel=120
    -1, 0, 4, 7, -6, 5, -7, -6, -2,
    -- layer=1 filter=234 channel=121
    -15, -7, 1, 0, 3, 4, 7, 5, -5,
    -- layer=1 filter=234 channel=122
    -4, 9, -8, -2, 2, 1, 10, 4, 1,
    -- layer=1 filter=234 channel=123
    -6, 6, 0, 10, 4, -9, 2, -3, -3,
    -- layer=1 filter=234 channel=124
    -2, 0, 3, -9, 0, -7, -9, 2, 7,
    -- layer=1 filter=234 channel=125
    3, -6, 2, -7, 7, 4, -10, 7, 10,
    -- layer=1 filter=234 channel=126
    7, -6, -12, -8, -1, -3, 8, 6, -4,
    -- layer=1 filter=234 channel=127
    -5, -11, -10, 1, 0, 10, 0, 0, -1,
    -- layer=1 filter=235 channel=0
    -1, -6, -6, -11, 2, -12, -5, 7, -2,
    -- layer=1 filter=235 channel=1
    0, 4, 0, -10, -5, 5, 7, -4, -4,
    -- layer=1 filter=235 channel=2
    1, 3, -10, 8, -6, 9, -8, 3, 5,
    -- layer=1 filter=235 channel=3
    -6, 9, 11, -9, -7, -5, 6, -2, 8,
    -- layer=1 filter=235 channel=4
    -12, 5, 6, -4, 5, 7, -6, 4, -3,
    -- layer=1 filter=235 channel=5
    -9, -5, -7, 5, -3, 8, -11, -9, 0,
    -- layer=1 filter=235 channel=6
    0, 3, -7, -4, -4, 8, -4, -8, 0,
    -- layer=1 filter=235 channel=7
    -4, -11, 6, 0, 6, 1, -9, -7, 4,
    -- layer=1 filter=235 channel=8
    -5, 0, -1, -10, 3, -10, 7, 0, 0,
    -- layer=1 filter=235 channel=9
    -9, -9, 8, -8, -2, 1, -3, -8, -11,
    -- layer=1 filter=235 channel=10
    -2, 9, -10, -6, 0, -9, -9, -3, 0,
    -- layer=1 filter=235 channel=11
    -8, 2, -4, -9, -9, 8, 3, 7, -5,
    -- layer=1 filter=235 channel=12
    -8, 9, 6, 0, 6, -8, 7, 1, -2,
    -- layer=1 filter=235 channel=13
    -10, -5, -2, 0, -8, 5, -10, 3, -2,
    -- layer=1 filter=235 channel=14
    7, 1, -2, -9, 5, -8, -3, 6, 10,
    -- layer=1 filter=235 channel=15
    -1, 5, -7, 0, -8, 4, 3, -7, -6,
    -- layer=1 filter=235 channel=16
    -5, -6, -6, 4, 8, 3, -1, 7, -7,
    -- layer=1 filter=235 channel=17
    3, -2, -7, 2, 3, -1, -6, 5, 6,
    -- layer=1 filter=235 channel=18
    2, 6, -4, -2, 2, -1, 9, 4, -3,
    -- layer=1 filter=235 channel=19
    3, 2, 6, -12, 8, 2, -5, 6, 3,
    -- layer=1 filter=235 channel=20
    1, -1, -10, -11, -7, -7, 0, 2, 7,
    -- layer=1 filter=235 channel=21
    4, 0, -7, 0, 5, 8, -2, -7, 8,
    -- layer=1 filter=235 channel=22
    -7, 5, 2, 0, 3, -4, -4, -1, 8,
    -- layer=1 filter=235 channel=23
    -1, -6, 6, 8, 3, 4, -2, -2, 1,
    -- layer=1 filter=235 channel=24
    9, -7, -9, -5, 2, -3, 0, -2, 4,
    -- layer=1 filter=235 channel=25
    0, -5, -6, 1, 12, -2, -3, 2, 3,
    -- layer=1 filter=235 channel=26
    7, -9, 0, 4, 11, -3, 6, -8, -11,
    -- layer=1 filter=235 channel=27
    1, 4, -8, 11, 0, 0, 1, 0, -6,
    -- layer=1 filter=235 channel=28
    -8, -7, 0, 7, 0, 8, -9, 0, -9,
    -- layer=1 filter=235 channel=29
    -6, 7, -3, 0, -3, 1, 4, 9, -2,
    -- layer=1 filter=235 channel=30
    7, -4, 11, 3, 6, -2, 2, -6, -2,
    -- layer=1 filter=235 channel=31
    -6, -5, 0, -10, -5, -2, -6, 4, -3,
    -- layer=1 filter=235 channel=32
    -8, 0, 4, 6, -4, -5, -2, -3, 2,
    -- layer=1 filter=235 channel=33
    -5, 8, -7, 1, 0, -7, 4, 1, -4,
    -- layer=1 filter=235 channel=34
    0, -4, 4, -9, -3, 0, -4, -7, 2,
    -- layer=1 filter=235 channel=35
    3, 4, -11, -3, 3, -10, 3, -9, 1,
    -- layer=1 filter=235 channel=36
    1, -10, 0, 0, -8, -10, 7, 4, 3,
    -- layer=1 filter=235 channel=37
    5, 0, 9, -6, -8, -11, -5, 0, 7,
    -- layer=1 filter=235 channel=38
    4, 5, 3, -8, 2, -9, -9, -9, 0,
    -- layer=1 filter=235 channel=39
    -8, -10, -4, -10, -10, 7, -4, 3, -4,
    -- layer=1 filter=235 channel=40
    -4, -8, 0, -11, 9, -4, -9, 9, -7,
    -- layer=1 filter=235 channel=41
    -6, -3, 0, -11, 5, 0, -9, -3, -5,
    -- layer=1 filter=235 channel=42
    8, -10, -10, 9, 8, -6, -10, 8, 3,
    -- layer=1 filter=235 channel=43
    -10, 5, 2, -6, 0, -1, -8, -4, -2,
    -- layer=1 filter=235 channel=44
    -4, 7, -4, -10, -2, 1, 3, -10, -1,
    -- layer=1 filter=235 channel=45
    -6, 4, -4, -4, -5, -8, -4, -4, 0,
    -- layer=1 filter=235 channel=46
    5, -6, -6, 8, -1, 8, -4, 7, 1,
    -- layer=1 filter=235 channel=47
    -9, 1, 0, -3, 7, 10, 0, -2, -5,
    -- layer=1 filter=235 channel=48
    -4, -11, -7, -9, 6, -6, 0, 0, -11,
    -- layer=1 filter=235 channel=49
    0, -6, -6, -3, 0, -3, -1, 9, -2,
    -- layer=1 filter=235 channel=50
    -6, -10, -7, -6, -3, -8, -4, -11, 3,
    -- layer=1 filter=235 channel=51
    -7, 0, -4, 0, 5, 8, -6, 8, 0,
    -- layer=1 filter=235 channel=52
    4, 1, 0, -2, 9, -1, 4, -3, 0,
    -- layer=1 filter=235 channel=53
    0, -3, -1, -6, 6, 0, -4, 7, 3,
    -- layer=1 filter=235 channel=54
    -5, 3, -4, -4, 2, -10, -1, -2, 8,
    -- layer=1 filter=235 channel=55
    -7, 7, -7, 2, 2, 7, -1, 9, 11,
    -- layer=1 filter=235 channel=56
    -2, -4, -2, 2, -2, -10, -4, 5, 1,
    -- layer=1 filter=235 channel=57
    -3, -4, -4, -8, 7, -3, 2, 6, -2,
    -- layer=1 filter=235 channel=58
    3, 10, -2, 8, -5, -6, -8, 10, 7,
    -- layer=1 filter=235 channel=59
    1, 2, -11, -2, -1, 4, -10, 7, 2,
    -- layer=1 filter=235 channel=60
    -3, -1, 10, -7, 5, 3, -2, -6, 4,
    -- layer=1 filter=235 channel=61
    3, 0, 9, -8, 4, -5, -1, 0, 1,
    -- layer=1 filter=235 channel=62
    0, 3, 1, -5, 0, 0, -9, 0, -3,
    -- layer=1 filter=235 channel=63
    -5, -10, 8, -8, 1, -2, -8, -7, -10,
    -- layer=1 filter=235 channel=64
    5, 0, 8, 5, -8, -8, -2, -3, 7,
    -- layer=1 filter=235 channel=65
    2, 2, -4, -5, -4, 6, 0, -4, -8,
    -- layer=1 filter=235 channel=66
    0, 0, -5, -2, -1, 2, 7, 3, -9,
    -- layer=1 filter=235 channel=67
    4, -1, -3, 1, -8, -4, -3, -3, 0,
    -- layer=1 filter=235 channel=68
    2, 4, -5, 8, 7, 3, -5, -4, -5,
    -- layer=1 filter=235 channel=69
    2, -5, 8, -5, -1, 1, -4, -3, -8,
    -- layer=1 filter=235 channel=70
    -1, -11, -4, 3, -1, -2, 8, 4, 0,
    -- layer=1 filter=235 channel=71
    5, -10, 2, 7, 4, 4, 5, -4, 2,
    -- layer=1 filter=235 channel=72
    -3, 1, -10, -8, -1, -1, -4, -11, 4,
    -- layer=1 filter=235 channel=73
    8, 3, -11, -10, -4, -4, -4, 3, 8,
    -- layer=1 filter=235 channel=74
    -2, 4, -9, 2, -5, -4, 6, -8, 3,
    -- layer=1 filter=235 channel=75
    -9, -10, -4, -1, 0, 1, -7, -5, -3,
    -- layer=1 filter=235 channel=76
    6, 7, 6, 5, 0, -12, 1, 3, -10,
    -- layer=1 filter=235 channel=77
    -5, -10, 0, -1, 3, 3, 0, -5, 0,
    -- layer=1 filter=235 channel=78
    -10, -10, 0, 1, 6, -10, 3, -8, -6,
    -- layer=1 filter=235 channel=79
    6, -11, 5, 6, -10, -2, -3, 5, -9,
    -- layer=1 filter=235 channel=80
    6, 5, 4, 9, -5, 0, -1, -7, -6,
    -- layer=1 filter=235 channel=81
    -10, -9, -1, 8, -4, -6, 0, 1, -5,
    -- layer=1 filter=235 channel=82
    -6, -2, -12, 8, -1, -4, 4, 7, 8,
    -- layer=1 filter=235 channel=83
    -5, -10, 0, 2, 6, 1, 4, -9, -3,
    -- layer=1 filter=235 channel=84
    -7, -10, -10, -4, -5, -8, 3, -11, -7,
    -- layer=1 filter=235 channel=85
    -12, -9, -5, 6, -4, 8, -12, -4, -11,
    -- layer=1 filter=235 channel=86
    -6, 0, -1, 7, 6, -5, -6, -6, -6,
    -- layer=1 filter=235 channel=87
    -10, -4, 0, 4, 4, -3, 4, -1, 0,
    -- layer=1 filter=235 channel=88
    -8, 7, -6, -1, -8, 0, -2, -10, -6,
    -- layer=1 filter=235 channel=89
    0, 6, 0, -8, 2, 7, -11, 1, -10,
    -- layer=1 filter=235 channel=90
    8, -10, -8, -9, -6, 2, -2, 4, -4,
    -- layer=1 filter=235 channel=91
    -6, 1, -10, -11, 0, 3, -6, 0, 2,
    -- layer=1 filter=235 channel=92
    1, -5, -10, -5, 0, -1, -8, 0, 2,
    -- layer=1 filter=235 channel=93
    -3, -6, 0, -5, -4, 0, 3, -11, 2,
    -- layer=1 filter=235 channel=94
    -8, -4, -4, -3, 1, 4, 8, 5, -1,
    -- layer=1 filter=235 channel=95
    -4, 3, -2, -7, -1, -6, 7, -9, 6,
    -- layer=1 filter=235 channel=96
    1, -10, -8, 2, -1, -6, -5, 6, -1,
    -- layer=1 filter=235 channel=97
    4, 0, -5, -10, -9, 0, 0, 5, 8,
    -- layer=1 filter=235 channel=98
    -9, 8, -2, -2, -1, -2, -7, 7, 8,
    -- layer=1 filter=235 channel=99
    -3, -12, -9, 1, -9, 7, 5, -7, -11,
    -- layer=1 filter=235 channel=100
    -4, -8, 4, 1, -9, 1, -11, 0, -11,
    -- layer=1 filter=235 channel=101
    7, -6, -1, -5, -7, 7, 5, -3, 2,
    -- layer=1 filter=235 channel=102
    -1, -4, 3, 6, -4, -5, -8, 7, -10,
    -- layer=1 filter=235 channel=103
    -3, -8, 7, 7, -4, -8, 0, -1, -8,
    -- layer=1 filter=235 channel=104
    2, -2, -5, 5, 5, -2, 0, -3, 1,
    -- layer=1 filter=235 channel=105
    1, -7, 0, 3, 1, 3, -5, -11, -1,
    -- layer=1 filter=235 channel=106
    6, 9, 5, -8, -8, -10, -2, 6, 0,
    -- layer=1 filter=235 channel=107
    -6, -8, -11, -1, 2, 1, -3, 1, 1,
    -- layer=1 filter=235 channel=108
    -8, -1, -6, 5, -1, 0, -2, -6, 11,
    -- layer=1 filter=235 channel=109
    0, -7, -7, -1, 4, 6, -1, -1, 1,
    -- layer=1 filter=235 channel=110
    -6, -1, -6, -7, -10, 1, -4, 3, -2,
    -- layer=1 filter=235 channel=111
    -1, -1, 5, -3, 9, 3, -6, -10, 6,
    -- layer=1 filter=235 channel=112
    1, 6, -10, 3, 5, 4, -8, -10, 7,
    -- layer=1 filter=235 channel=113
    -1, 3, -9, 0, 0, 8, 7, 0, -7,
    -- layer=1 filter=235 channel=114
    1, -5, 10, 0, 4, 2, -4, -7, -5,
    -- layer=1 filter=235 channel=115
    -6, -6, -8, 2, -7, -10, 0, -2, 2,
    -- layer=1 filter=235 channel=116
    5, -4, 6, -6, 4, -5, 6, 0, 9,
    -- layer=1 filter=235 channel=117
    -4, -5, -3, 7, 3, 0, 4, -1, 1,
    -- layer=1 filter=235 channel=118
    8, 9, -8, -4, 2, -4, -7, 0, -5,
    -- layer=1 filter=235 channel=119
    6, -2, -7, 8, 7, -1, -4, 1, -10,
    -- layer=1 filter=235 channel=120
    -9, 4, -11, 0, 0, -3, -3, -9, -7,
    -- layer=1 filter=235 channel=121
    -8, 0, 7, -2, -8, 6, 2, -8, 7,
    -- layer=1 filter=235 channel=122
    -7, -8, 4, -3, 9, 9, -7, -6, -2,
    -- layer=1 filter=235 channel=123
    5, 6, 1, -9, 3, -11, 4, 0, 1,
    -- layer=1 filter=235 channel=124
    -5, -9, 4, -10, 1, -3, 0, -11, 1,
    -- layer=1 filter=235 channel=125
    0, 8, -9, 0, -8, -8, -7, 0, -6,
    -- layer=1 filter=235 channel=126
    5, -6, -2, 0, -12, 2, 7, -5, 0,
    -- layer=1 filter=235 channel=127
    10, -1, 11, -2, -9, -4, 2, 2, -8,
    -- layer=1 filter=236 channel=0
    10, 10, 6, -5, -10, 0, 5, -9, -13,
    -- layer=1 filter=236 channel=1
    -4, -11, 20, 3, -9, -18, 8, 11, -11,
    -- layer=1 filter=236 channel=2
    -11, -28, -15, 22, -25, -1, 22, -9, 12,
    -- layer=1 filter=236 channel=3
    10, -13, -10, -9, -10, 0, 11, -9, 5,
    -- layer=1 filter=236 channel=4
    3, -1, 9, 6, 9, -9, 5, -4, -7,
    -- layer=1 filter=236 channel=5
    -6, -1, 17, 14, -21, -12, 2, 9, -7,
    -- layer=1 filter=236 channel=6
    -2, -14, -7, -11, -4, 3, -4, -8, -17,
    -- layer=1 filter=236 channel=7
    -2, -9, 16, 12, -12, 0, 2, -14, 15,
    -- layer=1 filter=236 channel=8
    -7, -10, 8, 16, -5, -16, 11, 22, 4,
    -- layer=1 filter=236 channel=9
    40, 20, -21, 8, -33, -9, -15, -8, -24,
    -- layer=1 filter=236 channel=10
    5, -12, 10, 22, -9, 0, 0, 6, 11,
    -- layer=1 filter=236 channel=11
    -7, -8, 5, -25, -13, 15, -15, 3, -12,
    -- layer=1 filter=236 channel=12
    -14, -14, -45, -6, -26, -4, -15, -2, 19,
    -- layer=1 filter=236 channel=13
    -7, 0, -11, 8, -3, 14, 3, 10, -14,
    -- layer=1 filter=236 channel=14
    -21, -22, 6, 7, 8, 0, 4, -8, -1,
    -- layer=1 filter=236 channel=15
    -5, 3, 1, -24, -33, -12, 19, 6, -2,
    -- layer=1 filter=236 channel=16
    0, 6, 11, -2, -23, -24, 13, 14, -3,
    -- layer=1 filter=236 channel=17
    -8, 13, 4, -12, -12, -15, 5, -10, -11,
    -- layer=1 filter=236 channel=18
    4, -15, 8, -5, 0, 26, 11, 2, 0,
    -- layer=1 filter=236 channel=19
    80, 109, 34, 61, 44, 33, 35, 55, 36,
    -- layer=1 filter=236 channel=20
    -7, 12, 9, 0, 0, 5, -2, 4, -8,
    -- layer=1 filter=236 channel=21
    2, -10, 3, 0, -4, -31, 7, -9, -11,
    -- layer=1 filter=236 channel=22
    -12, -9, 12, 0, 3, -13, 14, -1, -11,
    -- layer=1 filter=236 channel=23
    -1, 5, 16, -18, -44, -14, -9, -17, 25,
    -- layer=1 filter=236 channel=24
    19, 10, -8, -5, -34, -21, -12, -11, -10,
    -- layer=1 filter=236 channel=25
    14, 15, 19, 24, -3, -15, 7, 9, 15,
    -- layer=1 filter=236 channel=26
    3, 7, -15, 2, -19, 17, -8, 18, -9,
    -- layer=1 filter=236 channel=27
    42, 29, 28, 0, 13, 17, -20, -24, 3,
    -- layer=1 filter=236 channel=28
    10, 6, 32, 12, 10, -22, -19, 1, -11,
    -- layer=1 filter=236 channel=29
    29, 12, 18, -14, -15, -18, -19, -30, 2,
    -- layer=1 filter=236 channel=30
    15, -1, 13, 30, 10, 35, 23, 31, -5,
    -- layer=1 filter=236 channel=31
    -6, -14, 4, -12, -2, 15, -3, -5, -14,
    -- layer=1 filter=236 channel=32
    0, -10, -16, 12, -5, 15, 7, 9, 6,
    -- layer=1 filter=236 channel=33
    2, 16, 11, 7, 9, 13, 2, -8, -2,
    -- layer=1 filter=236 channel=34
    -2, -2, 10, 6, 4, -14, 11, 2, -12,
    -- layer=1 filter=236 channel=35
    4, 6, 0, 9, -2, -11, 5, 4, 3,
    -- layer=1 filter=236 channel=36
    -5, 12, 0, -14, -11, 6, -19, -11, -24,
    -- layer=1 filter=236 channel=37
    -2, 20, 9, 27, -5, -12, -1, 11, 9,
    -- layer=1 filter=236 channel=38
    -7, 6, 0, 12, 10, 8, -8, -14, -15,
    -- layer=1 filter=236 channel=39
    -5, 0, 3, 0, -17, -18, -24, -12, -16,
    -- layer=1 filter=236 channel=40
    -9, -13, 13, 8, 17, 27, 16, 9, -19,
    -- layer=1 filter=236 channel=41
    23, 13, -50, 41, -26, 23, -4, 20, -14,
    -- layer=1 filter=236 channel=42
    -44, -15, -19, -7, -9, -13, 7, 5, -5,
    -- layer=1 filter=236 channel=43
    -10, 12, 7, 1, -30, -48, 20, 23, 6,
    -- layer=1 filter=236 channel=44
    5, 1, -2, -4, -14, 17, -2, 16, -2,
    -- layer=1 filter=236 channel=45
    -5, 2, 0, 0, -22, -7, -1, 4, -1,
    -- layer=1 filter=236 channel=46
    74, 80, 55, 50, 22, 6, 26, 15, 40,
    -- layer=1 filter=236 channel=47
    -8, -15, -7, 21, -25, 20, 16, 2, 26,
    -- layer=1 filter=236 channel=48
    8, -2, -12, 3, -10, -2, 5, -22, -17,
    -- layer=1 filter=236 channel=49
    1, 0, -11, 1, -4, 3, 4, 0, -11,
    -- layer=1 filter=236 channel=50
    -4, 3, -4, -9, -1, -8, -7, -15, -17,
    -- layer=1 filter=236 channel=51
    4, -5, -1, 0, -6, 5, -2, -4, -1,
    -- layer=1 filter=236 channel=52
    8, -5, 7, -8, -9, -2, 4, 16, 19,
    -- layer=1 filter=236 channel=53
    6, 0, -12, -9, -21, -4, -21, 5, 13,
    -- layer=1 filter=236 channel=54
    20, 18, 15, 5, 2, -21, 4, 14, 6,
    -- layer=1 filter=236 channel=55
    0, -6, 0, -11, -11, 0, -4, -11, 4,
    -- layer=1 filter=236 channel=56
    1, -1, 0, 5, -5, -2, -9, -2, -5,
    -- layer=1 filter=236 channel=57
    0, -8, 7, 21, 16, -1, -5, 14, 15,
    -- layer=1 filter=236 channel=58
    17, 3, 9, 25, -16, 20, 3, -2, 40,
    -- layer=1 filter=236 channel=59
    10, 8, 3, -10, -9, -7, 1, 12, -11,
    -- layer=1 filter=236 channel=60
    23, 18, 4, 11, 12, 9, 5, 4, 5,
    -- layer=1 filter=236 channel=61
    -5, 0, -7, 11, -6, 14, 8, 14, -10,
    -- layer=1 filter=236 channel=62
    10, 32, 21, 11, -10, -18, 13, 16, 13,
    -- layer=1 filter=236 channel=63
    8, -1, 14, -6, -4, 9, -10, -5, -29,
    -- layer=1 filter=236 channel=64
    -10, -3, -7, -10, 3, -11, -13, -20, -6,
    -- layer=1 filter=236 channel=65
    9, -3, 3, -4, -10, -3, 9, -20, -15,
    -- layer=1 filter=236 channel=66
    -3, 18, 14, -5, -3, 1, -19, -18, -14,
    -- layer=1 filter=236 channel=67
    23, -3, -12, 11, -15, 0, -4, -23, 5,
    -- layer=1 filter=236 channel=68
    -2, 0, 3, 1, -6, 12, -7, 13, 16,
    -- layer=1 filter=236 channel=69
    1, -7, 2, -5, -30, -10, 8, 17, 16,
    -- layer=1 filter=236 channel=70
    9, -24, 0, -10, 5, 6, -4, 0, 12,
    -- layer=1 filter=236 channel=71
    8, 16, 13, 2, -9, -35, -6, -18, 2,
    -- layer=1 filter=236 channel=72
    38, 29, -14, 48, -2, 27, 20, 24, 13,
    -- layer=1 filter=236 channel=73
    5, -5, 4, -1, -7, -3, -14, 0, -17,
    -- layer=1 filter=236 channel=74
    14, -26, -12, -6, -5, 4, -6, 9, 1,
    -- layer=1 filter=236 channel=75
    -9, -25, 0, -15, -7, -9, 9, -10, -2,
    -- layer=1 filter=236 channel=76
    7, 0, 7, -13, -5, 12, -7, -6, -22,
    -- layer=1 filter=236 channel=77
    2, 3, 0, -13, -11, -27, 10, -6, -17,
    -- layer=1 filter=236 channel=78
    8, -3, 10, -5, 9, 1, -15, -4, -9,
    -- layer=1 filter=236 channel=79
    -11, 19, 21, 13, -27, -13, 17, 2, -2,
    -- layer=1 filter=236 channel=80
    10, -1, 3, 2, -7, -13, 8, -3, -2,
    -- layer=1 filter=236 channel=81
    18, 28, 8, -20, -34, -29, 0, -18, -3,
    -- layer=1 filter=236 channel=82
    -1, -4, -10, -17, -3, -23, -10, -24, -4,
    -- layer=1 filter=236 channel=83
    -4, -10, -5, 7, -16, -5, -9, 14, 6,
    -- layer=1 filter=236 channel=84
    24, 5, 4, 7, 18, 52, 34, 22, 5,
    -- layer=1 filter=236 channel=85
    9, 32, -4, 22, -31, -9, -10, -4, 2,
    -- layer=1 filter=236 channel=86
    3, 0, 21, -16, 0, -7, -21, -21, -15,
    -- layer=1 filter=236 channel=87
    71, 70, -12, 50, 1, -1, 2, 27, 26,
    -- layer=1 filter=236 channel=88
    -8, -6, -1, -4, -2, -2, 5, -13, -23,
    -- layer=1 filter=236 channel=89
    -4, 4, -6, 4, -12, -9, -7, -5, -21,
    -- layer=1 filter=236 channel=90
    -12, 0, -10, -7, -17, 5, 8, 31, 7,
    -- layer=1 filter=236 channel=91
    0, -1, -10, 0, 9, 17, 8, -7, 0,
    -- layer=1 filter=236 channel=92
    -14, -22, 0, -14, -54, 18, -22, 22, 28,
    -- layer=1 filter=236 channel=93
    0, 12, 3, -5, -17, -21, -11, -19, -18,
    -- layer=1 filter=236 channel=94
    10, 12, 20, -7, 12, 9, -11, -11, -14,
    -- layer=1 filter=236 channel=95
    13, -3, 25, 26, 34, 40, 27, 21, -9,
    -- layer=1 filter=236 channel=96
    3, 5, 12, -12, -10, -3, -16, -12, 0,
    -- layer=1 filter=236 channel=97
    12, 4, 13, -2, 0, -10, -18, -17, -4,
    -- layer=1 filter=236 channel=98
    0, 5, 9, 9, -17, -29, 19, 21, 23,
    -- layer=1 filter=236 channel=99
    2, -10, -4, -1, 9, -3, -5, 19, -8,
    -- layer=1 filter=236 channel=100
    13, -3, 0, -8, -11, 13, -10, -6, -17,
    -- layer=1 filter=236 channel=101
    0, -9, -2, -5, 0, 3, 1, -15, -8,
    -- layer=1 filter=236 channel=102
    2, 3, 3, 4, 14, 7, -3, -21, -14,
    -- layer=1 filter=236 channel=103
    0, 10, 2, -4, 3, 9, -6, -9, -3,
    -- layer=1 filter=236 channel=104
    2, -1, -5, 18, -24, 0, 3, 4, 21,
    -- layer=1 filter=236 channel=105
    13, 1, 16, -12, -10, -4, -11, -21, -15,
    -- layer=1 filter=236 channel=106
    -1, -12, -12, -7, 14, 15, 7, 3, -15,
    -- layer=1 filter=236 channel=107
    -7, -14, -17, -8, -29, -12, -13, -2, -6,
    -- layer=1 filter=236 channel=108
    -4, -14, -8, 2, -21, -11, 3, 20, -6,
    -- layer=1 filter=236 channel=109
    -4, -12, 7, 0, -6, 10, 4, 5, 5,
    -- layer=1 filter=236 channel=110
    7, 0, 8, 0, -10, -11, 0, 0, -2,
    -- layer=1 filter=236 channel=111
    17, -29, 5, 7, 2, 45, 15, 7, -21,
    -- layer=1 filter=236 channel=112
    -2, -24, 0, -18, 22, 4, 5, 17, 15,
    -- layer=1 filter=236 channel=113
    -21, -10, 20, -1, 3, -15, -25, -6, -28,
    -- layer=1 filter=236 channel=114
    -26, -9, 7, -16, -28, -11, 8, -10, -23,
    -- layer=1 filter=236 channel=115
    -4, 5, 21, -6, -14, -14, -22, -16, 1,
    -- layer=1 filter=236 channel=116
    -9, -4, -7, 3, -4, -3, 5, 7, -3,
    -- layer=1 filter=236 channel=117
    16, -37, 16, 14, 27, 48, 28, 28, 33,
    -- layer=1 filter=236 channel=118
    9, -13, 6, -5, 12, 14, 8, 25, -13,
    -- layer=1 filter=236 channel=119
    -1, 9, -4, 1, -17, 6, 14, 27, 9,
    -- layer=1 filter=236 channel=120
    -6, 2, -3, -4, -15, -24, 12, -1, 4,
    -- layer=1 filter=236 channel=121
    28, 29, 17, 6, 4, -6, -21, 11, -16,
    -- layer=1 filter=236 channel=122
    -4, -3, -4, 6, -2, -1, 1, 6, 4,
    -- layer=1 filter=236 channel=123
    8, 18, -9, -3, -9, -5, -19, -14, -20,
    -- layer=1 filter=236 channel=124
    0, 4, 0, 4, -10, 6, 8, 10, 10,
    -- layer=1 filter=236 channel=125
    -4, -28, -10, -10, 14, 7, -17, -5, -3,
    -- layer=1 filter=236 channel=126
    9, 7, -1, 26, 8, -8, 52, 34, 30,
    -- layer=1 filter=236 channel=127
    20, -5, 20, 13, 9, 31, 23, 37, 5,
    -- layer=1 filter=237 channel=0
    -36, -22, -39, 1, -13, -61, -14, -11, -38,
    -- layer=1 filter=237 channel=1
    21, -41, -54, -15, -21, -120, -57, -46, 50,
    -- layer=1 filter=237 channel=2
    2, 2, 16, 35, 55, 11, 31, 15, -44,
    -- layer=1 filter=237 channel=3
    1, -9, -1, 8, 5, -7, 2, -5, 8,
    -- layer=1 filter=237 channel=4
    16, 0, 13, 2, 6, 2, -7, -10, -11,
    -- layer=1 filter=237 channel=5
    -28, -38, -44, -18, -36, -51, 1, 0, 79,
    -- layer=1 filter=237 channel=6
    -27, -38, 20, -34, -41, -36, -27, -15, 3,
    -- layer=1 filter=237 channel=7
    1, -13, -8, -124, -39, 2, -53, -34, 120,
    -- layer=1 filter=237 channel=8
    2, -36, -70, -9, -37, -76, -30, -29, 65,
    -- layer=1 filter=237 channel=9
    -41, 2, 25, 10, -4, 33, 9, 25, -18,
    -- layer=1 filter=237 channel=10
    -31, -18, -24, -141, -35, -11, -27, -12, 133,
    -- layer=1 filter=237 channel=11
    -15, -2, -3, 15, 14, 0, 11, 13, 4,
    -- layer=1 filter=237 channel=12
    2, -21, 34, -13, -12, -18, 11, -3, -28,
    -- layer=1 filter=237 channel=13
    -9, -5, -7, 10, -29, -9, 22, 5, -79,
    -- layer=1 filter=237 channel=14
    8, 41, 45, -71, 47, -53, -62, -63, 1,
    -- layer=1 filter=237 channel=15
    -6, -7, -11, 58, -29, -21, 7, 43, 6,
    -- layer=1 filter=237 channel=16
    -10, -23, -41, -18, -71, -27, -27, -21, 94,
    -- layer=1 filter=237 channel=17
    -47, -28, -43, -9, -21, -28, -36, -64, -16,
    -- layer=1 filter=237 channel=18
    -46, -1, 0, -38, -34, -27, -7, -23, -62,
    -- layer=1 filter=237 channel=19
    -94, -36, -13, -106, -56, 64, 27, 78, 110,
    -- layer=1 filter=237 channel=20
    -30, -39, -6, 0, -25, -27, -19, -26, 29,
    -- layer=1 filter=237 channel=21
    -11, -38, -9, -15, -9, -26, -65, -37, -8,
    -- layer=1 filter=237 channel=22
    -8, -14, -25, 3, -15, -35, -36, -41, 19,
    -- layer=1 filter=237 channel=23
    4, -46, 0, -12, -46, 77, -13, 0, 115,
    -- layer=1 filter=237 channel=24
    -20, -6, 9, 3, -7, 27, 11, 34, -3,
    -- layer=1 filter=237 channel=25
    -8, -23, -35, -121, -41, 0, -14, -24, 161,
    -- layer=1 filter=237 channel=26
    -29, -5, 34, 26, -47, -21, 15, 10, -69,
    -- layer=1 filter=237 channel=27
    2, 13, 22, 16, 36, 5, 16, 25, 5,
    -- layer=1 filter=237 channel=28
    -21, -2, -21, -151, -39, -25, -75, -51, 93,
    -- layer=1 filter=237 channel=29
    -8, 3, 17, -17, 22, -21, -15, 23, -1,
    -- layer=1 filter=237 channel=30
    -78, 7, -29, -87, -45, -16, -8, 1, -44,
    -- layer=1 filter=237 channel=31
    -7, 3, 26, -26, 6, -33, 12, 9, -39,
    -- layer=1 filter=237 channel=32
    -18, 1, 26, 0, -50, 3, 9, 8, -41,
    -- layer=1 filter=237 channel=33
    -24, -10, -32, -23, -38, -2, -15, 0, 23,
    -- layer=1 filter=237 channel=34
    1, 9, 18, -2, -25, 7, -4, -1, 21,
    -- layer=1 filter=237 channel=35
    -4, -7, -1, 1, 2, -4, -6, -5, 6,
    -- layer=1 filter=237 channel=36
    -21, 7, -18, -10, -3, -24, 6, 10, -15,
    -- layer=1 filter=237 channel=37
    -56, -41, -49, -26, -40, -1, 1, 19, 111,
    -- layer=1 filter=237 channel=38
    -22, -19, 0, 1, -12, 1, 10, 1, -10,
    -- layer=1 filter=237 channel=39
    -24, -1, -14, 1, 5, -23, -23, -3, 34,
    -- layer=1 filter=237 channel=40
    -36, 7, 17, -29, 0, -31, 20, -8, 0,
    -- layer=1 filter=237 channel=41
    -31, 17, 50, -12, -46, 124, -9, 71, 10,
    -- layer=1 filter=237 channel=42
    6, 0, 3, 16, 45, 49, 37, 39, -28,
    -- layer=1 filter=237 channel=43
    -2, -39, -67, -46, -90, -43, -42, -21, 105,
    -- layer=1 filter=237 channel=44
    -18, -12, 14, 13, -35, -34, 20, 27, -52,
    -- layer=1 filter=237 channel=45
    0, -3, -2, 25, -3, -52, 10, 11, -26,
    -- layer=1 filter=237 channel=46
    -50, -20, 42, -41, -1, 37, 40, 103, 87,
    -- layer=1 filter=237 channel=47
    -3, -37, 22, 2, -32, 131, 9, 34, 46,
    -- layer=1 filter=237 channel=48
    -44, -31, -16, -29, -29, 16, 7, -25, 21,
    -- layer=1 filter=237 channel=49
    -9, -10, -11, -15, -14, 20, -9, 8, -46,
    -- layer=1 filter=237 channel=50
    -8, 15, -9, 17, 0, 0, 19, 44, 6,
    -- layer=1 filter=237 channel=51
    -42, -10, -11, -78, -23, -11, -39, -59, 99,
    -- layer=1 filter=237 channel=52
    -28, -14, 23, -55, -42, -43, -9, -5, -6,
    -- layer=1 filter=237 channel=53
    3, -4, -2, 3, 4, -9, -5, 0, -9,
    -- layer=1 filter=237 channel=54
    -42, -38, -30, -92, -26, 5, 20, 31, 195,
    -- layer=1 filter=237 channel=55
    3, 33, 28, 19, 14, 40, 18, 29, -5,
    -- layer=1 filter=237 channel=56
    0, -7, -8, 2, 8, -3, -3, 6, 2,
    -- layer=1 filter=237 channel=57
    -32, 7, -4, -92, -26, 14, -10, -8, 120,
    -- layer=1 filter=237 channel=58
    -6, -77, 4, -73, -83, 96, 15, 35, 146,
    -- layer=1 filter=237 channel=59
    -8, -3, 8, 4, -10, -7, -7, -3, 15,
    -- layer=1 filter=237 channel=60
    10, 10, 0, -31, -17, 4, 8, -30, -6,
    -- layer=1 filter=237 channel=61
    1, 8, 4, 6, -6, -7, -3, 3, -3,
    -- layer=1 filter=237 channel=62
    -35, -42, -43, -41, -86, -16, -34, -20, 116,
    -- layer=1 filter=237 channel=63
    -5, -1, 8, 1, 6, -7, 25, 14, -20,
    -- layer=1 filter=237 channel=64
    -31, -29, -2, -13, -2, -17, -17, -16, 20,
    -- layer=1 filter=237 channel=65
    -40, -33, -21, -28, -25, -40, -26, -66, 10,
    -- layer=1 filter=237 channel=66
    0, 11, -11, -1, 25, -18, -10, -15, 0,
    -- layer=1 filter=237 channel=67
    -6, 14, 28, -53, -21, 3, -12, -26, 0,
    -- layer=1 filter=237 channel=68
    -30, -7, 4, 30, -24, -25, 28, 7, -57,
    -- layer=1 filter=237 channel=69
    -12, 1, 21, 18, -33, -17, 7, 38, 44,
    -- layer=1 filter=237 channel=70
    -4, -3, 31, -20, -17, 0, -1, 23, 11,
    -- layer=1 filter=237 channel=71
    -10, -15, -4, -25, -6, -9, -25, 3, 54,
    -- layer=1 filter=237 channel=72
    -92, 14, -24, -84, -42, 29, -10, 46, -21,
    -- layer=1 filter=237 channel=73
    1, 1, -9, 0, -3, 6, -15, -7, 6,
    -- layer=1 filter=237 channel=74
    -4, -3, -24, -40, -20, -35, -10, -43, 12,
    -- layer=1 filter=237 channel=75
    -21, -7, 18, -35, 4, -20, -37, 0, -56,
    -- layer=1 filter=237 channel=76
    -39, -53, -15, -42, -35, -21, -6, -28, -8,
    -- layer=1 filter=237 channel=77
    -2, -14, -14, -23, -33, -41, -31, -37, -4,
    -- layer=1 filter=237 channel=78
    -4, -27, -46, -23, -23, -44, 12, -10, 52,
    -- layer=1 filter=237 channel=79
    -31, -39, -33, -26, -71, 14, -29, -1, 85,
    -- layer=1 filter=237 channel=80
    11, -1, 2, 5, 13, 15, -16, 0, 24,
    -- layer=1 filter=237 channel=81
    -15, -13, -24, -8, -35, 7, -21, 5, 37,
    -- layer=1 filter=237 channel=82
    -19, -21, -24, -13, -31, -27, -38, -24, -41,
    -- layer=1 filter=237 channel=83
    -13, 45, 2, 20, 2, -56, 6, 15, -36,
    -- layer=1 filter=237 channel=84
    -46, -11, -5, -22, -43, -39, 9, -30, -41,
    -- layer=1 filter=237 channel=85
    -30, -41, -47, -34, -68, 139, 5, 60, 123,
    -- layer=1 filter=237 channel=86
    14, 21, 0, -14, -15, -18, 6, 9, 15,
    -- layer=1 filter=237 channel=87
    -79, -18, 3, -40, -15, 76, 20, 84, 42,
    -- layer=1 filter=237 channel=88
    -4, 5, -15, -15, -21, 7, -1, -3, -27,
    -- layer=1 filter=237 channel=89
    -25, -36, -20, 4, -7, -71, -12, 12, -77,
    -- layer=1 filter=237 channel=90
    -15, 0, 37, 14, -37, -35, 19, 13, -63,
    -- layer=1 filter=237 channel=91
    -30, -9, 8, -14, -10, -4, 1, -25, 11,
    -- layer=1 filter=237 channel=92
    -8, -17, 41, 19, -20, -24, 17, 21, -59,
    -- layer=1 filter=237 channel=93
    -12, -45, -24, -11, -18, -35, -30, -29, 11,
    -- layer=1 filter=237 channel=94
    -23, -15, -48, -30, -24, -78, -16, -32, -49,
    -- layer=1 filter=237 channel=95
    -28, -25, -15, -74, -13, -37, -2, -41, -56,
    -- layer=1 filter=237 channel=96
    38, 30, 30, 26, 16, 15, 9, 5, 11,
    -- layer=1 filter=237 channel=97
    -26, -32, -48, -21, -22, -80, -25, -51, 21,
    -- layer=1 filter=237 channel=98
    0, -43, -73, -39, -95, -31, -63, -35, 92,
    -- layer=1 filter=237 channel=99
    -60, 12, -61, -117, -39, -85, -61, -61, 11,
    -- layer=1 filter=237 channel=100
    -11, 11, 12, 5, 20, 0, 30, 14, 4,
    -- layer=1 filter=237 channel=101
    -28, -34, -6, -12, -13, -22, -4, -12, -57,
    -- layer=1 filter=237 channel=102
    -47, -46, -48, -9, -25, -66, -24, -37, -48,
    -- layer=1 filter=237 channel=103
    10, 19, 7, 10, 29, 35, 22, 1, -6,
    -- layer=1 filter=237 channel=104
    -21, -26, -8, -34, -45, 69, -13, 1, 46,
    -- layer=1 filter=237 channel=105
    -46, -24, -50, -31, -31, -53, -17, -59, 28,
    -- layer=1 filter=237 channel=106
    -21, -28, 0, 23, -23, -41, 32, 16, -67,
    -- layer=1 filter=237 channel=107
    2, 7, -10, -10, -1, -10, -16, -18, -4,
    -- layer=1 filter=237 channel=108
    -26, -7, 28, 14, -30, 19, 5, -2, -53,
    -- layer=1 filter=237 channel=109
    4, 7, 0, 1, 6, -9, -2, -3, 7,
    -- layer=1 filter=237 channel=110
    -17, 7, -19, -22, 1, -5, -1, 3, -14,
    -- layer=1 filter=237 channel=111
    -55, 11, -12, -57, -44, -37, -17, -32, -65,
    -- layer=1 filter=237 channel=112
    -19, 1, 1, -51, 7, -52, 6, -23, -56,
    -- layer=1 filter=237 channel=113
    -7, 7, 6, 9, 19, 63, 10, 32, 53,
    -- layer=1 filter=237 channel=114
    -30, 0, -23, 14, -19, -43, -3, 43, 50,
    -- layer=1 filter=237 channel=115
    -12, 6, -13, -50, -24, -6, -21, -24, 74,
    -- layer=1 filter=237 channel=116
    8, -3, 7, 8, -6, -9, -8, 2, 3,
    -- layer=1 filter=237 channel=117
    -25, 0, 18, -104, -35, -106, 19, -108, -29,
    -- layer=1 filter=237 channel=118
    -53, -19, -20, -52, -62, -28, -3, -19, -64,
    -- layer=1 filter=237 channel=119
    -38, 18, 27, 0, -53, 33, 19, 17, -34,
    -- layer=1 filter=237 channel=120
    -16, -38, -30, -72, -47, 6, -38, -53, 101,
    -- layer=1 filter=237 channel=121
    -19, 4, 20, -22, 31, -3, 12, 42, -42,
    -- layer=1 filter=237 channel=122
    0, -9, 4, 5, 1, 7, 0, -3, 4,
    -- layer=1 filter=237 channel=123
    9, 16, 36, -19, 20, 42, 8, 50, 9,
    -- layer=1 filter=237 channel=124
    8, -5, 13, 15, -4, 7, 7, 2, 10,
    -- layer=1 filter=237 channel=125
    -10, 5, 21, -19, -22, 8, -26, 2, 57,
    -- layer=1 filter=237 channel=126
    16, -5, -59, 25, -27, -96, -61, -75, 44,
    -- layer=1 filter=237 channel=127
    -53, -15, -4, -67, -40, -49, -16, -19, -86,
    -- layer=1 filter=238 channel=0
    -6, -2, 7, 2, 10, -8, -12, -9, -12,
    -- layer=1 filter=238 channel=1
    0, 2, 0, -4, -10, -8, -7, 0, -2,
    -- layer=1 filter=238 channel=2
    6, 0, -6, 10, -5, 9, 7, 0, 5,
    -- layer=1 filter=238 channel=3
    4, -10, 5, -7, 6, 0, 3, -1, -6,
    -- layer=1 filter=238 channel=4
    -6, -3, 0, 3, -3, -10, -8, 1, -7,
    -- layer=1 filter=238 channel=5
    8, -8, 2, -4, -4, 5, -2, -3, -7,
    -- layer=1 filter=238 channel=6
    -7, 6, 3, -8, 2, -2, 9, 1, 9,
    -- layer=1 filter=238 channel=7
    2, 6, 6, 0, 0, 0, 5, 5, 3,
    -- layer=1 filter=238 channel=8
    1, -2, 6, 2, -9, -10, -7, -8, 0,
    -- layer=1 filter=238 channel=9
    -3, -7, -3, 5, 2, 3, 7, -11, 0,
    -- layer=1 filter=238 channel=10
    -1, 7, 1, -6, -8, -1, 2, 3, 5,
    -- layer=1 filter=238 channel=11
    -6, -12, 6, 4, 0, 4, -2, -5, 0,
    -- layer=1 filter=238 channel=12
    5, 8, 4, -7, 10, 6, 2, -2, 0,
    -- layer=1 filter=238 channel=13
    0, -2, -7, -3, -2, -4, 2, 0, -13,
    -- layer=1 filter=238 channel=14
    6, -7, 0, 6, -5, 4, -2, 6, 1,
    -- layer=1 filter=238 channel=15
    -6, 0, 9, 2, -7, 2, -6, -11, 4,
    -- layer=1 filter=238 channel=16
    6, -9, -4, -9, 9, -4, -11, -10, 1,
    -- layer=1 filter=238 channel=17
    -10, 4, -3, -2, -11, -10, 2, -8, 5,
    -- layer=1 filter=238 channel=18
    -9, 5, -1, 3, 6, 3, 0, 2, -6,
    -- layer=1 filter=238 channel=19
    -1, 11, 6, 0, -5, -1, 4, 0, -6,
    -- layer=1 filter=238 channel=20
    4, -9, -10, -13, 4, -12, -3, 7, 1,
    -- layer=1 filter=238 channel=21
    2, 9, -2, 4, 2, -5, 1, 1, 4,
    -- layer=1 filter=238 channel=22
    1, 0, 5, 1, 0, 6, 8, 8, -10,
    -- layer=1 filter=238 channel=23
    6, 7, -3, -4, -12, 10, -6, 6, 2,
    -- layer=1 filter=238 channel=24
    5, -9, 0, -2, 3, 3, 4, 0, 6,
    -- layer=1 filter=238 channel=25
    -5, -6, 1, -6, -5, 0, -10, 1, -7,
    -- layer=1 filter=238 channel=26
    3, 4, -13, -11, -2, 4, -14, 4, 7,
    -- layer=1 filter=238 channel=27
    3, 5, 8, -10, 1, -9, 4, -8, 9,
    -- layer=1 filter=238 channel=28
    -6, 8, 0, -5, -1, -7, -4, 0, 7,
    -- layer=1 filter=238 channel=29
    1, -7, -6, -4, 4, 0, -1, 1, 7,
    -- layer=1 filter=238 channel=30
    -8, 5, -5, -4, -4, -1, -10, 1, -10,
    -- layer=1 filter=238 channel=31
    0, 8, 1, 1, -6, -7, 5, -8, -5,
    -- layer=1 filter=238 channel=32
    -8, -8, -10, -5, -2, -8, 2, -6, 10,
    -- layer=1 filter=238 channel=33
    -6, 4, -1, -8, 4, 9, 5, 9, 0,
    -- layer=1 filter=238 channel=34
    1, -1, -1, -2, -4, 3, 7, -3, 5,
    -- layer=1 filter=238 channel=35
    4, -3, 0, -3, -2, -8, 8, -8, 7,
    -- layer=1 filter=238 channel=36
    -7, -5, -7, -4, 6, -9, 6, -3, -11,
    -- layer=1 filter=238 channel=37
    -11, 9, 1, 1, -8, -9, -8, 6, 0,
    -- layer=1 filter=238 channel=38
    4, 3, -3, -1, -10, -1, 8, -11, 7,
    -- layer=1 filter=238 channel=39
    -9, 2, 8, 2, -10, 0, -10, -3, -10,
    -- layer=1 filter=238 channel=40
    -6, -3, -4, -3, 7, -5, 3, 2, -10,
    -- layer=1 filter=238 channel=41
    0, 4, 2, 8, -1, 9, -2, 4, -1,
    -- layer=1 filter=238 channel=42
    2, 2, -2, 1, -5, -7, 8, -4, -2,
    -- layer=1 filter=238 channel=43
    5, 3, 2, 8, 4, 2, 3, 7, -11,
    -- layer=1 filter=238 channel=44
    0, 0, 3, 1, -4, 0, 2, -7, 2,
    -- layer=1 filter=238 channel=45
    -11, 0, -11, 8, 5, 3, 1, -3, 0,
    -- layer=1 filter=238 channel=46
    -6, 8, 0, -10, 5, 10, -7, 1, 0,
    -- layer=1 filter=238 channel=47
    8, -14, 5, 7, 2, 3, 0, -5, 6,
    -- layer=1 filter=238 channel=48
    -6, -9, -1, -2, -1, -7, -6, -7, -9,
    -- layer=1 filter=238 channel=49
    7, -1, -5, 4, -11, 0, 0, -6, 9,
    -- layer=1 filter=238 channel=50
    8, -6, 8, -1, 3, 4, -4, 6, -2,
    -- layer=1 filter=238 channel=51
    3, -6, 3, -5, -7, 3, -3, -1, 5,
    -- layer=1 filter=238 channel=52
    -10, 8, 2, -4, -10, 7, -3, 8, 0,
    -- layer=1 filter=238 channel=53
    -6, 3, 6, -9, 0, 6, 6, -5, -9,
    -- layer=1 filter=238 channel=54
    -1, 10, 8, 6, 5, 8, 6, 7, -1,
    -- layer=1 filter=238 channel=55
    4, -7, 3, -7, -10, -1, 4, 7, -8,
    -- layer=1 filter=238 channel=56
    0, 8, 7, 7, -5, -7, 0, 10, -5,
    -- layer=1 filter=238 channel=57
    -5, 1, -12, -2, 7, 0, 0, -11, -13,
    -- layer=1 filter=238 channel=58
    -5, 5, 5, 6, 1, -8, -2, 6, -8,
    -- layer=1 filter=238 channel=59
    2, 0, -9, -7, 4, -1, 5, 4, 0,
    -- layer=1 filter=238 channel=60
    -6, 1, -3, -2, 0, 10, 6, -3, 3,
    -- layer=1 filter=238 channel=61
    9, 3, 10, -5, 5, 11, -1, -5, 0,
    -- layer=1 filter=238 channel=62
    -6, 9, 2, -7, -7, -3, -3, -8, 0,
    -- layer=1 filter=238 channel=63
    5, 1, 9, -2, -13, -9, -4, -5, -3,
    -- layer=1 filter=238 channel=64
    2, -7, -7, -2, -8, -6, 3, 0, 7,
    -- layer=1 filter=238 channel=65
    -9, -7, 3, -3, 5, -4, -5, -1, -9,
    -- layer=1 filter=238 channel=66
    -13, -11, 3, 4, 1, 5, 0, -9, -8,
    -- layer=1 filter=238 channel=67
    -11, -1, -5, 0, 0, -2, -6, 0, -8,
    -- layer=1 filter=238 channel=68
    -10, -6, -4, -2, -6, 5, -7, -3, -8,
    -- layer=1 filter=238 channel=69
    2, 0, -3, -4, 1, 7, 4, -1, -11,
    -- layer=1 filter=238 channel=70
    -4, 9, -3, -3, -7, 0, 1, 10, -1,
    -- layer=1 filter=238 channel=71
    -9, -6, 0, -6, -8, -7, -8, -5, -3,
    -- layer=1 filter=238 channel=72
    -1, 10, -8, 2, -2, -5, 6, 7, 5,
    -- layer=1 filter=238 channel=73
    -3, 9, 2, 7, -4, 8, 0, 0, -9,
    -- layer=1 filter=238 channel=74
    4, 0, -6, 3, 8, 3, 7, 5, 0,
    -- layer=1 filter=238 channel=75
    -9, 9, -1, -2, 5, -7, -2, -9, 4,
    -- layer=1 filter=238 channel=76
    -9, 0, -6, 2, 1, -3, -7, -7, 6,
    -- layer=1 filter=238 channel=77
    0, -2, 3, -12, 3, 0, 8, 6, -1,
    -- layer=1 filter=238 channel=78
    1, 3, -3, -10, 1, 0, 0, -9, 7,
    -- layer=1 filter=238 channel=79
    -11, -7, 2, 0, 1, 5, -2, 0, -10,
    -- layer=1 filter=238 channel=80
    -5, -5, 9, 8, -5, 0, 9, -6, -3,
    -- layer=1 filter=238 channel=81
    -7, -8, 5, -10, 8, 4, 0, 0, -3,
    -- layer=1 filter=238 channel=82
    3, -7, -9, -2, -2, -9, -6, 2, -2,
    -- layer=1 filter=238 channel=83
    6, -7, 8, 7, -4, 0, -12, 7, -2,
    -- layer=1 filter=238 channel=84
    6, -7, -6, 8, -1, -3, 1, -1, 0,
    -- layer=1 filter=238 channel=85
    -1, 0, -8, -3, -12, -10, -5, 0, -1,
    -- layer=1 filter=238 channel=86
    4, -4, 2, -3, -9, -11, 5, -8, 1,
    -- layer=1 filter=238 channel=87
    -4, 7, -3, -10, 6, -3, 5, 1, 2,
    -- layer=1 filter=238 channel=88
    1, -2, -1, 2, -6, -7, -6, 8, 4,
    -- layer=1 filter=238 channel=89
    -1, -5, 3, 3, 4, 5, -8, -1, 0,
    -- layer=1 filter=238 channel=90
    -1, 2, -9, -2, 1, -2, -10, 8, 4,
    -- layer=1 filter=238 channel=91
    1, -8, -11, -2, -5, -4, -2, 7, -3,
    -- layer=1 filter=238 channel=92
    2, -5, -6, 7, 1, 0, 5, 2, 2,
    -- layer=1 filter=238 channel=93
    -10, -10, -12, 1, 7, 0, -11, -8, -6,
    -- layer=1 filter=238 channel=94
    -8, -8, -10, -2, 6, 0, -8, 1, 0,
    -- layer=1 filter=238 channel=95
    -4, 2, -6, 0, -14, -9, -1, -4, -1,
    -- layer=1 filter=238 channel=96
    -11, -3, -6, -5, 3, -9, -7, 8, 0,
    -- layer=1 filter=238 channel=97
    -11, -11, -12, -8, -8, -6, 3, 8, 1,
    -- layer=1 filter=238 channel=98
    -14, 3, -6, -6, 3, -4, -11, 3, 2,
    -- layer=1 filter=238 channel=99
    2, -6, 8, -1, -9, -9, -11, 5, 7,
    -- layer=1 filter=238 channel=100
    -8, -4, -1, 5, 1, -5, -8, -7, -2,
    -- layer=1 filter=238 channel=101
    -9, 2, -13, -9, -6, -3, -12, 4, -3,
    -- layer=1 filter=238 channel=102
    -6, -10, 7, -12, -6, 3, -4, 5, -10,
    -- layer=1 filter=238 channel=103
    -5, 4, 0, -7, -11, 9, -9, -6, 10,
    -- layer=1 filter=238 channel=104
    0, 8, -4, 6, -2, 3, -7, -4, -5,
    -- layer=1 filter=238 channel=105
    -16, 3, -12, 0, -8, 6, 4, 4, -6,
    -- layer=1 filter=238 channel=106
    3, 2, 8, 8, -4, -1, -12, 0, -3,
    -- layer=1 filter=238 channel=107
    0, -7, 6, 3, -5, 2, -2, 0, 5,
    -- layer=1 filter=238 channel=108
    7, -10, -12, -11, -7, -12, 6, -1, -12,
    -- layer=1 filter=238 channel=109
    1, 6, -5, 6, -1, -2, 2, -2, 3,
    -- layer=1 filter=238 channel=110
    -5, 8, 0, -2, -7, -1, 8, -4, 1,
    -- layer=1 filter=238 channel=111
    -8, 5, 2, -4, -3, 9, -15, 3, -2,
    -- layer=1 filter=238 channel=112
    4, -9, 6, -6, 5, -3, -9, -8, -5,
    -- layer=1 filter=238 channel=113
    0, -4, -9, -2, -3, 4, -9, 9, -6,
    -- layer=1 filter=238 channel=114
    -6, 0, 6, -4, -9, -3, -5, 0, -5,
    -- layer=1 filter=238 channel=115
    3, 5, 3, -7, -6, -12, -11, -7, -5,
    -- layer=1 filter=238 channel=116
    8, -2, -2, 0, -1, 0, 3, 4, 1,
    -- layer=1 filter=238 channel=117
    -4, -11, 7, -5, 7, 4, -9, -9, 1,
    -- layer=1 filter=238 channel=118
    -10, -11, -4, 0, 0, 6, -10, -5, -3,
    -- layer=1 filter=238 channel=119
    -4, -12, -3, 3, 0, -9, -6, -10, 9,
    -- layer=1 filter=238 channel=120
    -10, -5, 2, -11, -9, -7, -8, -6, 8,
    -- layer=1 filter=238 channel=121
    -9, -3, 0, 2, 1, 3, 0, -6, 3,
    -- layer=1 filter=238 channel=122
    5, 4, 7, 7, 7, -5, -10, -8, -9,
    -- layer=1 filter=238 channel=123
    2, 3, -11, 5, -3, -2, -9, -10, 1,
    -- layer=1 filter=238 channel=124
    0, 10, 7, -4, 8, -4, 0, 0, 0,
    -- layer=1 filter=238 channel=125
    -3, 6, -5, -1, -2, -10, 5, 1, 6,
    -- layer=1 filter=238 channel=126
    -3, 5, -11, 5, -8, -6, 0, -8, 1,
    -- layer=1 filter=238 channel=127
    -3, -8, 7, -6, 4, 7, 3, 2, 0,
    -- layer=1 filter=239 channel=0
    -9, -27, -10, -8, -16, -61, -51, -35, -37,
    -- layer=1 filter=239 channel=1
    -95, -42, -12, -1, 1, 33, 18, 2, 30,
    -- layer=1 filter=239 channel=2
    69, 48, 38, 80, 86, 88, 37, 34, 27,
    -- layer=1 filter=239 channel=3
    0, 2, 5, -11, -6, -5, 10, -7, 0,
    -- layer=1 filter=239 channel=4
    5, 5, 1, -4, -5, 5, 3, 0, -4,
    -- layer=1 filter=239 channel=5
    -53, -82, -37, 14, 41, 42, 17, 23, 65,
    -- layer=1 filter=239 channel=6
    -30, -9, -45, 20, 12, 17, -33, -7, -5,
    -- layer=1 filter=239 channel=7
    -6, 13, -12, -33, -50, -54, -20, 37, -65,
    -- layer=1 filter=239 channel=8
    -91, -78, -39, 9, 24, 27, 18, 22, 55,
    -- layer=1 filter=239 channel=9
    40, 34, 49, 68, 9, 80, -9, 25, 2,
    -- layer=1 filter=239 channel=10
    -19, 15, 5, -25, -21, -51, -14, 65, -35,
    -- layer=1 filter=239 channel=11
    0, -10, 16, -21, -53, -68, -44, -68, -57,
    -- layer=1 filter=239 channel=12
    46, 116, 68, -22, 9, 32, -8, 10, 33,
    -- layer=1 filter=239 channel=13
    -31, -27, -31, 8, 13, 15, 22, -2, 38,
    -- layer=1 filter=239 channel=14
    18, 95, 44, -10, 7, 30, -25, 6, -39,
    -- layer=1 filter=239 channel=15
    -19, -77, 7, 27, 29, 44, 36, 12, 81,
    -- layer=1 filter=239 channel=16
    -71, -61, -68, 12, 51, 26, 42, 42, 71,
    -- layer=1 filter=239 channel=17
    -32, -48, -35, -41, -15, -12, -20, -45, -25,
    -- layer=1 filter=239 channel=18
    21, 52, 53, -28, -12, 14, -15, -18, -4,
    -- layer=1 filter=239 channel=19
    -9, -15, -31, 2, 19, 18, 27, 45, 52,
    -- layer=1 filter=239 channel=20
    -44, -72, -37, -9, 4, 2, 22, 1, 26,
    -- layer=1 filter=239 channel=21
    -56, -44, -52, -20, -26, -18, 26, 33, 0,
    -- layer=1 filter=239 channel=22
    -67, -64, -33, -16, -5, 18, 20, 9, 41,
    -- layer=1 filter=239 channel=23
    11, -8, -49, 1, -23, -20, 13, -8, -4,
    -- layer=1 filter=239 channel=24
    -16, -49, -36, 15, -5, -12, 21, 29, 42,
    -- layer=1 filter=239 channel=25
    -13, -27, -19, 6, 18, -30, 10, 52, 9,
    -- layer=1 filter=239 channel=26
    17, -45, 0, 22, -17, 7, 17, -32, 21,
    -- layer=1 filter=239 channel=27
    -10, -8, -15, 15, 19, 4, -13, -20, -5,
    -- layer=1 filter=239 channel=28
    -43, 13, -29, -39, -16, -67, -27, 36, -39,
    -- layer=1 filter=239 channel=29
    23, 6, -13, -32, 15, -15, -18, -27, 3,
    -- layer=1 filter=239 channel=30
    -3, 29, 35, -12, -26, 33, -21, -55, -26,
    -- layer=1 filter=239 channel=31
    14, 69, 18, 12, 23, 59, -1, 2, 30,
    -- layer=1 filter=239 channel=32
    33, -12, 13, 34, -17, -36, 30, -2, -15,
    -- layer=1 filter=239 channel=33
    -26, -8, -9, 10, -2, 16, -21, -29, -31,
    -- layer=1 filter=239 channel=34
    -41, -11, -6, 19, 2, 5, -30, -18, -11,
    -- layer=1 filter=239 channel=35
    0, -9, 11, -7, -6, 9, 3, -11, 0,
    -- layer=1 filter=239 channel=36
    -7, -24, -3, -33, -74, -76, -51, -75, -66,
    -- layer=1 filter=239 channel=37
    -53, -60, -75, 16, 43, 27, 25, 51, 70,
    -- layer=1 filter=239 channel=38
    -38, -30, -33, -15, -1, 12, 9, 24, 16,
    -- layer=1 filter=239 channel=39
    -52, -44, -51, -4, -19, 17, -41, -27, -11,
    -- layer=1 filter=239 channel=40
    1, 56, 48, 19, 35, 46, -46, -21, 18,
    -- layer=1 filter=239 channel=41
    27, -8, 20, 48, -40, 19, 39, 50, -19,
    -- layer=1 filter=239 channel=42
    57, 49, 30, 73, 90, 84, 59, 44, 44,
    -- layer=1 filter=239 channel=43
    -70, -43, -34, 28, 35, 15, 18, 33, 46,
    -- layer=1 filter=239 channel=44
    12, -49, 6, 19, -71, -46, 17, -34, 0,
    -- layer=1 filter=239 channel=45
    -49, -83, -45, -16, -7, -4, 32, 15, 81,
    -- layer=1 filter=239 channel=46
    21, 19, -21, 55, 64, 74, 36, 37, 139,
    -- layer=1 filter=239 channel=47
    7, -30, 2, 20, 28, -9, 22, 43, 21,
    -- layer=1 filter=239 channel=48
    -39, -52, -9, -31, -33, -68, -26, 22, -38,
    -- layer=1 filter=239 channel=49
    13, -2, -24, 34, 20, 14, 10, 38, 6,
    -- layer=1 filter=239 channel=50
    -14, -16, 5, -8, -24, 5, -11, -8, -7,
    -- layer=1 filter=239 channel=51
    -24, -3, 14, -16, -4, -24, -25, 15, -34,
    -- layer=1 filter=239 channel=52
    2, -17, -2, 31, -7, 38, 20, 15, 6,
    -- layer=1 filter=239 channel=53
    -4, -2, -12, 1, 18, -1, -9, -1, -3,
    -- layer=1 filter=239 channel=54
    -21, -41, -55, 26, 32, -19, 38, 79, 28,
    -- layer=1 filter=239 channel=55
    -24, -34, -11, 5, -28, -25, -44, -26, -27,
    -- layer=1 filter=239 channel=56
    4, 2, 2, 9, -6, 9, -3, 7, 3,
    -- layer=1 filter=239 channel=57
    -11, 8, 8, -22, -18, -23, -27, 36, -35,
    -- layer=1 filter=239 channel=58
    -3, -21, -12, 0, -37, -21, 12, 78, -38,
    -- layer=1 filter=239 channel=59
    -4, 2, 1, -1, 0, -7, -7, -11, 0,
    -- layer=1 filter=239 channel=60
    -18, 0, 3, 0, 5, 3, -4, 5, 10,
    -- layer=1 filter=239 channel=61
    1, -12, 3, -9, -2, 10, 5, -4, -7,
    -- layer=1 filter=239 channel=62
    -63, -67, -64, 14, 34, 4, 26, 37, 72,
    -- layer=1 filter=239 channel=63
    9, 15, 27, -27, -59, -46, -36, -61, -66,
    -- layer=1 filter=239 channel=64
    -32, -38, -25, -4, -36, -31, 2, 17, -15,
    -- layer=1 filter=239 channel=65
    -42, -35, -55, -38, -37, -51, -16, -18, -34,
    -- layer=1 filter=239 channel=66
    0, -21, -36, -28, -59, -63, -66, -45, -40,
    -- layer=1 filter=239 channel=67
    23, 20, 18, 16, -1, 16, 19, -33, 15,
    -- layer=1 filter=239 channel=68
    11, -38, -9, 1, -60, -44, 1, -26, -3,
    -- layer=1 filter=239 channel=69
    -11, -66, -27, 15, 34, 30, 43, 9, 73,
    -- layer=1 filter=239 channel=70
    -52, -13, -42, -10, -21, 27, 16, 10, 38,
    -- layer=1 filter=239 channel=71
    -29, -56, -62, -29, -9, -20, 7, 11, 6,
    -- layer=1 filter=239 channel=72
    26, 26, -3, 2, 6, 41, 30, -3, 8,
    -- layer=1 filter=239 channel=73
    -1, 11, -10, 18, 0, -2, -4, 0, 0,
    -- layer=1 filter=239 channel=74
    12, 13, 1, 18, 10, 7, -10, -3, 3,
    -- layer=1 filter=239 channel=75
    33, 85, 14, -19, 30, 63, -19, -22, -7,
    -- layer=1 filter=239 channel=76
    -2, -9, 6, 32, -12, -22, 5, -31, -6,
    -- layer=1 filter=239 channel=77
    -46, -36, -55, -43, -59, -82, -28, 31, -4,
    -- layer=1 filter=239 channel=78
    -3, -10, -11, 19, -22, -20, 5, 12, -39,
    -- layer=1 filter=239 channel=79
    -79, -86, -59, 2, 25, 12, 27, 30, 52,
    -- layer=1 filter=239 channel=80
    18, 21, 10, 37, -10, 6, -1, 0, 5,
    -- layer=1 filter=239 channel=81
    -56, -66, -76, -13, -28, -43, -4, 21, 23,
    -- layer=1 filter=239 channel=82
    -50, -64, -56, -47, -30, -53, -1, 14, -7,
    -- layer=1 filter=239 channel=83
    -45, -70, -7, -20, -44, 13, -19, -37, 35,
    -- layer=1 filter=239 channel=84
    24, 43, 60, 34, 4, 3, -12, -53, -34,
    -- layer=1 filter=239 channel=85
    24, -18, 5, 34, 7, 5, 49, 57, -7,
    -- layer=1 filter=239 channel=86
    -36, -34, -51, -60, -55, -47, -62, -54, -33,
    -- layer=1 filter=239 channel=87
    19, 20, -15, 14, 11, 43, 56, 66, 53,
    -- layer=1 filter=239 channel=88
    -7, -23, -26, 0, -1, -22, -18, 6, -15,
    -- layer=1 filter=239 channel=89
    -24, -28, -43, -12, -39, -31, -18, -19, -24,
    -- layer=1 filter=239 channel=90
    -4, -64, -5, 12, -74, -25, 23, -40, 8,
    -- layer=1 filter=239 channel=91
    -23, -21, -10, -22, -10, -12, -36, -8, -25,
    -- layer=1 filter=239 channel=92
    -4, -34, 24, 36, -22, -50, 15, -1, 31,
    -- layer=1 filter=239 channel=93
    -61, -78, -60, -68, -53, -76, 0, -8, -16,
    -- layer=1 filter=239 channel=94
    -38, -12, -12, -49, -29, -48, -53, -22, -20,
    -- layer=1 filter=239 channel=95
    22, 40, 37, 6, -12, 9, -12, -62, -40,
    -- layer=1 filter=239 channel=96
    12, 9, -9, 28, 11, -4, -6, -33, -16,
    -- layer=1 filter=239 channel=97
    -28, -23, -32, -57, -71, -70, -27, -23, -13,
    -- layer=1 filter=239 channel=98
    -112, -74, -71, -10, 36, -10, 12, 44, 43,
    -- layer=1 filter=239 channel=99
    -64, 21, 0, -46, -28, -62, -66, 23, -39,
    -- layer=1 filter=239 channel=100
    0, -8, -10, -25, -20, -28, 5, -46, -33,
    -- layer=1 filter=239 channel=101
    -53, -21, -15, -15, -29, -34, -11, -6, -26,
    -- layer=1 filter=239 channel=102
    -14, -25, -19, 3, -20, -31, -42, -52, -21,
    -- layer=1 filter=239 channel=103
    5, -2, 14, -44, -78, -36, -18, -55, -8,
    -- layer=1 filter=239 channel=104
    17, 23, 0, 14, -11, -10, 1, 8, -5,
    -- layer=1 filter=239 channel=105
    -25, -13, 1, -75, -77, -110, -48, -15, -65,
    -- layer=1 filter=239 channel=106
    3, -20, -2, 4, -15, -29, 17, -4, 6,
    -- layer=1 filter=239 channel=107
    -9, -4, -11, -9, -7, -5, 15, 14, 17,
    -- layer=1 filter=239 channel=108
    22, -57, 19, 40, -58, -8, 36, -16, 21,
    -- layer=1 filter=239 channel=109
    5, -6, 4, -8, 1, 1, -11, -10, 1,
    -- layer=1 filter=239 channel=110
    2, 2, 2, -6, -23, -20, -20, 7, -10,
    -- layer=1 filter=239 channel=111
    1, 29, 54, -6, -20, -17, -42, -59, -63,
    -- layer=1 filter=239 channel=112
    10, 45, 57, 11, 4, -29, -11, -26, -28,
    -- layer=1 filter=239 channel=113
    7, 1, -1, 45, 94, 38, 50, 47, 51,
    -- layer=1 filter=239 channel=114
    -5, -36, -20, 42, 59, 63, 6, 1, 82,
    -- layer=1 filter=239 channel=115
    -55, -9, -23, -65, -40, -61, -56, -1, -35,
    -- layer=1 filter=239 channel=116
    8, -6, 7, 0, -9, 0, -3, 8, -6,
    -- layer=1 filter=239 channel=117
    5, 73, 87, -8, -11, -14, -7, -67, -51,
    -- layer=1 filter=239 channel=118
    13, 22, 30, 19, 8, 17, -26, -77, -30,
    -- layer=1 filter=239 channel=119
    16, -70, 8, 25, -68, -51, 23, -39, -13,
    -- layer=1 filter=239 channel=120
    -39, -71, -45, -16, -16, -37, 8, 36, -6,
    -- layer=1 filter=239 channel=121
    15, 41, -6, -10, -6, 50, -33, -18, -37,
    -- layer=1 filter=239 channel=122
    -5, -7, -10, 7, 8, 3, 4, 1, 0,
    -- layer=1 filter=239 channel=123
    8, 31, -14, -26, -5, 14, -20, -31, -41,
    -- layer=1 filter=239 channel=124
    -4, 1, 2, 4, 20, 6, 2, 7, -2,
    -- layer=1 filter=239 channel=125
    -53, -18, -4, -8, -8, -14, 11, 50, 28,
    -- layer=1 filter=239 channel=126
    -92, -77, -59, -29, -12, -18, -3, 25, 26,
    -- layer=1 filter=239 channel=127
    26, 40, 36, 11, 16, 22, -20, -58, -16,
    -- layer=1 filter=240 channel=0
    13, 15, -3, -59, -53, -40, -48, -55, -30,
    -- layer=1 filter=240 channel=1
    -67, -22, -71, -2, -17, -3, -7, -54, -88,
    -- layer=1 filter=240 channel=2
    -76, -54, -3, -32, -24, 8, -10, -10, -4,
    -- layer=1 filter=240 channel=3
    8, 10, -8, 0, -5, 8, 6, -9, 8,
    -- layer=1 filter=240 channel=4
    -1, 2, -3, 21, 46, 10, -1, -4, -10,
    -- layer=1 filter=240 channel=5
    -43, -24, -104, -42, -7, 1, -20, -51, -71,
    -- layer=1 filter=240 channel=6
    -11, 13, 32, 14, 19, 24, -36, -13, -12,
    -- layer=1 filter=240 channel=7
    10, -71, -38, 32, -34, -43, -52, 29, -44,
    -- layer=1 filter=240 channel=8
    -49, -21, -64, -31, -21, -3, -11, -52, -90,
    -- layer=1 filter=240 channel=9
    -31, -49, 43, 24, 79, 26, -77, -59, -8,
    -- layer=1 filter=240 channel=10
    27, -59, -56, 17, 7, -19, -47, 15, -39,
    -- layer=1 filter=240 channel=11
    15, -2, 22, -7, -4, -23, -3, -14, 14,
    -- layer=1 filter=240 channel=12
    -22, 5, 49, 60, 11, 2, -74, -30, -92,
    -- layer=1 filter=240 channel=13
    15, 21, 28, -19, -25, 5, 12, 6, 14,
    -- layer=1 filter=240 channel=14
    -12, -48, -39, 53, -39, -1, -47, 0, -44,
    -- layer=1 filter=240 channel=15
    20, -13, -39, -51, -43, -39, 32, -1, -35,
    -- layer=1 filter=240 channel=16
    -61, -59, -94, -20, -28, -6, -21, -41, -46,
    -- layer=1 filter=240 channel=17
    18, 13, 3, -69, -51, -47, -35, -21, -30,
    -- layer=1 filter=240 channel=18
    31, 31, 49, 36, 21, -10, -75, -24, -36,
    -- layer=1 filter=240 channel=19
    -97, -117, 3, 23, 72, 26, -86, -29, -13,
    -- layer=1 filter=240 channel=20
    -3, -5, -32, -15, -32, -27, -13, -6, -17,
    -- layer=1 filter=240 channel=21
    -45, -27, -11, -17, -44, -8, -21, -2, -22,
    -- layer=1 filter=240 channel=22
    19, 17, 12, -40, -69, -30, 29, 17, 1,
    -- layer=1 filter=240 channel=23
    -15, -6, 4, -14, 10, -29, 10, 18, -8,
    -- layer=1 filter=240 channel=24
    -36, -55, 5, -41, -6, 17, 0, -36, 2,
    -- layer=1 filter=240 channel=25
    -3, -71, -20, -18, 12, -16, -50, -16, -58,
    -- layer=1 filter=240 channel=26
    1, -5, 38, -2, -1, 14, 27, -4, 7,
    -- layer=1 filter=240 channel=27
    -14, 8, 4, -44, -76, -55, -41, -15, -3,
    -- layer=1 filter=240 channel=28
    4, -63, -8, 23, -55, -30, -23, 11, -42,
    -- layer=1 filter=240 channel=29
    5, -12, 0, -21, -26, -16, -47, -30, -14,
    -- layer=1 filter=240 channel=30
    24, 4, 36, 54, 52, 5, -108, -61, -62,
    -- layer=1 filter=240 channel=31
    1, 7, 17, 46, 20, 17, -71, -49, -63,
    -- layer=1 filter=240 channel=32
    -10, 21, 64, 14, 17, 7, 24, -12, -22,
    -- layer=1 filter=240 channel=33
    12, 7, -8, -16, -22, -12, -15, 9, 19,
    -- layer=1 filter=240 channel=34
    5, -8, -19, 5, -33, -8, -36, -28, 19,
    -- layer=1 filter=240 channel=35
    -1, 2, -16, -12, 3, -18, -12, -13, -11,
    -- layer=1 filter=240 channel=36
    0, 4, -3, -1, -7, -13, -20, -30, 10,
    -- layer=1 filter=240 channel=37
    -34, -60, -119, -18, 11, 17, -51, -48, -38,
    -- layer=1 filter=240 channel=38
    1, -10, -2, 0, 4, -4, -26, -6, 11,
    -- layer=1 filter=240 channel=39
    -19, -26, -41, -27, -19, -23, -22, -53, -10,
    -- layer=1 filter=240 channel=40
    35, 26, 40, 43, 8, -10, -36, -20, -25,
    -- layer=1 filter=240 channel=41
    -47, -3, 43, 6, 60, 21, 10, -19, 17,
    -- layer=1 filter=240 channel=42
    -66, -42, -24, 2, -14, 11, -4, 8, 13,
    -- layer=1 filter=240 channel=43
    -59, -55, -67, -28, 1, -19, -26, -36, -76,
    -- layer=1 filter=240 channel=44
    -33, 4, 31, -33, -22, 10, 20, -13, -23,
    -- layer=1 filter=240 channel=45
    -27, -16, -43, -13, -47, -33, 12, -24, -34,
    -- layer=1 filter=240 channel=46
    -105, -123, -57, 25, 38, 37, -59, -20, -24,
    -- layer=1 filter=240 channel=47
    -18, -1, 7, -38, 0, -30, 11, -29, 19,
    -- layer=1 filter=240 channel=48
    20, -2, 6, -45, -23, -29, -44, -30, -10,
    -- layer=1 filter=240 channel=49
    -10, -23, -22, -37, -8, -20, -36, -9, 4,
    -- layer=1 filter=240 channel=50
    28, 13, -4, 1, 53, 16, -9, -3, -7,
    -- layer=1 filter=240 channel=51
    12, -8, -10, 13, -11, -19, -49, -11, -35,
    -- layer=1 filter=240 channel=52
    6, -4, -6, -20, -9, 10, 8, 4, -3,
    -- layer=1 filter=240 channel=53
    9, -4, 0, 5, 10, -1, -1, 11, 1,
    -- layer=1 filter=240 channel=54
    20, -51, -25, -54, 24, -3, -66, -2, -45,
    -- layer=1 filter=240 channel=55
    -51, -39, -31, -26, 0, 7, 28, -1, 5,
    -- layer=1 filter=240 channel=56
    7, -6, 0, -3, -8, -5, -4, -9, 1,
    -- layer=1 filter=240 channel=57
    15, -44, -44, 0, 7, -22, -35, 13, -25,
    -- layer=1 filter=240 channel=58
    7, -51, -18, -40, 64, -51, -54, -5, -31,
    -- layer=1 filter=240 channel=59
    -9, -12, -6, 6, 2, -3, -9, -4, -8,
    -- layer=1 filter=240 channel=60
    0, -1, 13, -1, 2, -19, -4, 0, 11,
    -- layer=1 filter=240 channel=61
    -9, -3, 5, -7, -6, 3, 4, 4, 1,
    -- layer=1 filter=240 channel=62
    -57, -54, -90, -42, -16, 2, -36, -44, -63,
    -- layer=1 filter=240 channel=63
    0, 20, 11, 20, -13, -27, -3, -8, 6,
    -- layer=1 filter=240 channel=64
    -13, 27, 6, -15, -39, -15, -13, 1, 3,
    -- layer=1 filter=240 channel=65
    -12, 3, -9, -2, -21, -3, -35, -14, -7,
    -- layer=1 filter=240 channel=66
    -4, -7, -34, -34, -38, -41, -26, -28, -28,
    -- layer=1 filter=240 channel=67
    -17, -21, -11, -72, -27, -33, -55, -31, -11,
    -- layer=1 filter=240 channel=68
    -9, 22, 52, -11, -1, 10, 15, -14, -10,
    -- layer=1 filter=240 channel=69
    -47, -46, -71, -34, -32, -11, 10, -23, -47,
    -- layer=1 filter=240 channel=70
    16, 12, -13, 0, 14, 9, -53, -17, -22,
    -- layer=1 filter=240 channel=71
    -26, 8, -4, 1, -17, -8, -20, -1, -17,
    -- layer=1 filter=240 channel=72
    -54, -37, 54, 65, 57, 25, -94, -62, -38,
    -- layer=1 filter=240 channel=73
    -13, 2, 2, -8, -5, -7, -3, 6, -7,
    -- layer=1 filter=240 channel=74
    17, 58, 54, 35, 28, 21, -57, -83, -27,
    -- layer=1 filter=240 channel=75
    -25, 8, 34, 51, 24, 0, -74, -32, -41,
    -- layer=1 filter=240 channel=76
    8, 17, 51, -8, -6, -22, -28, -44, -28,
    -- layer=1 filter=240 channel=77
    -20, -20, -4, 2, -1, 14, -46, -51, -33,
    -- layer=1 filter=240 channel=78
    23, -29, -43, 21, 10, -4, -24, -6, -23,
    -- layer=1 filter=240 channel=79
    -39, -51, -93, -26, -19, -21, -19, -32, -51,
    -- layer=1 filter=240 channel=80
    1, -20, -16, -25, -20, -34, -14, -4, -32,
    -- layer=1 filter=240 channel=81
    -56, -53, -33, -13, -16, 6, -31, -40, -17,
    -- layer=1 filter=240 channel=82
    -2, 15, 5, -46, -45, -15, -33, -8, -19,
    -- layer=1 filter=240 channel=83
    -5, -37, -39, -15, -23, -14, -2, -20, -91,
    -- layer=1 filter=240 channel=84
    42, 38, 73, 21, 18, -18, -37, -30, -22,
    -- layer=1 filter=240 channel=85
    0, -41, 18, -31, 45, -18, -49, 10, -28,
    -- layer=1 filter=240 channel=86
    -21, -15, -46, 9, -7, -13, -22, -25, -30,
    -- layer=1 filter=240 channel=87
    -72, -99, 21, 31, 78, 30, -70, -35, 31,
    -- layer=1 filter=240 channel=88
    -25, -31, -21, -40, -10, 2, -48, 0, -19,
    -- layer=1 filter=240 channel=89
    -4, 37, 40, -14, -40, 9, -18, -19, -6,
    -- layer=1 filter=240 channel=90
    -19, -22, 16, -19, -9, 32, 27, -27, -34,
    -- layer=1 filter=240 channel=91
    39, 23, 10, 1, -3, -13, -32, -15, -15,
    -- layer=1 filter=240 channel=92
    -7, 21, -13, -36, 14, -3, 26, 8, -25,
    -- layer=1 filter=240 channel=93
    -12, -7, -31, -51, -51, -30, -28, -29, -36,
    -- layer=1 filter=240 channel=94
    36, 13, 2, -9, -14, -29, -29, -35, -13,
    -- layer=1 filter=240 channel=95
    22, 34, 37, 43, 35, 10, -63, -62, -40,
    -- layer=1 filter=240 channel=96
    2, -2, 1, -39, 1, -14, -10, -21, -31,
    -- layer=1 filter=240 channel=97
    -5, 5, -17, -65, -87, -45, -47, -46, -52,
    -- layer=1 filter=240 channel=98
    -32, -65, -71, -29, -17, -8, -20, -22, -62,
    -- layer=1 filter=240 channel=99
    36, -35, -51, -22, -42, 1, 7, -27, 10,
    -- layer=1 filter=240 channel=100
    -10, 25, 42, 40, 18, 0, -10, -13, 8,
    -- layer=1 filter=240 channel=101
    27, 36, 3, -17, -28, -19, -22, -16, -24,
    -- layer=1 filter=240 channel=102
    49, 51, 32, -12, -27, -10, -65, -41, -44,
    -- layer=1 filter=240 channel=103
    13, 19, 55, 14, 14, -13, -20, -16, 17,
    -- layer=1 filter=240 channel=104
    4, -9, 27, -9, 55, -13, -5, -17, -1,
    -- layer=1 filter=240 channel=105
    22, 5, -11, -38, -35, -44, -45, -18, -35,
    -- layer=1 filter=240 channel=106
    31, 29, 32, -22, -5, -2, 18, -30, -13,
    -- layer=1 filter=240 channel=107
    4, 0, -5, -2, -9, -5, 0, 8, 5,
    -- layer=1 filter=240 channel=108
    -30, -27, 32, -42, -4, 12, 38, 2, -6,
    -- layer=1 filter=240 channel=109
    -3, 8, -9, 6, -6, -9, -2, -6, 4,
    -- layer=1 filter=240 channel=110
    18, 33, 3, 3, -6, -11, 10, -7, -14,
    -- layer=1 filter=240 channel=111
    53, 40, 46, 26, 19, -13, -86, -61, -51,
    -- layer=1 filter=240 channel=112
    43, 63, 37, -2, 0, -17, 23, 22, 2,
    -- layer=1 filter=240 channel=113
    16, 7, -6, -17, -35, 8, -15, -6, 7,
    -- layer=1 filter=240 channel=114
    -27, 1, -89, -36, -23, -9, 0, -49, -65,
    -- layer=1 filter=240 channel=115
    28, -11, -43, 17, 2, -36, -33, 16, -33,
    -- layer=1 filter=240 channel=116
    0, 7, -2, -8, 0, -6, -8, -4, 9,
    -- layer=1 filter=240 channel=117
    74, 61, 19, -8, 21, -28, 16, 28, 9,
    -- layer=1 filter=240 channel=118
    31, 35, 42, 42, 36, 7, -66, -84, -45,
    -- layer=1 filter=240 channel=119
    -28, -4, 55, -6, 2, 19, 16, -26, 0,
    -- layer=1 filter=240 channel=120
    -28, -52, -30, -40, -16, -24, -44, -10, -45,
    -- layer=1 filter=240 channel=121
    -43, -67, -4, 58, 65, 17, -51, -3, 10,
    -- layer=1 filter=240 channel=122
    0, 0, -10, -9, -4, 0, 6, 0, -6,
    -- layer=1 filter=240 channel=123
    -35, -35, -5, 38, 33, -3, -20, -4, -2,
    -- layer=1 filter=240 channel=124
    8, 1, 8, -2, -8, -1, 3, 0, -1,
    -- layer=1 filter=240 channel=125
    27, -5, -5, -29, -5, -3, -15, -40, -11,
    -- layer=1 filter=240 channel=126
    -40, -61, -44, -20, -7, 3, 4, -20, -59,
    -- layer=1 filter=240 channel=127
    27, 32, 45, 56, 41, 14, -92, -60, -49,
    -- layer=1 filter=241 channel=0
    2, 4, -1, 0, -9, 0, -7, 1, -8,
    -- layer=1 filter=241 channel=1
    2, -1, -2, -6, -3, 3, 8, 1, 0,
    -- layer=1 filter=241 channel=2
    3, 11, -7, -7, -2, -8, 6, -8, 0,
    -- layer=1 filter=241 channel=3
    -1, 10, 5, 7, -5, -3, -6, 0, 1,
    -- layer=1 filter=241 channel=4
    -2, 3, 1, -1, 5, 8, -11, 0, 3,
    -- layer=1 filter=241 channel=5
    -4, -12, 5, 6, 5, 6, 3, 2, -2,
    -- layer=1 filter=241 channel=6
    1, -7, -10, 0, 1, -8, -11, 0, 10,
    -- layer=1 filter=241 channel=7
    -3, 4, -3, -3, -6, -8, 5, -4, 1,
    -- layer=1 filter=241 channel=8
    6, 4, -4, 0, 0, -10, -7, 2, -2,
    -- layer=1 filter=241 channel=9
    -7, -8, -4, 2, -6, 0, -10, -11, 0,
    -- layer=1 filter=241 channel=10
    7, 6, 5, -11, -12, 10, 9, -2, -4,
    -- layer=1 filter=241 channel=11
    -4, 7, -2, 0, 3, -4, -4, -8, -2,
    -- layer=1 filter=241 channel=12
    7, 7, 9, 0, 0, -2, 9, 9, 7,
    -- layer=1 filter=241 channel=13
    -7, 9, -7, 4, 5, 1, -6, 2, -10,
    -- layer=1 filter=241 channel=14
    4, 5, -7, -9, -5, -1, 6, 0, -6,
    -- layer=1 filter=241 channel=15
    -2, 0, -7, 3, -3, -6, -3, 4, 3,
    -- layer=1 filter=241 channel=16
    4, 5, -8, 0, -7, 0, -1, 3, 0,
    -- layer=1 filter=241 channel=17
    5, -3, -3, 8, 7, 0, 1, -1, -2,
    -- layer=1 filter=241 channel=18
    -7, 2, -12, -6, -10, 0, 1, -6, -10,
    -- layer=1 filter=241 channel=19
    -5, -10, -11, -12, 4, 6, 5, 5, 0,
    -- layer=1 filter=241 channel=20
    -8, 0, 2, 2, -3, -5, -5, -10, 8,
    -- layer=1 filter=241 channel=21
    -7, -3, 8, 4, 3, 2, 4, -12, -3,
    -- layer=1 filter=241 channel=22
    -7, 0, -2, 8, 6, 4, -10, -12, -9,
    -- layer=1 filter=241 channel=23
    2, 2, -4, -8, -2, 3, -8, -3, 7,
    -- layer=1 filter=241 channel=24
    9, -11, 3, 0, -8, 0, -1, -11, -3,
    -- layer=1 filter=241 channel=25
    4, -5, 6, 4, 2, 1, 0, 8, -1,
    -- layer=1 filter=241 channel=26
    -4, 9, 4, 9, -8, 7, 8, 4, 0,
    -- layer=1 filter=241 channel=27
    -7, -10, -3, -3, 4, 1, -9, -5, 0,
    -- layer=1 filter=241 channel=28
    4, -12, -3, 1, -12, -1, -6, 7, -6,
    -- layer=1 filter=241 channel=29
    -8, -12, -6, -4, -6, 4, -1, 1, 4,
    -- layer=1 filter=241 channel=30
    7, -1, 6, 9, -11, -3, 1, 2, 2,
    -- layer=1 filter=241 channel=31
    -7, -9, -9, -3, 0, -3, -6, 6, 1,
    -- layer=1 filter=241 channel=32
    2, 2, -1, -1, -5, 3, -4, -5, 5,
    -- layer=1 filter=241 channel=33
    -9, 6, 3, 4, 5, 5, -4, -2, -1,
    -- layer=1 filter=241 channel=34
    -9, 0, 4, -2, -3, -12, -3, 8, -1,
    -- layer=1 filter=241 channel=35
    -4, -5, -5, 7, -6, -2, 9, -1, 4,
    -- layer=1 filter=241 channel=36
    -8, 5, 5, -2, 2, 2, 7, -4, -6,
    -- layer=1 filter=241 channel=37
    5, -5, 3, 7, 6, 7, 7, 9, -3,
    -- layer=1 filter=241 channel=38
    5, -6, 0, -1, -7, -5, 0, 0, -8,
    -- layer=1 filter=241 channel=39
    -5, 3, -12, -10, -5, -3, -8, 0, -2,
    -- layer=1 filter=241 channel=40
    5, 1, 4, -1, -5, -8, -4, -3, -9,
    -- layer=1 filter=241 channel=41
    6, 4, -4, 0, -10, -11, 1, -6, -4,
    -- layer=1 filter=241 channel=42
    -8, -2, -8, 0, -6, -7, 1, 0, 8,
    -- layer=1 filter=241 channel=43
    -10, -8, -5, -2, -8, -12, 8, -9, 2,
    -- layer=1 filter=241 channel=44
    -8, 0, -5, -4, -4, 0, 3, 0, -4,
    -- layer=1 filter=241 channel=45
    1, 6, 8, 8, 0, 0, -5, -11, -9,
    -- layer=1 filter=241 channel=46
    -4, 1, 6, -3, 8, 0, -1, 0, 10,
    -- layer=1 filter=241 channel=47
    3, -9, 9, -10, 5, -10, -9, -1, 0,
    -- layer=1 filter=241 channel=48
    7, -4, 6, -8, -10, -2, -2, -7, -3,
    -- layer=1 filter=241 channel=49
    -9, 8, -8, -6, -6, 5, 4, -3, -2,
    -- layer=1 filter=241 channel=50
    -5, -2, -10, 7, -12, -8, -5, -6, -2,
    -- layer=1 filter=241 channel=51
    -1, 5, -4, 6, -10, -9, 0, -6, -11,
    -- layer=1 filter=241 channel=52
    -1, 3, 6, -6, 1, 6, 5, -7, 11,
    -- layer=1 filter=241 channel=53
    5, -7, -11, -9, 2, 8, -5, -7, -1,
    -- layer=1 filter=241 channel=54
    -2, -3, -9, 10, 8, 2, -9, -9, 1,
    -- layer=1 filter=241 channel=55
    -3, -1, 0, -7, 3, 3, -5, -10, 3,
    -- layer=1 filter=241 channel=56
    -6, -7, -12, 3, -9, -7, 0, -2, -3,
    -- layer=1 filter=241 channel=57
    -7, -10, 5, -5, -4, -2, 6, -12, -10,
    -- layer=1 filter=241 channel=58
    7, 0, 6, 9, -5, 3, -8, 8, -2,
    -- layer=1 filter=241 channel=59
    -4, 4, 0, -3, -10, -9, 5, -3, 0,
    -- layer=1 filter=241 channel=60
    5, -2, -9, -8, 0, 9, -2, 9, 7,
    -- layer=1 filter=241 channel=61
    8, -5, -3, -8, 11, -7, 7, -3, 3,
    -- layer=1 filter=241 channel=62
    2, 8, 9, 5, -2, -5, -1, 1, -4,
    -- layer=1 filter=241 channel=63
    -5, 7, 6, 1, 5, -6, -9, 2, -11,
    -- layer=1 filter=241 channel=64
    -7, 7, -12, 6, -4, 2, -6, 2, 7,
    -- layer=1 filter=241 channel=65
    -8, -7, -1, -3, -5, 7, -8, -8, 3,
    -- layer=1 filter=241 channel=66
    6, -5, -7, 5, -2, -3, -5, -4, 5,
    -- layer=1 filter=241 channel=67
    7, -2, -8, 7, 2, -5, 6, 2, 5,
    -- layer=1 filter=241 channel=68
    -4, -1, 3, -9, -12, -3, 1, 2, 9,
    -- layer=1 filter=241 channel=69
    0, 6, 6, -9, -3, 3, 1, 2, 2,
    -- layer=1 filter=241 channel=70
    4, -8, 8, 0, 5, -4, 11, 5, 5,
    -- layer=1 filter=241 channel=71
    -6, -8, 0, -11, -4, -4, -3, -7, -5,
    -- layer=1 filter=241 channel=72
    -7, 5, 0, 4, -6, -11, -2, 6, 0,
    -- layer=1 filter=241 channel=73
    -6, 0, -4, -10, 1, -1, -11, -5, 2,
    -- layer=1 filter=241 channel=74
    -5, -7, -8, 0, -12, 3, -9, -10, 0,
    -- layer=1 filter=241 channel=75
    6, 9, 3, -8, -7, -2, 0, -2, 5,
    -- layer=1 filter=241 channel=76
    -1, 4, -4, 5, -11, 2, -11, -9, -8,
    -- layer=1 filter=241 channel=77
    -5, -8, -4, -3, -12, -1, 4, -12, -2,
    -- layer=1 filter=241 channel=78
    1, 3, 1, 5, -1, 4, 0, 6, 1,
    -- layer=1 filter=241 channel=79
    0, -5, 2, -1, -6, -2, 2, -8, -1,
    -- layer=1 filter=241 channel=80
    5, 3, 6, -9, -5, -2, 10, 2, 2,
    -- layer=1 filter=241 channel=81
    -4, 5, -12, 4, 7, -6, 5, 4, -3,
    -- layer=1 filter=241 channel=82
    0, 1, -4, 0, -2, -6, 6, -2, 3,
    -- layer=1 filter=241 channel=83
    8, 6, 0, -1, 1, -6, 3, -3, 2,
    -- layer=1 filter=241 channel=84
    0, 9, -6, -2, -9, -10, -7, 5, -9,
    -- layer=1 filter=241 channel=85
    4, -5, 6, -12, 0, -10, -2, -3, -10,
    -- layer=1 filter=241 channel=86
    2, -4, -1, 6, 2, -2, -5, 8, -10,
    -- layer=1 filter=241 channel=87
    2, -7, -10, -11, -10, 5, 2, -3, 6,
    -- layer=1 filter=241 channel=88
    8, -6, 5, 9, -4, -11, 0, -5, -10,
    -- layer=1 filter=241 channel=89
    -8, 5, -8, 3, 3, -4, 2, -9, 7,
    -- layer=1 filter=241 channel=90
    7, 4, -6, 6, -5, 4, 6, -5, -11,
    -- layer=1 filter=241 channel=91
    0, -5, 2, -3, -1, -7, 5, -1, 1,
    -- layer=1 filter=241 channel=92
    -1, 6, 7, -8, 4, 3, 6, -11, -5,
    -- layer=1 filter=241 channel=93
    -9, 3, 5, 3, -10, -1, -7, 1, 0,
    -- layer=1 filter=241 channel=94
    -4, -1, 3, 7, -2, 3, 0, -1, -12,
    -- layer=1 filter=241 channel=95
    7, -5, -5, 7, 4, -11, -1, 8, -4,
    -- layer=1 filter=241 channel=96
    -3, -11, -7, 4, -4, -9, -6, -1, 0,
    -- layer=1 filter=241 channel=97
    -10, -8, 8, -1, 6, 7, 0, 7, 4,
    -- layer=1 filter=241 channel=98
    3, -9, -3, -6, 0, 7, 4, -6, -8,
    -- layer=1 filter=241 channel=99
    4, -5, 4, -7, 0, 7, -9, -6, 3,
    -- layer=1 filter=241 channel=100
    -5, 5, -2, -12, 0, -3, 6, 0, -2,
    -- layer=1 filter=241 channel=101
    -6, 3, -11, 3, 0, -10, -2, 2, 0,
    -- layer=1 filter=241 channel=102
    1, -11, 4, -1, 1, -3, 2, -5, 7,
    -- layer=1 filter=241 channel=103
    8, 4, 3, -1, -4, 8, 1, -3, 1,
    -- layer=1 filter=241 channel=104
    4, 3, -3, -11, 1, -8, -1, 4, 6,
    -- layer=1 filter=241 channel=105
    -1, 3, -7, -5, -4, -12, -4, -8, -1,
    -- layer=1 filter=241 channel=106
    -7, -5, 6, 1, 2, 9, -1, 5, 1,
    -- layer=1 filter=241 channel=107
    5, -1, 7, -2, 2, 5, -1, -11, -3,
    -- layer=1 filter=241 channel=108
    -5, 5, -10, -3, 5, 6, -13, -2, -9,
    -- layer=1 filter=241 channel=109
    8, 0, 5, 2, 4, -9, -1, -8, -1,
    -- layer=1 filter=241 channel=110
    2, 5, -5, -8, -7, -5, -3, -6, 1,
    -- layer=1 filter=241 channel=111
    0, 5, 9, 0, -6, -4, 3, 2, 6,
    -- layer=1 filter=241 channel=112
    -2, -9, 5, -12, -2, 0, -4, -1, -12,
    -- layer=1 filter=241 channel=113
    7, 9, 8, 1, -9, 0, -8, -5, -8,
    -- layer=1 filter=241 channel=114
    -11, 6, -12, -5, 0, 8, -4, 5, 9,
    -- layer=1 filter=241 channel=115
    5, -3, -10, -11, 1, 7, -4, 1, -4,
    -- layer=1 filter=241 channel=116
    8, -9, 2, -7, 5, 7, 1, -6, 7,
    -- layer=1 filter=241 channel=117
    -8, 1, -1, 4, 8, -4, 8, -8, 5,
    -- layer=1 filter=241 channel=118
    2, -6, -7, -5, 4, 3, -5, 0, 8,
    -- layer=1 filter=241 channel=119
    4, -3, -2, -4, -9, -12, 4, 8, -3,
    -- layer=1 filter=241 channel=120
    8, 5, 3, -6, 6, 1, 3, 7, 3,
    -- layer=1 filter=241 channel=121
    -9, -4, 1, 8, -10, -4, -1, -6, -10,
    -- layer=1 filter=241 channel=122
    4, -4, 2, -5, -3, 7, 10, -3, -9,
    -- layer=1 filter=241 channel=123
    -3, 5, 4, 3, -4, 0, -7, 0, -1,
    -- layer=1 filter=241 channel=124
    -2, 3, -4, -6, -1, -10, -5, 4, -1,
    -- layer=1 filter=241 channel=125
    -10, 1, -7, 9, 7, 7, 0, -7, -10,
    -- layer=1 filter=241 channel=126
    3, 8, 4, 2, 3, -5, 0, 0, 0,
    -- layer=1 filter=241 channel=127
    -12, 0, -6, 2, -1, 0, -3, 0, 5,
    -- layer=1 filter=242 channel=0
    -11, -23, -21, -5, 0, -11, 4, 4, -7,
    -- layer=1 filter=242 channel=1
    -2, 6, 6, 10, -16, 14, 23, 11, 19,
    -- layer=1 filter=242 channel=2
    -15, -9, 36, -17, 3, 44, 1, 26, 20,
    -- layer=1 filter=242 channel=3
    0, -5, 2, -2, -1, -4, -12, -6, 2,
    -- layer=1 filter=242 channel=4
    -8, -1, -10, 1, 3, -6, 0, -10, -5,
    -- layer=1 filter=242 channel=5
    0, 2, 3, 2, -8, 35, 32, 10, 11,
    -- layer=1 filter=242 channel=6
    5, -24, 2, -5, -5, -1, -26, -4, 2,
    -- layer=1 filter=242 channel=7
    -51, -69, -32, -46, -76, -39, -38, -38, 16,
    -- layer=1 filter=242 channel=8
    2, 12, 11, 25, -17, 29, 11, 8, 18,
    -- layer=1 filter=242 channel=9
    -6, 8, 7, -27, -21, 21, -9, 5, 36,
    -- layer=1 filter=242 channel=10
    -71, -53, -46, -45, -76, -14, -24, -7, 6,
    -- layer=1 filter=242 channel=11
    -18, -15, -14, -8, -13, -14, -33, -15, -29,
    -- layer=1 filter=242 channel=12
    -79, -44, -26, -48, -40, 30, -24, -23, -6,
    -- layer=1 filter=242 channel=13
    2, 1, -1, -11, 6, 15, -6, -8, 9,
    -- layer=1 filter=242 channel=14
    -69, -44, -14, -51, -45, -63, -27, -54, 9,
    -- layer=1 filter=242 channel=15
    -27, 0, 13, -2, -33, 17, -50, -43, 4,
    -- layer=1 filter=242 channel=16
    -3, 11, 1, -2, -8, 25, -1, -7, 14,
    -- layer=1 filter=242 channel=17
    -5, -6, -21, 8, -12, -2, 6, -3, 2,
    -- layer=1 filter=242 channel=18
    -9, -17, -14, -17, -39, -2, -22, -13, 13,
    -- layer=1 filter=242 channel=19
    -30, 8, 2, 14, 3, 62, 2, 33, 36,
    -- layer=1 filter=242 channel=20
    11, 0, -1, 1, 0, 18, 0, -3, 10,
    -- layer=1 filter=242 channel=21
    -3, -18, 0, 8, -5, -7, -3, 9, 10,
    -- layer=1 filter=242 channel=22
    -1, 11, 16, -8, 0, 15, 1, -4, 16,
    -- layer=1 filter=242 channel=23
    -2, -45, 9, -19, -31, -3, -1, -7, 12,
    -- layer=1 filter=242 channel=24
    -5, 21, 9, 12, 12, 28, -9, 19, 15,
    -- layer=1 filter=242 channel=25
    -45, -29, -17, -25, -42, 6, -10, 23, 24,
    -- layer=1 filter=242 channel=26
    -15, 7, 16, -14, -4, 19, -7, -1, 7,
    -- layer=1 filter=242 channel=27
    -18, -18, 15, -6, 4, -2, -20, -22, -33,
    -- layer=1 filter=242 channel=28
    -41, -40, -18, -52, -42, -28, -28, -3, 0,
    -- layer=1 filter=242 channel=29
    -6, -12, -5, -4, -9, -14, -8, -18, -6,
    -- layer=1 filter=242 channel=30
    -15, -25, -28, 4, -21, 13, -7, 16, 28,
    -- layer=1 filter=242 channel=31
    -30, -16, 16, -25, -1, -13, 6, 9, 12,
    -- layer=1 filter=242 channel=32
    -11, -19, 11, -26, -20, 13, -15, 17, 24,
    -- layer=1 filter=242 channel=33
    -10, -7, 10, 2, -7, 3, -2, 21, 4,
    -- layer=1 filter=242 channel=34
    -18, -19, 5, -22, -7, -13, -13, -19, -8,
    -- layer=1 filter=242 channel=35
    2, 1, 11, 15, 1, 8, 13, 3, 8,
    -- layer=1 filter=242 channel=36
    -29, -24, -25, -10, -17, -18, -27, -10, -27,
    -- layer=1 filter=242 channel=37
    -8, -13, 2, 0, 2, 20, 11, -2, 3,
    -- layer=1 filter=242 channel=38
    4, 1, 0, 9, 3, 10, 5, 18, 10,
    -- layer=1 filter=242 channel=39
    -4, -3, -4, -19, -4, -10, 2, -5, -19,
    -- layer=1 filter=242 channel=40
    6, -25, 7, 11, -4, -20, -21, -4, 0,
    -- layer=1 filter=242 channel=41
    -32, 7, 35, 0, -22, -6, -22, 32, 60,
    -- layer=1 filter=242 channel=42
    -26, -13, 22, -4, -4, 24, 0, -3, 27,
    -- layer=1 filter=242 channel=43
    -11, 7, 0, 3, 0, 18, 2, 2, 4,
    -- layer=1 filter=242 channel=44
    -6, -19, 13, -22, -20, 21, 18, -2, 24,
    -- layer=1 filter=242 channel=45
    0, 15, -1, 0, 7, 29, 0, -3, 10,
    -- layer=1 filter=242 channel=46
    -34, -12, 8, -3, 0, 27, 1, -11, 5,
    -- layer=1 filter=242 channel=47
    -16, -30, 30, -22, -4, -1, -15, 15, 46,
    -- layer=1 filter=242 channel=48
    -7, -4, -27, 10, 0, -4, 4, 22, 8,
    -- layer=1 filter=242 channel=49
    -13, -8, 17, -14, 1, 19, 3, 14, 30,
    -- layer=1 filter=242 channel=50
    -17, -5, 8, -18, -11, -3, -8, 11, 0,
    -- layer=1 filter=242 channel=51
    -16, -15, -27, -2, -21, -31, 0, 8, -2,
    -- layer=1 filter=242 channel=52
    -8, 4, 1, 4, 11, 5, -3, 6, 7,
    -- layer=1 filter=242 channel=53
    0, -8, -21, -23, -7, -19, -13, -4, -12,
    -- layer=1 filter=242 channel=54
    -36, -21, -16, -17, -39, 22, -9, 32, 10,
    -- layer=1 filter=242 channel=55
    4, -3, 15, -3, -12, 2, -6, 4, -3,
    -- layer=1 filter=242 channel=56
    11, -2, -11, 8, -10, -9, 0, -8, -1,
    -- layer=1 filter=242 channel=57
    -46, -40, -29, -7, -63, -15, -23, -16, -3,
    -- layer=1 filter=242 channel=58
    -42, -39, -1, -12, -32, 36, -45, 22, 11,
    -- layer=1 filter=242 channel=59
    5, 8, 1, 0, 6, -4, 2, 0, -1,
    -- layer=1 filter=242 channel=60
    0, 18, 14, 13, 11, 1, 9, -2, -3,
    -- layer=1 filter=242 channel=61
    -5, -14, 8, -2, 4, -1, -2, -9, 0,
    -- layer=1 filter=242 channel=62
    4, 3, -5, 9, -11, 33, 18, 24, 9,
    -- layer=1 filter=242 channel=63
    -4, -6, -21, -2, 10, 0, 9, 10, -2,
    -- layer=1 filter=242 channel=64
    9, 5, 0, 1, -6, -4, -2, 8, 8,
    -- layer=1 filter=242 channel=65
    -1, -8, -21, 1, 0, -20, 14, 5, -5,
    -- layer=1 filter=242 channel=66
    6, 6, -9, 12, 2, -7, 17, 8, 10,
    -- layer=1 filter=242 channel=67
    -14, -6, -9, -23, -35, -32, -33, -31, -57,
    -- layer=1 filter=242 channel=68
    -22, -8, 8, -30, -14, 32, 9, 0, 20,
    -- layer=1 filter=242 channel=69
    -20, 0, 27, 1, -30, 35, -9, -26, 15,
    -- layer=1 filter=242 channel=70
    -25, -37, -12, -19, -34, -25, -18, -19, -16,
    -- layer=1 filter=242 channel=71
    -10, -1, -4, 0, 0, -4, 10, 6, 1,
    -- layer=1 filter=242 channel=72
    -17, -4, -11, -3, -20, 31, -11, 22, 24,
    -- layer=1 filter=242 channel=73
    12, -2, 2, 1, -2, -3, 6, 0, -4,
    -- layer=1 filter=242 channel=74
    13, -17, -4, -14, 15, 22, 9, 22, 7,
    -- layer=1 filter=242 channel=75
    -20, -31, -10, -51, -10, 0, -15, -2, -30,
    -- layer=1 filter=242 channel=76
    -3, -26, -22, -13, -14, 3, 8, 13, -4,
    -- layer=1 filter=242 channel=77
    4, -7, -19, 0, -8, -24, -6, 13, 0,
    -- layer=1 filter=242 channel=78
    -21, -6, -6, 10, 4, 1, -10, -4, -10,
    -- layer=1 filter=242 channel=79
    7, 3, 9, 0, -13, 39, 3, 0, 14,
    -- layer=1 filter=242 channel=80
    -1, -6, -7, 5, 2, 0, -1, -15, 1,
    -- layer=1 filter=242 channel=81
    13, -2, -7, 4, 15, -8, -4, 5, -4,
    -- layer=1 filter=242 channel=82
    11, -8, -7, -3, 10, -9, 6, 4, 1,
    -- layer=1 filter=242 channel=83
    -7, -27, 4, 0, -21, 0, 2, -45, -10,
    -- layer=1 filter=242 channel=84
    9, -11, 0, -21, 7, 15, 10, 40, 24,
    -- layer=1 filter=242 channel=85
    -41, -24, 4, -2, -11, 32, -18, 20, 23,
    -- layer=1 filter=242 channel=86
    11, -5, -9, -3, -4, -15, -10, -20, -15,
    -- layer=1 filter=242 channel=87
    -33, 10, 41, -20, 12, 40, 17, 13, 40,
    -- layer=1 filter=242 channel=88
    -4, -10, -6, -15, 3, -12, 0, -3, -11,
    -- layer=1 filter=242 channel=89
    4, -5, 1, 0, -2, 2, 13, 2, -7,
    -- layer=1 filter=242 channel=90
    -28, -21, 0, -22, -30, 7, 6, -10, 9,
    -- layer=1 filter=242 channel=91
    -2, -6, -8, 5, -4, 9, -8, 14, 8,
    -- layer=1 filter=242 channel=92
    -37, -19, -2, -26, -14, -25, -33, 9, 32,
    -- layer=1 filter=242 channel=93
    5, 10, -10, 11, 4, -1, 22, 24, 7,
    -- layer=1 filter=242 channel=94
    -25, -16, -20, -3, -2, -5, -6, 1, 0,
    -- layer=1 filter=242 channel=95
    -8, -28, 3, -20, 8, 10, 12, 36, 20,
    -- layer=1 filter=242 channel=96
    2, -4, -5, -3, -2, -1, -1, -6, -7,
    -- layer=1 filter=242 channel=97
    -5, 3, 1, 7, 7, -3, 5, 5, 4,
    -- layer=1 filter=242 channel=98
    -4, -3, -8, -7, 0, 20, -14, 0, 15,
    -- layer=1 filter=242 channel=99
    -43, -21, -27, -54, -65, -33, -13, 18, 16,
    -- layer=1 filter=242 channel=100
    -6, -21, -24, -13, -13, -18, 6, 11, -6,
    -- layer=1 filter=242 channel=101
    0, -2, -12, 8, 8, 5, 13, 16, 20,
    -- layer=1 filter=242 channel=102
    -9, -15, -14, -11, -15, -10, 1, 9, 0,
    -- layer=1 filter=242 channel=103
    -14, -14, 12, 1, 9, 15, -7, 16, 0,
    -- layer=1 filter=242 channel=104
    -4, -11, 24, -11, -10, 15, -3, 17, 2,
    -- layer=1 filter=242 channel=105
    0, -1, -5, 1, -9, -8, 14, 12, 2,
    -- layer=1 filter=242 channel=106
    0, 5, 11, -4, 8, 3, 14, 14, 23,
    -- layer=1 filter=242 channel=107
    4, 8, -5, 0, -1, 3, -10, -7, 5,
    -- layer=1 filter=242 channel=108
    -18, -17, 10, -25, -27, 24, -8, 0, 25,
    -- layer=1 filter=242 channel=109
    -6, 9, -7, 8, -1, 7, -5, -8, -8,
    -- layer=1 filter=242 channel=110
    -4, -13, -15, 0, -3, -5, -4, -2, 2,
    -- layer=1 filter=242 channel=111
    -9, -34, -27, 10, -34, 22, -13, 19, 27,
    -- layer=1 filter=242 channel=112
    8, -22, 4, 0, 5, 21, 11, 32, 21,
    -- layer=1 filter=242 channel=113
    -27, -23, 9, -5, -13, 1, -3, -1, 15,
    -- layer=1 filter=242 channel=114
    -51, -41, -27, -31, -45, -33, -5, -29, -29,
    -- layer=1 filter=242 channel=115
    -6, -22, -21, -11, -22, -3, -6, -7, -16,
    -- layer=1 filter=242 channel=116
    -9, -5, -5, 0, 0, 5, -6, -8, -7,
    -- layer=1 filter=242 channel=117
    -44, -42, -6, -11, -22, 11, -35, -6, -9,
    -- layer=1 filter=242 channel=118
    -8, -6, -22, 9, 2, 33, 11, 37, 16,
    -- layer=1 filter=242 channel=119
    -26, 1, 11, -25, -14, 26, 0, -4, 17,
    -- layer=1 filter=242 channel=120
    0, -2, -1, 0, -2, -6, 8, 12, 17,
    -- layer=1 filter=242 channel=121
    -28, -24, -11, -39, -49, 1, -14, -10, -11,
    -- layer=1 filter=242 channel=122
    -5, 3, -6, -5, -6, 2, -6, 0, 0,
    -- layer=1 filter=242 channel=123
    -7, -35, -14, -24, -23, -5, -13, -5, -1,
    -- layer=1 filter=242 channel=124
    4, -5, 5, 4, 4, -10, -14, -10, -7,
    -- layer=1 filter=242 channel=125
    -9, -33, -13, -12, -22, -26, -9, -10, -2,
    -- layer=1 filter=242 channel=126
    27, 7, 14, 3, -1, 15, 18, -4, 28,
    -- layer=1 filter=242 channel=127
    13, -22, -19, -7, -6, 22, 5, 27, 20,
    -- layer=1 filter=243 channel=0
    0, 7, 7, 10, 9, 6, 15, 17, 6,
    -- layer=1 filter=243 channel=1
    -7, -58, -24, -21, -22, 7, -40, -11, 33,
    -- layer=1 filter=243 channel=2
    4, 1, 5, 13, 28, 25, 23, 19, 28,
    -- layer=1 filter=243 channel=3
    2, 0, 11, -9, 2, -5, 5, -9, -7,
    -- layer=1 filter=243 channel=4
    1, 10, 0, -9, 4, -2, -2, 14, 1,
    -- layer=1 filter=243 channel=5
    -8, -45, -10, -87, -55, -33, -13, 18, 48,
    -- layer=1 filter=243 channel=6
    0, 1, -7, -31, -14, -27, 9, -9, -3,
    -- layer=1 filter=243 channel=7
    -62, -112, -96, -79, -126, -109, 18, -41, -48,
    -- layer=1 filter=243 channel=8
    -41, -75, -25, -61, -65, -13, -20, 32, 45,
    -- layer=1 filter=243 channel=9
    -6, 0, 15, -37, 31, -1, 41, 28, 36,
    -- layer=1 filter=243 channel=10
    -79, -101, -77, -65, -122, -65, 62, -50, -33,
    -- layer=1 filter=243 channel=11
    1, 11, 9, 20, 18, 7, 10, 6, -7,
    -- layer=1 filter=243 channel=12
    -30, 3, 3, -70, 11, 39, 2, 27, 29,
    -- layer=1 filter=243 channel=13
    -11, 0, 3, -5, 1, 3, 3, 0, 19,
    -- layer=1 filter=243 channel=14
    -15, -40, 2, -48, -66, -34, 11, -58, -64,
    -- layer=1 filter=243 channel=15
    12, -9, 3, -41, -60, 6, -28, 10, 26,
    -- layer=1 filter=243 channel=16
    -42, -64, -12, -59, -49, 6, 23, 50, 58,
    -- layer=1 filter=243 channel=17
    0, 16, 2, 22, -1, 2, 8, 22, 7,
    -- layer=1 filter=243 channel=18
    -42, -32, -7, 0, 33, 23, 31, -8, 13,
    -- layer=1 filter=243 channel=19
    -33, -28, -22, -47, -98, -8, 49, 21, 45,
    -- layer=1 filter=243 channel=20
    -2, 0, 6, -9, 0, 6, -6, 32, 23,
    -- layer=1 filter=243 channel=21
    -23, -14, 0, -19, 4, 0, -1, 12, 32,
    -- layer=1 filter=243 channel=22
    17, 1, 28, 25, 10, 19, 17, 21, 33,
    -- layer=1 filter=243 channel=23
    4, -13, -31, -39, -26, -28, -51, -29, 0,
    -- layer=1 filter=243 channel=24
    -26, -21, -8, -35, -15, 15, 4, 24, 33,
    -- layer=1 filter=243 channel=25
    -68, -74, -82, -79, -104, -36, 8, 32, 4,
    -- layer=1 filter=243 channel=26
    -16, -42, 13, -19, -24, 16, -32, 25, 9,
    -- layer=1 filter=243 channel=27
    25, 38, 23, 49, 59, 34, 39, 28, 26,
    -- layer=1 filter=243 channel=28
    -23, -52, -65, -36, -63, -43, 38, -23, -21,
    -- layer=1 filter=243 channel=29
    29, 42, 25, 18, 35, 41, -5, 0, -3,
    -- layer=1 filter=243 channel=30
    -90, -105, -12, -10, -27, 2, 18, -23, 7,
    -- layer=1 filter=243 channel=31
    -10, -23, 7, -5, 29, 13, -2, -4, 2,
    -- layer=1 filter=243 channel=32
    -22, -91, 11, -37, -52, 12, -77, -35, 7,
    -- layer=1 filter=243 channel=33
    -13, 2, -16, 2, -8, 0, -1, 14, 0,
    -- layer=1 filter=243 channel=34
    14, 25, 14, 22, 19, 35, 24, 21, -4,
    -- layer=1 filter=243 channel=35
    -9, 0, -1, -4, 1, -6, -2, -1, 1,
    -- layer=1 filter=243 channel=36
    25, 8, 8, 22, 33, 19, 12, 6, -7,
    -- layer=1 filter=243 channel=37
    -16, -35, -6, -74, -57, 0, 11, 44, 52,
    -- layer=1 filter=243 channel=38
    -5, -5, -3, -1, -3, 13, 16, 12, 14,
    -- layer=1 filter=243 channel=39
    3, 21, -3, 8, 10, -3, 13, 13, 0,
    -- layer=1 filter=243 channel=40
    -37, -20, -25, -19, -15, -14, 47, -17, -11,
    -- layer=1 filter=243 channel=41
    13, -11, 14, -23, 31, 28, 7, -3, 24,
    -- layer=1 filter=243 channel=42
    6, 21, 1, 9, 16, 8, 29, 14, 12,
    -- layer=1 filter=243 channel=43
    -42, -101, -34, -61, -64, -13, -26, 34, 37,
    -- layer=1 filter=243 channel=44
    -63, -91, 5, -70, -50, 19, -73, -7, 18,
    -- layer=1 filter=243 channel=45
    -8, -30, -12, -19, -24, 9, -22, 13, 40,
    -- layer=1 filter=243 channel=46
    -25, -2, 39, -125, -71, -16, 69, 51, 64,
    -- layer=1 filter=243 channel=47
    1, -16, -32, -49, -31, -26, -49, -53, -10,
    -- layer=1 filter=243 channel=48
    -26, -7, 0, -16, 4, 10, -5, -7, -1,
    -- layer=1 filter=243 channel=49
    -22, -11, -24, -9, -9, 16, 1, 10, 4,
    -- layer=1 filter=243 channel=50
    -10, -15, -17, -1, -1, -1, -23, -9, -12,
    -- layer=1 filter=243 channel=51
    -38, -6, -20, -10, -8, -4, 47, 10, 3,
    -- layer=1 filter=243 channel=52
    22, -7, 4, -2, -7, -9, 8, 13, -1,
    -- layer=1 filter=243 channel=53
    -23, -20, -8, -22, -17, -4, -23, -12, -14,
    -- layer=1 filter=243 channel=54
    -45, -54, -55, -87, -69, -27, 39, 48, 34,
    -- layer=1 filter=243 channel=55
    7, 20, 6, 22, 29, -1, 0, 9, -8,
    -- layer=1 filter=243 channel=56
    1, -3, 3, 7, 0, -4, 0, -5, -1,
    -- layer=1 filter=243 channel=57
    -63, -49, -69, -45, -75, -50, 89, -30, -26,
    -- layer=1 filter=243 channel=58
    -69, -97, -69, -148, -121, -46, 17, 0, -36,
    -- layer=1 filter=243 channel=59
    -6, -1, -7, -2, 1, -1, -9, -13, 1,
    -- layer=1 filter=243 channel=60
    -1, 11, 17, -1, -2, 8, -6, -5, 11,
    -- layer=1 filter=243 channel=61
    10, -4, -5, -7, 10, 6, 9, 4, -1,
    -- layer=1 filter=243 channel=62
    -75, -82, -30, -100, -76, -8, 1, 43, 55,
    -- layer=1 filter=243 channel=63
    4, 9, -2, 31, 17, 12, 5, 11, -15,
    -- layer=1 filter=243 channel=64
    16, 14, 6, 5, 14, 10, -2, 10, 26,
    -- layer=1 filter=243 channel=65
    -7, 0, 1, -16, 11, 9, 11, 1, 12,
    -- layer=1 filter=243 channel=66
    20, 12, -3, 21, 12, 13, 5, -5, -14,
    -- layer=1 filter=243 channel=67
    -34, -38, -59, -37, -36, -21, -8, -19, -8,
    -- layer=1 filter=243 channel=68
    -56, -99, 19, -64, -30, 30, -61, 3, 18,
    -- layer=1 filter=243 channel=69
    14, -19, -2, -43, -55, -8, 17, 59, 60,
    -- layer=1 filter=243 channel=70
    -38, -27, -49, -3, 5, -2, 51, 10, -22,
    -- layer=1 filter=243 channel=71
    -15, -9, -1, -22, -12, 0, -10, 15, 8,
    -- layer=1 filter=243 channel=72
    -42, -25, 18, -43, -18, 1, 15, -1, 19,
    -- layer=1 filter=243 channel=73
    -10, 0, -2, -9, 0, 1, 6, 8, 8,
    -- layer=1 filter=243 channel=74
    -65, -52, 61, -24, -21, 32, -31, -9, 30,
    -- layer=1 filter=243 channel=75
    -55, -41, 27, -36, 13, 38, -14, 13, 17,
    -- layer=1 filter=243 channel=76
    -15, -24, 12, 5, 7, 29, -13, 25, 19,
    -- layer=1 filter=243 channel=77
    -33, -17, -15, -10, -7, 0, -15, -16, 7,
    -- layer=1 filter=243 channel=78
    5, -3, -21, -10, -17, -12, 3, -6, -7,
    -- layer=1 filter=243 channel=79
    -21, -42, 10, -55, -27, 5, 11, 41, 64,
    -- layer=1 filter=243 channel=80
    -2, 8, -3, 8, 11, 14, -5, 1, -5,
    -- layer=1 filter=243 channel=81
    -6, -12, -8, -15, -3, 4, -10, 20, 13,
    -- layer=1 filter=243 channel=82
    -19, -8, -2, -2, -7, 5, 0, 13, 22,
    -- layer=1 filter=243 channel=83
    -7, -22, 5, -2, -10, 14, -21, 1, 23,
    -- layer=1 filter=243 channel=84
    -114, -89, 11, -13, 14, 33, -3, 5, 25,
    -- layer=1 filter=243 channel=85
    1, -25, -15, -59, -19, -16, -20, -11, -25,
    -- layer=1 filter=243 channel=86
    22, 17, 12, 21, 8, 9, 3, -1, -13,
    -- layer=1 filter=243 channel=87
    -28, -25, -2, -54, -14, 0, 89, 20, 59,
    -- layer=1 filter=243 channel=88
    -5, -8, -2, 5, 12, 1, 21, 17, 13,
    -- layer=1 filter=243 channel=89
    -13, -24, 8, 0, -5, 3, -18, -7, 33,
    -- layer=1 filter=243 channel=90
    -55, -88, -14, -97, -65, 13, -57, -19, 8,
    -- layer=1 filter=243 channel=91
    3, 5, 6, 9, -10, 9, 26, 17, 9,
    -- layer=1 filter=243 channel=92
    5, 2, 12, -10, 1, 27, 19, 36, 5,
    -- layer=1 filter=243 channel=93
    -12, 6, 5, -10, 2, 1, -1, 19, 19,
    -- layer=1 filter=243 channel=94
    12, 1, 8, 21, 2, 16, 7, 14, 7,
    -- layer=1 filter=243 channel=95
    -123, -94, 6, -24, -16, -1, -32, -18, 24,
    -- layer=1 filter=243 channel=96
    21, 21, 8, 19, 12, 7, 8, 11, 15,
    -- layer=1 filter=243 channel=97
    0, 4, -1, 14, 10, 14, 11, 19, -1,
    -- layer=1 filter=243 channel=98
    -28, -46, -8, -16, -9, 1, -23, 22, 51,
    -- layer=1 filter=243 channel=99
    -54, -65, -18, 17, -107, -49, 53, -59, -22,
    -- layer=1 filter=243 channel=100
    0, 15, 14, 9, 32, 17, 0, -13, -19,
    -- layer=1 filter=243 channel=101
    0, 2, 8, -11, 10, -5, 0, 13, 32,
    -- layer=1 filter=243 channel=102
    6, 15, 10, 14, 14, 20, 20, 19, 15,
    -- layer=1 filter=243 channel=103
    13, 15, 9, 18, 45, 19, -5, 2, -5,
    -- layer=1 filter=243 channel=104
    -10, 7, -27, -20, 9, -26, -20, -7, -17,
    -- layer=1 filter=243 channel=105
    -1, 6, 3, 15, 12, 12, 11, -2, 0,
    -- layer=1 filter=243 channel=106
    -27, -13, -2, 0, -20, -2, -18, -8, 10,
    -- layer=1 filter=243 channel=107
    -3, -1, 0, 9, 5, -4, 13, 14, 6,
    -- layer=1 filter=243 channel=108
    -43, -113, -18, -74, -99, -2, -60, -32, 24,
    -- layer=1 filter=243 channel=109
    1, -9, -2, -10, 7, -2, 3, 3, 8,
    -- layer=1 filter=243 channel=110
    -1, -1, -2, 3, 0, 3, 14, -7, 5,
    -- layer=1 filter=243 channel=111
    -91, -76, 4, -13, 15, 17, 37, 9, 37,
    -- layer=1 filter=243 channel=112
    -36, -20, 1, 11, 31, 38, 3, 24, 29,
    -- layer=1 filter=243 channel=113
    -2, -10, -13, -21, -2, -3, 7, 11, -2,
    -- layer=1 filter=243 channel=114
    20, -1, 4, 7, -10, 10, 12, 51, 59,
    -- layer=1 filter=243 channel=115
    5, 12, -1, -1, 7, 4, 34, 5, 10,
    -- layer=1 filter=243 channel=116
    10, -9, 9, 5, -5, 8, -1, 2, 3,
    -- layer=1 filter=243 channel=117
    -74, -62, 12, 13, 23, 36, 52, 41, 19,
    -- layer=1 filter=243 channel=118
    -77, -77, 3, -4, 0, 23, 2, -17, 28,
    -- layer=1 filter=243 channel=119
    -29, -78, -17, -56, -68, 13, -64, -40, 18,
    -- layer=1 filter=243 channel=120
    -7, -11, -8, -15, -7, 8, 23, 22, 31,
    -- layer=1 filter=243 channel=121
    6, 17, 22, -11, 16, 12, 6, -18, -32,
    -- layer=1 filter=243 channel=122
    -10, 1, -5, 0, -3, -3, -7, -2, 5,
    -- layer=1 filter=243 channel=123
    11, 34, 12, 6, 36, 14, 16, 6, -2,
    -- layer=1 filter=243 channel=124
    -12, -7, 3, -4, -7, -8, 6, -6, -8,
    -- layer=1 filter=243 channel=125
    -47, -53, -44, -5, -19, -35, 39, 11, -21,
    -- layer=1 filter=243 channel=126
    -77, -87, -32, -51, -50, -26, -62, -15, 6,
    -- layer=1 filter=243 channel=127
    -87, -75, 20, -2, -1, 8, -11, -8, 32,
    -- layer=1 filter=244 channel=0
    7, -4, -6, -2, 6, 6, -3, 0, 7,
    -- layer=1 filter=244 channel=1
    -10, -10, 3, -7, -4, -2, 2, -8, 5,
    -- layer=1 filter=244 channel=2
    3, 4, 10, 8, 8, 8, 7, 0, 9,
    -- layer=1 filter=244 channel=3
    -10, 10, 6, 7, -5, -1, 2, 0, 6,
    -- layer=1 filter=244 channel=4
    0, -11, -6, -7, -3, 2, -2, -2, -4,
    -- layer=1 filter=244 channel=5
    -8, 1, 0, -8, 5, 1, -4, -1, 0,
    -- layer=1 filter=244 channel=6
    5, 2, 9, -8, 2, 0, 0, -9, -7,
    -- layer=1 filter=244 channel=7
    0, -2, -1, -7, -2, 4, 5, -11, 9,
    -- layer=1 filter=244 channel=8
    -7, -2, -10, 8, 2, -9, -8, 3, 0,
    -- layer=1 filter=244 channel=9
    8, 1, -7, -8, 1, -11, -5, 7, -6,
    -- layer=1 filter=244 channel=10
    -6, -7, 8, -7, -7, -9, -12, 7, 3,
    -- layer=1 filter=244 channel=11
    -2, -7, 4, -1, -11, -1, -9, -5, -4,
    -- layer=1 filter=244 channel=12
    7, 7, 4, -9, 0, 9, -9, 6, 5,
    -- layer=1 filter=244 channel=13
    -1, -4, 0, -11, 1, -9, -6, -8, 7,
    -- layer=1 filter=244 channel=14
    -1, -8, -7, 1, 6, -1, 7, -1, -7,
    -- layer=1 filter=244 channel=15
    -6, -8, 4, 10, 0, -3, 11, -1, -2,
    -- layer=1 filter=244 channel=16
    5, -10, -6, -12, -4, 5, 7, -8, -4,
    -- layer=1 filter=244 channel=17
    -1, -2, -10, 1, -5, 8, 1, 7, -10,
    -- layer=1 filter=244 channel=18
    -1, 6, -2, -12, -8, 0, -4, 8, 9,
    -- layer=1 filter=244 channel=19
    0, 2, 0, 8, -1, 7, 1, -10, -6,
    -- layer=1 filter=244 channel=20
    7, 4, 0, -9, 7, 2, 6, -3, 0,
    -- layer=1 filter=244 channel=21
    -9, 5, -6, -4, -1, -11, -5, 3, 1,
    -- layer=1 filter=244 channel=22
    7, -10, -7, -2, -11, 1, 1, -3, -8,
    -- layer=1 filter=244 channel=23
    6, -1, 5, -6, 5, -8, 8, -12, -1,
    -- layer=1 filter=244 channel=24
    -8, 3, 1, -8, -1, 4, -6, -12, 3,
    -- layer=1 filter=244 channel=25
    -11, 3, 7, -3, 0, -10, 5, 3, -2,
    -- layer=1 filter=244 channel=26
    2, 1, -5, -1, -8, -9, 4, 0, -2,
    -- layer=1 filter=244 channel=27
    6, -5, 0, -7, -5, -9, 5, -8, 5,
    -- layer=1 filter=244 channel=28
    6, -5, -7, -6, 8, -12, -1, 5, 1,
    -- layer=1 filter=244 channel=29
    -5, 0, -11, -9, 10, -6, 9, -10, -6,
    -- layer=1 filter=244 channel=30
    7, 0, 0, -8, 6, 0, -4, -1, -3,
    -- layer=1 filter=244 channel=31
    -8, 3, -6, -11, 0, 0, -9, -8, -2,
    -- layer=1 filter=244 channel=32
    3, -8, -1, 1, 4, 1, 0, -3, -2,
    -- layer=1 filter=244 channel=33
    -2, -7, -8, 8, 0, -6, -3, 0, -7,
    -- layer=1 filter=244 channel=34
    7, -6, 2, 5, -2, 7, 7, -2, -6,
    -- layer=1 filter=244 channel=35
    -7, -9, 6, 7, 6, 5, -5, -12, 2,
    -- layer=1 filter=244 channel=36
    1, -5, 3, 5, -1, 1, 5, 2, -7,
    -- layer=1 filter=244 channel=37
    -1, 6, -6, 0, 4, 8, 0, 0, 0,
    -- layer=1 filter=244 channel=38
    5, 7, -3, -2, -6, -2, 4, -8, -1,
    -- layer=1 filter=244 channel=39
    -2, -7, -7, 2, -8, -11, 4, 6, 8,
    -- layer=1 filter=244 channel=40
    -11, 1, -6, -1, -5, 2, 0, 3, -4,
    -- layer=1 filter=244 channel=41
    8, -12, -3, -1, -8, 3, 0, -9, -4,
    -- layer=1 filter=244 channel=42
    3, 1, 5, 0, 8, -2, -3, 5, -4,
    -- layer=1 filter=244 channel=43
    6, -8, 3, -8, 5, 6, 8, -10, -6,
    -- layer=1 filter=244 channel=44
    -2, -8, -5, -3, 1, 2, 2, -6, 0,
    -- layer=1 filter=244 channel=45
    3, -5, -8, 1, -1, -9, -8, 0, -6,
    -- layer=1 filter=244 channel=46
    2, 0, 5, 2, 6, 8, 10, -6, 9,
    -- layer=1 filter=244 channel=47
    -4, -2, 1, -3, -9, 8, 3, 1, -10,
    -- layer=1 filter=244 channel=48
    6, -3, -3, -10, 4, -6, 5, 0, 0,
    -- layer=1 filter=244 channel=49
    0, -7, -10, -7, -11, 9, 0, 7, -7,
    -- layer=1 filter=244 channel=50
    7, 6, -9, 0, -3, -10, -11, -1, 0,
    -- layer=1 filter=244 channel=51
    0, 0, -6, 2, 2, 5, -7, 3, -1,
    -- layer=1 filter=244 channel=52
    2, -9, -4, -9, -9, 9, -7, 9, 0,
    -- layer=1 filter=244 channel=53
    -9, 5, 4, 0, -8, -8, -12, -1, 8,
    -- layer=1 filter=244 channel=54
    -3, -9, -7, -2, -12, 3, -4, 4, -2,
    -- layer=1 filter=244 channel=55
    8, 2, -5, -8, 3, 1, -11, -10, 8,
    -- layer=1 filter=244 channel=56
    -11, 0, 4, 7, -2, 6, -8, -4, 3,
    -- layer=1 filter=244 channel=57
    6, -9, -6, 4, -7, 5, -10, -9, -12,
    -- layer=1 filter=244 channel=58
    0, 9, 1, -9, 3, 11, -9, -7, -9,
    -- layer=1 filter=244 channel=59
    -11, 7, 7, 4, 5, -7, -11, -3, 6,
    -- layer=1 filter=244 channel=60
    9, 0, 7, 0, -2, 3, -2, 11, -7,
    -- layer=1 filter=244 channel=61
    2, 8, 7, 10, 1, -7, 3, 7, -11,
    -- layer=1 filter=244 channel=62
    5, 2, -10, 6, 5, -7, 6, -12, 2,
    -- layer=1 filter=244 channel=63
    -5, 4, 5, -3, 7, -9, -8, 5, -5,
    -- layer=1 filter=244 channel=64
    2, -9, 8, -11, -4, 8, -1, -1, -1,
    -- layer=1 filter=244 channel=65
    6, -8, -8, 1, 5, 7, 2, 8, 1,
    -- layer=1 filter=244 channel=66
    -7, 7, 0, 0, -4, -6, -1, -9, 4,
    -- layer=1 filter=244 channel=67
    1, -1, 3, -8, 2, 1, 4, -5, 2,
    -- layer=1 filter=244 channel=68
    0, 0, 4, -10, -9, 0, 0, -8, -11,
    -- layer=1 filter=244 channel=69
    -8, -8, -6, -3, -1, -4, -7, 2, 7,
    -- layer=1 filter=244 channel=70
    8, 5, -3, 0, -6, 8, 4, -1, -3,
    -- layer=1 filter=244 channel=71
    -9, 6, 0, 5, -11, -3, -3, -10, -11,
    -- layer=1 filter=244 channel=72
    -2, 0, -7, -10, -10, -5, -11, -11, 1,
    -- layer=1 filter=244 channel=73
    -2, -9, -6, -8, 6, 4, 5, -8, -6,
    -- layer=1 filter=244 channel=74
    2, 4, -1, 6, 1, 4, -2, -6, -3,
    -- layer=1 filter=244 channel=75
    0, 1, -7, 7, 3, 6, -9, -2, 2,
    -- layer=1 filter=244 channel=76
    9, -4, 4, -10, 7, 1, -4, -11, -11,
    -- layer=1 filter=244 channel=77
    -10, -2, -1, 1, 4, 8, 5, 5, -3,
    -- layer=1 filter=244 channel=78
    -9, 4, 8, -10, 0, 4, -8, 6, 4,
    -- layer=1 filter=244 channel=79
    2, -7, 9, -6, 5, -5, -9, 9, -6,
    -- layer=1 filter=244 channel=80
    2, -7, -11, -8, 6, 4, -6, -3, 3,
    -- layer=1 filter=244 channel=81
    -2, -9, 3, 6, 8, -6, -2, 7, -10,
    -- layer=1 filter=244 channel=82
    -4, 1, 4, -5, -1, -3, -2, 3, 0,
    -- layer=1 filter=244 channel=83
    7, 1, -8, 0, -5, -10, -8, -1, 1,
    -- layer=1 filter=244 channel=84
    -4, 0, -4, 0, -7, -4, 1, 8, -7,
    -- layer=1 filter=244 channel=85
    -1, 7, -7, -7, -2, 9, -1, -1, -5,
    -- layer=1 filter=244 channel=86
    -1, -2, -2, 0, 5, 0, -2, 4, 3,
    -- layer=1 filter=244 channel=87
    -5, -9, 7, 5, -7, 4, -4, 4, 0,
    -- layer=1 filter=244 channel=88
    2, 2, 0, -2, -12, -8, 7, -4, 7,
    -- layer=1 filter=244 channel=89
    -5, -1, -2, -10, 7, 0, -10, 0, -5,
    -- layer=1 filter=244 channel=90
    4, -3, -1, -10, 1, 8, -1, -6, -1,
    -- layer=1 filter=244 channel=91
    -5, 0, -2, 7, 8, -7, -12, 0, -1,
    -- layer=1 filter=244 channel=92
    -6, -2, -1, 1, 2, -8, 2, -5, -3,
    -- layer=1 filter=244 channel=93
    8, -8, 1, -6, -9, 0, -7, -5, 4,
    -- layer=1 filter=244 channel=94
    -11, -11, -11, 1, -11, 4, 1, 8, -8,
    -- layer=1 filter=244 channel=95
    -4, 0, -5, -1, 0, 5, 1, 0, 3,
    -- layer=1 filter=244 channel=96
    -9, 0, 5, 3, 7, 0, -7, -1, -10,
    -- layer=1 filter=244 channel=97
    -3, 3, 6, 6, 4, -6, 7, 7, 0,
    -- layer=1 filter=244 channel=98
    2, 2, 10, 7, -7, -7, 1, -5, 2,
    -- layer=1 filter=244 channel=99
    2, 7, 2, -3, 0, 0, 3, 7, -5,
    -- layer=1 filter=244 channel=100
    7, 3, 0, -10, -4, -10, 6, -1, 2,
    -- layer=1 filter=244 channel=101
    0, 2, -2, -10, -8, -2, -5, -1, 4,
    -- layer=1 filter=244 channel=102
    0, -10, 3, 7, -3, 6, 8, -3, -5,
    -- layer=1 filter=244 channel=103
    1, -3, 3, -7, -3, -1, 0, 4, -6,
    -- layer=1 filter=244 channel=104
    3, -3, -4, 0, -5, -5, -2, 1, -1,
    -- layer=1 filter=244 channel=105
    7, -5, -10, 6, 3, -6, 5, -5, 2,
    -- layer=1 filter=244 channel=106
    -7, 6, 1, 0, 7, 8, 2, -4, -3,
    -- layer=1 filter=244 channel=107
    -11, -8, -8, 6, -9, 4, 3, 4, -9,
    -- layer=1 filter=244 channel=108
    -9, 1, -7, -5, 3, -5, 6, -1, -7,
    -- layer=1 filter=244 channel=109
    -8, 1, 0, -1, 9, 11, 10, 5, -6,
    -- layer=1 filter=244 channel=110
    5, -1, -10, 8, -10, -8, -5, -3, -7,
    -- layer=1 filter=244 channel=111
    -2, 5, 2, 7, 3, 10, -4, -6, 7,
    -- layer=1 filter=244 channel=112
    0, 7, -6, -6, -2, 0, 0, -7, 0,
    -- layer=1 filter=244 channel=113
    -6, -6, 11, 0, 0, 8, -10, 0, 8,
    -- layer=1 filter=244 channel=114
    1, -4, 8, 6, -3, -8, -11, 0, 0,
    -- layer=1 filter=244 channel=115
    0, -6, -1, 6, -3, -3, 6, -11, -9,
    -- layer=1 filter=244 channel=116
    -9, 1, -6, 2, 4, 4, -9, -5, 9,
    -- layer=1 filter=244 channel=117
    7, -6, -2, 0, 0, -3, 0, -1, 5,
    -- layer=1 filter=244 channel=118
    9, -11, 5, 0, 8, -4, 1, -2, -3,
    -- layer=1 filter=244 channel=119
    0, 4, -6, 5, -11, 11, 0, -2, 2,
    -- layer=1 filter=244 channel=120
    1, 4, -6, 0, 2, 7, 7, -2, -3,
    -- layer=1 filter=244 channel=121
    -2, -7, 0, 9, 3, -10, -3, -5, -4,
    -- layer=1 filter=244 channel=122
    4, -8, -6, -9, 1, 6, 4, 1, -1,
    -- layer=1 filter=244 channel=123
    -8, 7, 7, 1, -6, 6, -2, -3, 4,
    -- layer=1 filter=244 channel=124
    -4, -1, 5, 1, -12, 0, -7, -9, 4,
    -- layer=1 filter=244 channel=125
    -3, 8, 0, 0, -5, -5, -11, 7, 4,
    -- layer=1 filter=244 channel=126
    -7, 6, -1, -11, 4, 0, -1, 6, 6,
    -- layer=1 filter=244 channel=127
    -7, -5, 6, -12, 2, 0, 7, -2, 0,
    -- layer=1 filter=245 channel=0
    0, -21, -26, -2, -13, -19, 4, 18, 17,
    -- layer=1 filter=245 channel=1
    9, 2, 7, -6, -5, 20, -8, 12, -7,
    -- layer=1 filter=245 channel=2
    40, 22, 2, -8, -15, -28, -23, -51, -64,
    -- layer=1 filter=245 channel=3
    10, 8, 13, 0, -14, -3, 4, -11, -3,
    -- layer=1 filter=245 channel=4
    -6, -5, -13, -3, -19, -6, -8, -4, -13,
    -- layer=1 filter=245 channel=5
    8, -3, -10, 28, 31, 21, 30, 21, 19,
    -- layer=1 filter=245 channel=6
    0, 22, 25, 6, 31, 11, -18, -26, -27,
    -- layer=1 filter=245 channel=7
    -59, -9, -12, -25, -4, 1, -14, -4, -6,
    -- layer=1 filter=245 channel=8
    29, 26, 14, 2, -8, -8, 0, 11, -17,
    -- layer=1 filter=245 channel=9
    19, 11, 10, -12, -61, -7, -3, -17, 28,
    -- layer=1 filter=245 channel=10
    -40, -34, -6, -8, 16, -13, 0, 12, -10,
    -- layer=1 filter=245 channel=11
    -27, -51, -35, -12, -32, -35, 13, 3, 10,
    -- layer=1 filter=245 channel=12
    17, 48, 21, -14, 4, -3, -11, -48, -27,
    -- layer=1 filter=245 channel=13
    16, 39, 57, 10, 31, 13, -31, -26, -33,
    -- layer=1 filter=245 channel=14
    -36, -13, -43, -41, -3, -36, -6, 5, -23,
    -- layer=1 filter=245 channel=15
    59, 46, 58, 7, 37, 10, 7, 0, -12,
    -- layer=1 filter=245 channel=16
    14, 11, 22, -8, 1, 3, 5, 3, 13,
    -- layer=1 filter=245 channel=17
    18, 54, 47, 31, 44, 18, -22, -17, -15,
    -- layer=1 filter=245 channel=18
    -34, -25, -10, 0, 9, -18, -4, 1, 12,
    -- layer=1 filter=245 channel=19
    32, 15, 14, -28, 8, 0, 2, -1, 29,
    -- layer=1 filter=245 channel=20
    34, 48, 45, 35, 52, 27, -22, -7, -25,
    -- layer=1 filter=245 channel=21
    -53, -44, -31, -22, -51, -10, -21, -15, -4,
    -- layer=1 filter=245 channel=22
    35, 65, 64, 23, 37, 46, -41, -11, -32,
    -- layer=1 filter=245 channel=23
    -18, 1, -12, -52, -46, -45, 14, 14, 23,
    -- layer=1 filter=245 channel=24
    -54, -74, -52, -32, -53, -38, 22, -1, 46,
    -- layer=1 filter=245 channel=25
    -33, 4, -2, 4, 13, 23, 0, 17, -3,
    -- layer=1 filter=245 channel=26
    35, 53, 44, 17, 12, 26, -18, -7, -21,
    -- layer=1 filter=245 channel=27
    42, 18, 16, 37, 22, 20, 51, 51, 41,
    -- layer=1 filter=245 channel=28
    -33, 4, -1, -55, -15, -12, -48, -14, -5,
    -- layer=1 filter=245 channel=29
    -8, -2, 11, 12, -3, -5, -7, -7, 5,
    -- layer=1 filter=245 channel=30
    -32, -41, -19, -22, 3, -25, -8, 8, 11,
    -- layer=1 filter=245 channel=31
    15, 47, 42, 30, 48, 52, -2, 7, 0,
    -- layer=1 filter=245 channel=32
    -35, -25, -35, 2, -16, -12, 18, -19, 23,
    -- layer=1 filter=245 channel=33
    19, 7, 12, 7, 19, 5, -12, -6, -13,
    -- layer=1 filter=245 channel=34
    -18, 2, -9, 0, 11, -9, -17, -24, -17,
    -- layer=1 filter=245 channel=35
    0, -7, -12, -18, -23, -8, 0, 6, -19,
    -- layer=1 filter=245 channel=36
    -1, -54, -45, -12, -52, -41, 24, 6, 16,
    -- layer=1 filter=245 channel=37
    0, -2, 19, 43, 61, 58, 30, 50, 43,
    -- layer=1 filter=245 channel=38
    17, 27, 22, 10, 30, 13, -15, -12, -19,
    -- layer=1 filter=245 channel=39
    8, -9, -6, -25, -44, -39, 15, 2, 4,
    -- layer=1 filter=245 channel=40
    36, 45, 42, 39, 50, 20, -30, -12, -24,
    -- layer=1 filter=245 channel=41
    -63, -64, -41, -3, -37, 4, 0, -19, 59,
    -- layer=1 filter=245 channel=42
    66, 64, 53, 3, 2, -7, -46, -32, -42,
    -- layer=1 filter=245 channel=43
    -1, 2, -5, -18, -20, -5, -2, 3, -12,
    -- layer=1 filter=245 channel=44
    12, 18, 24, 23, 17, 15, 13, -9, -11,
    -- layer=1 filter=245 channel=45
    -6, -25, -26, 12, 9, -4, 11, -1, 1,
    -- layer=1 filter=245 channel=46
    26, 16, -8, -1, 0, -11, -22, -29, -33,
    -- layer=1 filter=245 channel=47
    -32, -11, 8, -7, 36, 41, 7, 14, 37,
    -- layer=1 filter=245 channel=48
    -46, -34, -16, -21, -34, -33, -36, -40, -36,
    -- layer=1 filter=245 channel=49
    4, 0, 0, 20, 22, 0, -11, -13, -37,
    -- layer=1 filter=245 channel=50
    30, 17, 24, 15, 3, 0, -16, -14, -15,
    -- layer=1 filter=245 channel=51
    -27, -19, 2, -16, 0, -4, -26, -4, -18,
    -- layer=1 filter=245 channel=52
    -10, 19, 8, 17, 15, 9, 2, 2, 16,
    -- layer=1 filter=245 channel=53
    5, -10, 2, 4, -21, 8, 0, -5, 7,
    -- layer=1 filter=245 channel=54
    -38, -25, -16, -2, 36, 30, 8, 28, 27,
    -- layer=1 filter=245 channel=55
    -23, -56, -38, -24, -65, -49, 46, 34, 42,
    -- layer=1 filter=245 channel=56
    0, 0, -8, 5, 5, 0, 3, 5, -3,
    -- layer=1 filter=245 channel=57
    27, 56, 52, 43, 74, 34, 3, 1, -4,
    -- layer=1 filter=245 channel=58
    -23, -9, 2, -43, 14, -7, -5, -8, 19,
    -- layer=1 filter=245 channel=59
    -3, 4, -18, -35, -37, -34, -3, 5, -1,
    -- layer=1 filter=245 channel=60
    -17, -5, -12, -13, -12, -28, -17, -10, -4,
    -- layer=1 filter=245 channel=61
    -3, 0, 8, 1, 4, 1, 9, 5, -12,
    -- layer=1 filter=245 channel=62
    1, 21, 14, -10, 8, -13, 13, 6, 6,
    -- layer=1 filter=245 channel=63
    -49, -64, -38, -16, -34, -34, 42, 17, 35,
    -- layer=1 filter=245 channel=64
    -19, 5, 11, -16, 11, 19, -31, -16, -14,
    -- layer=1 filter=245 channel=65
    -33, -22, -10, -44, -33, -41, -46, -38, -15,
    -- layer=1 filter=245 channel=66
    5, -34, -59, 6, -31, -37, 35, 30, 32,
    -- layer=1 filter=245 channel=67
    -44, -54, -54, -69, -56, -52, -24, -54, -48,
    -- layer=1 filter=245 channel=68
    -16, -23, -31, 17, -17, 3, 16, -27, -5,
    -- layer=1 filter=245 channel=69
    14, 12, 18, -22, 5, -8, 13, -2, -7,
    -- layer=1 filter=245 channel=70
    11, 16, 0, 4, 31, 11, 0, 1, 0,
    -- layer=1 filter=245 channel=71
    -35, -59, -71, -31, -92, -38, 14, 18, 13,
    -- layer=1 filter=245 channel=72
    11, 0, 11, 6, 2, 11, 11, 17, 8,
    -- layer=1 filter=245 channel=73
    -9, -10, -13, 4, -13, -13, 2, -11, 0,
    -- layer=1 filter=245 channel=74
    1, 5, 10, 21, 5, 10, -14, -19, -7,
    -- layer=1 filter=245 channel=75
    -28, -16, -36, -25, -15, -36, 11, -25, -38,
    -- layer=1 filter=245 channel=76
    -32, -33, -15, 0, -13, -12, 13, -37, 17,
    -- layer=1 filter=245 channel=77
    -73, -73, -49, -37, -61, -30, 0, 1, 2,
    -- layer=1 filter=245 channel=78
    10, 10, -3, 23, 49, 15, 14, 23, 3,
    -- layer=1 filter=245 channel=79
    24, 40, 33, 2, 14, -5, -10, -2, -9,
    -- layer=1 filter=245 channel=80
    -10, 0, -13, -22, -4, -18, -16, -12, -12,
    -- layer=1 filter=245 channel=81
    -16, -40, -16, -59, -73, -72, 31, -5, 34,
    -- layer=1 filter=245 channel=82
    -65, -57, -40, -54, -39, -30, -29, -36, -25,
    -- layer=1 filter=245 channel=83
    -18, -25, 18, -21, -13, 0, 16, 3, -27,
    -- layer=1 filter=245 channel=84
    14, 21, 36, 19, 21, 14, 7, -21, -7,
    -- layer=1 filter=245 channel=85
    0, -23, 12, -4, 2, -4, -3, -5, 31,
    -- layer=1 filter=245 channel=86
    43, 18, 19, 20, 32, 6, 9, 4, 9,
    -- layer=1 filter=245 channel=87
    19, 8, 1, -2, 20, 3, 16, 1, 17,
    -- layer=1 filter=245 channel=88
    -29, -30, -35, -16, -17, -22, -23, -23, -20,
    -- layer=1 filter=245 channel=89
    -51, -65, -54, -35, -53, -42, -31, -49, -42,
    -- layer=1 filter=245 channel=90
    -17, -20, 6, 0, -23, -13, 9, -24, -12,
    -- layer=1 filter=245 channel=91
    0, 29, 24, 16, 41, 30, -24, 2, -13,
    -- layer=1 filter=245 channel=92
    -81, -56, -6, -65, -25, -9, 5, -26, 19,
    -- layer=1 filter=245 channel=93
    -64, -74, -56, -40, -72, -46, 0, -1, 14,
    -- layer=1 filter=245 channel=94
    16, 21, 4, 4, 7, -7, 0, 7, -8,
    -- layer=1 filter=245 channel=95
    -34, -6, -1, -4, 0, -12, -3, -20, 2,
    -- layer=1 filter=245 channel=96
    12, -7, 0, 12, 0, 16, -3, -10, 8,
    -- layer=1 filter=245 channel=97
    -4, -16, -11, -24, -41, -22, -2, -3, 0,
    -- layer=1 filter=245 channel=98
    27, 43, 53, 0, 10, -2, -11, -8, -8,
    -- layer=1 filter=245 channel=99
    -31, -41, -29, -49, -25, -30, -32, -12, -37,
    -- layer=1 filter=245 channel=100
    -38, -33, -13, 14, 4, -15, 58, 29, 59,
    -- layer=1 filter=245 channel=101
    -4, 17, 5, 21, 26, 22, -15, -12, -21,
    -- layer=1 filter=245 channel=102
    -11, 10, -3, 5, 13, 9, -19, -7, -4,
    -- layer=1 filter=245 channel=103
    -1, -24, -9, 22, 4, -15, 14, 13, 15,
    -- layer=1 filter=245 channel=104
    -24, 0, 1, -7, 24, 13, 15, -8, 13,
    -- layer=1 filter=245 channel=105
    -13, -42, -43, -26, -46, -48, 5, 1, 3,
    -- layer=1 filter=245 channel=106
    12, 34, 9, 21, 21, 26, -17, -18, -17,
    -- layer=1 filter=245 channel=107
    2, -2, -11, 2, -3, 9, -1, -8, 0,
    -- layer=1 filter=245 channel=108
    1, -12, 1, 9, -14, -24, 20, -10, -16,
    -- layer=1 filter=245 channel=109
    3, -10, 5, -6, 6, -1, -7, 7, 6,
    -- layer=1 filter=245 channel=110
    -22, -7, -23, -7, -14, -7, -16, -10, -23,
    -- layer=1 filter=245 channel=111
    -29, -37, 15, -8, 3, -48, -20, -34, -3,
    -- layer=1 filter=245 channel=112
    -53, -21, -19, 5, -2, -14, 0, -19, 13,
    -- layer=1 filter=245 channel=113
    33, 55, 53, 34, 46, 32, -25, -2, -25,
    -- layer=1 filter=245 channel=114
    -8, -59, -21, -34, -30, -31, 27, 4, -5,
    -- layer=1 filter=245 channel=115
    27, 40, 15, 30, 25, 8, 2, -5, -6,
    -- layer=1 filter=245 channel=116
    7, -4, 6, 11, -11, 9, -9, -4, -2,
    -- layer=1 filter=245 channel=117
    -2, -11, 13, 1, 26, -24, -11, 0, -3,
    -- layer=1 filter=245 channel=118
    -15, -32, 0, -9, -17, -21, -18, -22, -10,
    -- layer=1 filter=245 channel=119
    -40, -79, -57, -17, -43, -28, 15, -30, 7,
    -- layer=1 filter=245 channel=120
    -37, -12, -3, -16, -7, 0, -2, -7, 14,
    -- layer=1 filter=245 channel=121
    -4, -27, -26, -7, -23, -24, 12, 13, 18,
    -- layer=1 filter=245 channel=122
    10, -4, -8, -9, -1, 4, 5, -5, 10,
    -- layer=1 filter=245 channel=123
    -12, -68, -78, 21, -23, -25, 57, 30, 13,
    -- layer=1 filter=245 channel=124
    -20, -18, -20, 2, -8, -8, -2, 7, -7,
    -- layer=1 filter=245 channel=125
    -20, 9, 6, 5, 32, 5, -17, -17, -4,
    -- layer=1 filter=245 channel=126
    -36, 17, 27, -23, -19, 1, -10, 15, -5,
    -- layer=1 filter=245 channel=127
    -17, -24, 6, 0, 7, -13, 1, 7, 24,
    -- layer=1 filter=246 channel=0
    -6, -2, -4, 3, 2, 0, -5, -3, 0,
    -- layer=1 filter=246 channel=1
    -5, -1, 7, -9, 5, 0, 3, -10, 2,
    -- layer=1 filter=246 channel=2
    1, 8, -9, 0, 8, -5, -10, -10, 5,
    -- layer=1 filter=246 channel=3
    0, 5, 11, 1, -5, 1, -10, -3, 6,
    -- layer=1 filter=246 channel=4
    0, 5, -12, -2, 1, -1, -8, -9, -11,
    -- layer=1 filter=246 channel=5
    0, -11, -7, 5, -9, -9, 2, 3, 6,
    -- layer=1 filter=246 channel=6
    -4, -6, -11, 7, -11, -5, 0, -7, 6,
    -- layer=1 filter=246 channel=7
    -5, -2, 6, -4, -2, 0, -4, 7, -1,
    -- layer=1 filter=246 channel=8
    2, 1, -10, -9, 2, 6, -2, 5, 5,
    -- layer=1 filter=246 channel=9
    1, 4, 10, 0, -2, 6, 3, 7, -4,
    -- layer=1 filter=246 channel=10
    2, 0, 7, -8, 7, 2, 3, 7, 7,
    -- layer=1 filter=246 channel=11
    -6, -3, -5, -1, -11, -10, -9, 1, 5,
    -- layer=1 filter=246 channel=12
    5, -9, -4, 10, -7, -5, -7, 10, -8,
    -- layer=1 filter=246 channel=13
    8, -7, 7, 2, 1, 0, 2, -8, -2,
    -- layer=1 filter=246 channel=14
    -7, 0, 9, -3, -11, 1, 1, 0, -8,
    -- layer=1 filter=246 channel=15
    0, -1, 0, 3, -9, -3, 6, 0, -12,
    -- layer=1 filter=246 channel=16
    -11, 0, 2, 5, -4, -7, -6, 3, 2,
    -- layer=1 filter=246 channel=17
    -10, -8, -12, 0, -7, 2, -5, -2, 3,
    -- layer=1 filter=246 channel=18
    -7, -11, 6, 7, -12, 4, 2, -5, -8,
    -- layer=1 filter=246 channel=19
    -8, -3, -12, -9, -4, 6, 8, -5, -9,
    -- layer=1 filter=246 channel=20
    -9, -11, -7, -6, 2, 6, 6, 4, -7,
    -- layer=1 filter=246 channel=21
    8, 1, -8, 8, -10, -8, -6, 0, -5,
    -- layer=1 filter=246 channel=22
    -10, -3, 7, 0, -1, -8, -11, -5, 1,
    -- layer=1 filter=246 channel=23
    -12, -6, -7, 3, 0, 6, -10, 3, 0,
    -- layer=1 filter=246 channel=24
    -1, 1, -11, 4, -3, -5, -8, -9, 7,
    -- layer=1 filter=246 channel=25
    -6, -12, -10, 3, 0, -10, 7, -2, -3,
    -- layer=1 filter=246 channel=26
    -4, 2, 5, 0, -3, 6, -6, 3, -13,
    -- layer=1 filter=246 channel=27
    -7, -5, -9, -3, -1, 2, -10, -8, -6,
    -- layer=1 filter=246 channel=28
    -7, -1, -11, 4, -5, 2, 2, -12, 2,
    -- layer=1 filter=246 channel=29
    3, 8, -2, 5, 3, 2, 0, -11, -6,
    -- layer=1 filter=246 channel=30
    3, -4, 0, 3, -7, -1, -2, -10, -8,
    -- layer=1 filter=246 channel=31
    -6, 6, 6, -4, 2, 3, -11, 5, -10,
    -- layer=1 filter=246 channel=32
    -6, 1, 1, -2, -8, -15, 3, -4, -1,
    -- layer=1 filter=246 channel=33
    5, -9, -7, 0, 10, 0, 7, 4, -4,
    -- layer=1 filter=246 channel=34
    -2, -8, -6, -2, -2, 6, 2, 0, -7,
    -- layer=1 filter=246 channel=35
    -5, -8, 1, 3, 4, 4, -9, 2, -12,
    -- layer=1 filter=246 channel=36
    -1, -3, -5, 5, -7, 0, -3, -5, 8,
    -- layer=1 filter=246 channel=37
    -12, -15, 5, -6, 6, -4, 7, -4, -8,
    -- layer=1 filter=246 channel=38
    3, -3, -3, 3, 0, 8, -10, -7, -4,
    -- layer=1 filter=246 channel=39
    -5, 0, -1, -11, 1, 3, 8, 8, 6,
    -- layer=1 filter=246 channel=40
    -1, 4, 8, -8, 0, 8, 1, -14, -2,
    -- layer=1 filter=246 channel=41
    -5, -12, -10, 2, 2, 3, -6, 4, 2,
    -- layer=1 filter=246 channel=42
    -3, 4, -9, 2, -4, -9, 0, -6, 8,
    -- layer=1 filter=246 channel=43
    4, 4, 3, 5, -3, 0, -6, -8, -9,
    -- layer=1 filter=246 channel=44
    -11, -12, -5, 3, 4, -3, -6, 0, 3,
    -- layer=1 filter=246 channel=45
    3, 5, -5, 0, 0, -7, -2, 8, -7,
    -- layer=1 filter=246 channel=46
    -9, -9, 5, 5, 8, -6, 2, 7, 4,
    -- layer=1 filter=246 channel=47
    -3, 1, 0, -3, -5, -15, 2, 8, -3,
    -- layer=1 filter=246 channel=48
    -2, 3, -8, 6, 4, -10, -2, 4, -6,
    -- layer=1 filter=246 channel=49
    -3, -8, 8, -10, -3, 5, -11, 0, -1,
    -- layer=1 filter=246 channel=50
    -5, 3, -1, -2, 0, -12, 8, 0, 8,
    -- layer=1 filter=246 channel=51
    -5, 9, 9, 3, -11, -1, -9, -6, -5,
    -- layer=1 filter=246 channel=52
    -4, 0, 6, 6, 3, 8, 1, -1, 0,
    -- layer=1 filter=246 channel=53
    -12, 7, -3, -3, 0, -2, -4, 7, -4,
    -- layer=1 filter=246 channel=54
    -4, -9, 2, -8, -7, 7, -4, -11, 6,
    -- layer=1 filter=246 channel=55
    3, -6, 5, 14, 7, -4, -1, 1, -5,
    -- layer=1 filter=246 channel=56
    0, -6, 1, 3, -11, 1, -2, -5, -7,
    -- layer=1 filter=246 channel=57
    5, 2, 2, 3, -1, -6, -2, 5, -7,
    -- layer=1 filter=246 channel=58
    -9, -3, 8, 8, 2, 3, 8, -2, 0,
    -- layer=1 filter=246 channel=59
    3, 4, -1, 4, 0, 3, -10, -8, -1,
    -- layer=1 filter=246 channel=60
    10, -7, -6, -5, 5, -4, -3, 7, -5,
    -- layer=1 filter=246 channel=61
    -8, 3, 7, 6, -5, -2, 5, -3, -4,
    -- layer=1 filter=246 channel=62
    -11, -13, 2, 3, -7, -13, -10, -10, 13,
    -- layer=1 filter=246 channel=63
    4, -10, -4, 2, 3, -9, 4, -7, -4,
    -- layer=1 filter=246 channel=64
    3, -11, 1, 7, 6, 8, -2, 7, -10,
    -- layer=1 filter=246 channel=65
    -1, -11, 7, -8, -11, -11, -10, -6, 7,
    -- layer=1 filter=246 channel=66
    0, 2, 6, 2, 6, -1, 4, -12, -7,
    -- layer=1 filter=246 channel=67
    6, 6, 6, -7, -11, -2, 2, -3, 7,
    -- layer=1 filter=246 channel=68
    0, 5, -8, -7, 3, 0, -2, 3, -9,
    -- layer=1 filter=246 channel=69
    -15, -5, 9, 7, 0, -10, 4, 4, 9,
    -- layer=1 filter=246 channel=70
    -7, -8, -7, 0, -5, -5, -1, 4, 7,
    -- layer=1 filter=246 channel=71
    -1, -8, 5, -7, 0, -8, 8, -3, -6,
    -- layer=1 filter=246 channel=72
    0, 6, 8, 7, -4, 2, 1, 4, 4,
    -- layer=1 filter=246 channel=73
    7, -8, 7, 0, 6, -2, -11, 2, 0,
    -- layer=1 filter=246 channel=74
    6, 6, 5, -7, 1, 4, -6, -9, -4,
    -- layer=1 filter=246 channel=75
    0, -1, -2, 8, -6, -1, -7, -9, -10,
    -- layer=1 filter=246 channel=76
    0, 5, -11, 0, 7, 0, -10, 5, 3,
    -- layer=1 filter=246 channel=77
    -5, 3, -3, -1, 9, -9, 6, 0, -1,
    -- layer=1 filter=246 channel=78
    6, 2, -5, -1, 2, 5, 2, 8, 5,
    -- layer=1 filter=246 channel=79
    0, 2, -1, -7, -4, 1, 7, 1, -1,
    -- layer=1 filter=246 channel=80
    -6, -11, -6, 2, -8, -5, 3, -3, -3,
    -- layer=1 filter=246 channel=81
    0, 5, -11, 4, -10, -5, -9, 4, -7,
    -- layer=1 filter=246 channel=82
    0, 2, 4, -10, -4, -10, -2, -9, -10,
    -- layer=1 filter=246 channel=83
    7, 3, 2, 1, -4, -13, -11, -10, -1,
    -- layer=1 filter=246 channel=84
    0, 1, 2, -1, 4, -1, -8, 7, 0,
    -- layer=1 filter=246 channel=85
    -12, 2, 6, 8, -6, 1, 2, -1, 5,
    -- layer=1 filter=246 channel=86
    -3, -1, -13, -4, -1, 5, -2, 0, 6,
    -- layer=1 filter=246 channel=87
    -6, -9, -2, -7, -6, -5, -11, 0, 8,
    -- layer=1 filter=246 channel=88
    5, -4, -2, 7, -8, 1, 7, -2, -3,
    -- layer=1 filter=246 channel=89
    -10, -6, 7, 0, 8, -6, -1, -11, 4,
    -- layer=1 filter=246 channel=90
    0, 3, -5, -6, 0, 6, 6, -5, -6,
    -- layer=1 filter=246 channel=91
    -9, -11, 9, -2, 4, -12, 5, 2, -4,
    -- layer=1 filter=246 channel=92
    4, -6, 2, -9, 2, -9, -4, 1, -6,
    -- layer=1 filter=246 channel=93
    0, 5, -11, -5, -2, 6, 1, -10, 2,
    -- layer=1 filter=246 channel=94
    -3, 0, -8, 5, -13, -9, -7, -1, 3,
    -- layer=1 filter=246 channel=95
    -6, 6, -4, 5, 6, 7, 6, -3, -3,
    -- layer=1 filter=246 channel=96
    -4, -1, -6, 0, 1, -11, 4, -1, -4,
    -- layer=1 filter=246 channel=97
    2, -1, 2, 0, 0, -4, 5, 7, -5,
    -- layer=1 filter=246 channel=98
    5, -12, 8, -10, 8, 4, -5, -9, 0,
    -- layer=1 filter=246 channel=99
    -7, 6, 1, -11, -9, 0, -11, 2, -6,
    -- layer=1 filter=246 channel=100
    -11, -3, -9, -7, 3, 6, -8, -7, 4,
    -- layer=1 filter=246 channel=101
    0, 6, -4, -10, -9, 5, 0, 2, -3,
    -- layer=1 filter=246 channel=102
    1, -12, -2, 1, -6, -5, 6, -3, 6,
    -- layer=1 filter=246 channel=103
    -9, -3, 7, -6, -11, 5, 7, 8, -7,
    -- layer=1 filter=246 channel=104
    -12, 3, 6, -5, 5, -9, -12, 0, -1,
    -- layer=1 filter=246 channel=105
    -9, 5, -12, 5, -1, -11, -9, 6, -9,
    -- layer=1 filter=246 channel=106
    -3, -11, -5, 3, -6, 2, 9, -6, -6,
    -- layer=1 filter=246 channel=107
    -4, -8, 4, -8, -11, -3, 0, 5, -10,
    -- layer=1 filter=246 channel=108
    -9, -13, -5, 14, -10, -8, 7, 4, -9,
    -- layer=1 filter=246 channel=109
    -5, -2, -8, 7, -2, -6, 6, -3, -9,
    -- layer=1 filter=246 channel=110
    -3, 1, 4, -2, 2, 8, -8, 0, -4,
    -- layer=1 filter=246 channel=111
    -12, 1, 1, 1, -13, -8, -9, -13, -4,
    -- layer=1 filter=246 channel=112
    3, 2, -7, -7, -3, 5, -9, 0, -2,
    -- layer=1 filter=246 channel=113
    -8, 8, -3, 1, -9, -10, -2, 0, -9,
    -- layer=1 filter=246 channel=114
    -4, -13, -10, 1, -3, 1, -2, -3, 0,
    -- layer=1 filter=246 channel=115
    -11, 0, 0, -2, -3, -10, 5, 0, -4,
    -- layer=1 filter=246 channel=116
    8, 1, 5, -7, 1, -2, 9, -8, -5,
    -- layer=1 filter=246 channel=117
    7, -2, -7, -8, 0, -10, -8, -4, -6,
    -- layer=1 filter=246 channel=118
    0, -7, 0, 4, -7, -4, 7, -12, -5,
    -- layer=1 filter=246 channel=119
    -2, -4, 4, 6, -7, 5, -9, -4, -7,
    -- layer=1 filter=246 channel=120
    7, 5, -1, 2, -1, 6, 8, -10, -6,
    -- layer=1 filter=246 channel=121
    5, 0, 9, -6, 9, -6, 7, -1, 4,
    -- layer=1 filter=246 channel=122
    -8, 0, 4, 0, 8, 2, 3, 3, -1,
    -- layer=1 filter=246 channel=123
    -8, -3, 5, 6, -7, 2, -4, 5, 0,
    -- layer=1 filter=246 channel=124
    -8, -12, -9, 6, -11, 8, 1, -5, -1,
    -- layer=1 filter=246 channel=125
    -1, 3, 4, 2, 5, -9, 0, 8, 4,
    -- layer=1 filter=246 channel=126
    1, -14, -11, 6, -4, 0, 2, -6, -10,
    -- layer=1 filter=246 channel=127
    0, 0, -9, -1, -13, -3, 0, -3, -11,
    -- layer=1 filter=247 channel=0
    6, -1, -11, -9, -6, -1, -12, -6, 6,
    -- layer=1 filter=247 channel=1
    -8, -12, 0, -10, 8, 6, 0, 6, -8,
    -- layer=1 filter=247 channel=2
    -10, -12, 1, -2, -2, -6, 5, -8, 6,
    -- layer=1 filter=247 channel=3
    5, 0, 8, 2, -7, 9, 9, -8, 3,
    -- layer=1 filter=247 channel=4
    0, -2, -12, 3, -6, -5, 0, 0, -7,
    -- layer=1 filter=247 channel=5
    3, -3, -1, -5, 0, 6, -5, 7, 2,
    -- layer=1 filter=247 channel=6
    -2, -2, -7, -8, 3, -8, 6, -13, 0,
    -- layer=1 filter=247 channel=7
    -1, 2, -6, -4, 7, -10, 10, -5, -3,
    -- layer=1 filter=247 channel=8
    -1, -1, 5, -6, 3, 6, 8, -9, 8,
    -- layer=1 filter=247 channel=9
    -7, -4, -8, -11, -10, -2, 0, -3, -1,
    -- layer=1 filter=247 channel=10
    -4, 12, 4, -8, -7, -11, -3, -8, -12,
    -- layer=1 filter=247 channel=11
    -2, -11, 4, -3, -5, 3, -3, -11, -5,
    -- layer=1 filter=247 channel=12
    -10, -11, 0, -10, 0, 7, 2, 7, -2,
    -- layer=1 filter=247 channel=13
    -11, 8, -2, -5, -7, -1, 4, 5, 7,
    -- layer=1 filter=247 channel=14
    -7, 0, -8, -4, 5, -7, 0, -9, 4,
    -- layer=1 filter=247 channel=15
    -6, -2, 2, 4, 0, 3, 2, 7, 6,
    -- layer=1 filter=247 channel=16
    3, -10, -2, -7, 5, -9, -6, 9, -9,
    -- layer=1 filter=247 channel=17
    3, 3, 4, -5, 6, 5, -5, -11, -12,
    -- layer=1 filter=247 channel=18
    0, -7, -1, 1, -11, -2, -8, 4, 5,
    -- layer=1 filter=247 channel=19
    -3, -8, 3, 0, 2, -5, -11, 2, 1,
    -- layer=1 filter=247 channel=20
    -1, -10, -2, -12, 7, -12, -2, -10, 0,
    -- layer=1 filter=247 channel=21
    4, -6, 0, 0, -1, 5, -3, 0, -9,
    -- layer=1 filter=247 channel=22
    -11, -8, 5, 2, -10, 0, 6, -4, 5,
    -- layer=1 filter=247 channel=23
    4, -5, 0, 1, -4, 0, -11, -1, -8,
    -- layer=1 filter=247 channel=24
    3, -2, -7, 0, 7, 7, -7, -7, -6,
    -- layer=1 filter=247 channel=25
    -2, -1, 0, -11, 2, 1, -3, 0, -1,
    -- layer=1 filter=247 channel=26
    -7, 4, -11, -14, 0, -10, 7, -2, -6,
    -- layer=1 filter=247 channel=27
    -3, -8, 1, 2, -7, 4, 6, 5, -10,
    -- layer=1 filter=247 channel=28
    1, -2, -4, 3, -8, 0, -6, -1, -10,
    -- layer=1 filter=247 channel=29
    -4, -12, -2, 6, -1, -4, 0, -9, -5,
    -- layer=1 filter=247 channel=30
    -2, 7, 2, 0, -4, -2, 2, -14, 3,
    -- layer=1 filter=247 channel=31
    -1, 3, -15, -9, 0, -1, 6, -4, -10,
    -- layer=1 filter=247 channel=32
    4, -3, 1, 0, 5, -3, 5, -6, 6,
    -- layer=1 filter=247 channel=33
    3, 8, 0, -6, -6, 7, 0, 9, 6,
    -- layer=1 filter=247 channel=34
    7, -3, -8, 5, -5, 4, 0, 3, -4,
    -- layer=1 filter=247 channel=35
    -2, -4, -7, -6, 0, -7, -9, -3, -7,
    -- layer=1 filter=247 channel=36
    -2, 3, -10, 3, -1, -3, 1, -3, 3,
    -- layer=1 filter=247 channel=37
    7, 1, -9, 3, -13, -14, -12, -7, -1,
    -- layer=1 filter=247 channel=38
    -6, -8, 2, -2, -9, 0, -11, 5, 0,
    -- layer=1 filter=247 channel=39
    -12, -3, -6, -11, -3, -10, -8, 5, 6,
    -- layer=1 filter=247 channel=40
    -4, 3, -3, -12, 0, -2, 0, 6, 3,
    -- layer=1 filter=247 channel=41
    -4, -4, -5, -8, 3, -11, 8, -10, -4,
    -- layer=1 filter=247 channel=42
    8, 2, 6, 9, -4, -6, 9, -3, -10,
    -- layer=1 filter=247 channel=43
    -5, -7, -11, 5, 2, 1, 0, -9, -6,
    -- layer=1 filter=247 channel=44
    -2, -10, -1, -5, -4, 5, 0, 3, 0,
    -- layer=1 filter=247 channel=45
    4, -1, -6, 2, -1, 8, -7, 6, 1,
    -- layer=1 filter=247 channel=46
    -5, -10, 3, 2, -4, -2, 8, 9, -7,
    -- layer=1 filter=247 channel=47
    -6, 5, -1, -4, -2, -11, -7, -2, -11,
    -- layer=1 filter=247 channel=48
    6, 9, -3, -4, -9, 3, -3, -7, 7,
    -- layer=1 filter=247 channel=49
    0, -6, 3, -4, 6, -11, -10, 4, 0,
    -- layer=1 filter=247 channel=50
    -7, 0, 1, -8, -11, -3, 0, 8, -7,
    -- layer=1 filter=247 channel=51
    -4, -1, 5, -4, -10, -11, -10, -1, 8,
    -- layer=1 filter=247 channel=52
    -5, -9, -3, -8, 9, 0, -2, 6, 4,
    -- layer=1 filter=247 channel=53
    8, 7, -4, 7, 6, 4, -3, 7, -11,
    -- layer=1 filter=247 channel=54
    -3, 0, 0, 4, 7, 0, 2, 4, 5,
    -- layer=1 filter=247 channel=55
    2, -11, -5, -12, -3, 1, 4, -3, 3,
    -- layer=1 filter=247 channel=56
    -1, 1, -4, 5, 8, 4, -12, 0, 1,
    -- layer=1 filter=247 channel=57
    -1, 4, 4, -4, -6, 3, 5, -2, -7,
    -- layer=1 filter=247 channel=58
    -6, 9, -4, -3, -2, -6, -3, -6, 0,
    -- layer=1 filter=247 channel=59
    8, -12, -10, -10, 8, 0, -1, 1, 3,
    -- layer=1 filter=247 channel=60
    -8, 1, 8, -9, 8, -2, -8, 11, 10,
    -- layer=1 filter=247 channel=61
    0, 9, -8, -9, 7, -9, 4, -4, -9,
    -- layer=1 filter=247 channel=62
    -5, 0, 3, 6, 0, 4, -17, 0, -7,
    -- layer=1 filter=247 channel=63
    -1, -9, -2, 0, -13, 6, 0, -9, -1,
    -- layer=1 filter=247 channel=64
    -2, 1, -7, -12, 0, 5, -1, -6, 9,
    -- layer=1 filter=247 channel=65
    -7, -12, 4, 0, -2, 7, 4, -9, -2,
    -- layer=1 filter=247 channel=66
    -4, 5, 2, -1, -7, 6, -5, -1, -1,
    -- layer=1 filter=247 channel=67
    -2, 8, -2, -6, 5, -4, -9, -11, -14,
    -- layer=1 filter=247 channel=68
    1, -9, -8, -6, 7, 3, 5, 7, -1,
    -- layer=1 filter=247 channel=69
    4, -6, 2, -12, 1, -9, 0, 1, 6,
    -- layer=1 filter=247 channel=70
    4, 0, -5, -11, -1, -9, -9, -4, -9,
    -- layer=1 filter=247 channel=71
    -11, -4, 3, -1, -6, 0, -9, -3, 8,
    -- layer=1 filter=247 channel=72
    2, 7, 5, -2, 5, -3, 3, -9, -2,
    -- layer=1 filter=247 channel=73
    2, -11, -6, -11, 7, -8, 8, 6, -4,
    -- layer=1 filter=247 channel=74
    3, -7, 2, 7, -4, 4, 7, 0, 3,
    -- layer=1 filter=247 channel=75
    0, -2, -12, -10, -14, 1, -5, 4, -13,
    -- layer=1 filter=247 channel=76
    0, 0, -4, 3, -11, 5, -10, 1, -9,
    -- layer=1 filter=247 channel=77
    2, 5, -11, 0, 3, -4, 0, -4, -8,
    -- layer=1 filter=247 channel=78
    0, -2, -8, -6, 5, -5, -12, 5, -3,
    -- layer=1 filter=247 channel=79
    -3, -10, 0, -8, -5, 0, -11, -3, -9,
    -- layer=1 filter=247 channel=80
    0, 3, 1, 5, -1, 3, -5, -5, 6,
    -- layer=1 filter=247 channel=81
    -5, 4, -12, 7, 1, 5, 1, 5, 3,
    -- layer=1 filter=247 channel=82
    -6, 6, -8, 8, -3, -3, -6, -3, 8,
    -- layer=1 filter=247 channel=83
    3, -1, -5, -7, 5, 3, 0, 2, 7,
    -- layer=1 filter=247 channel=84
    8, -9, -3, 6, -10, 2, -3, 0, 5,
    -- layer=1 filter=247 channel=85
    -11, 4, -1, 4, 4, 0, 7, 7, -10,
    -- layer=1 filter=247 channel=86
    3, 0, 4, -7, -8, -8, -9, -10, -3,
    -- layer=1 filter=247 channel=87
    -12, 8, 5, 2, -1, 7, 5, -1, -11,
    -- layer=1 filter=247 channel=88
    -8, -8, 3, 3, -5, -12, 0, 0, -4,
    -- layer=1 filter=247 channel=89
    -8, -5, -1, 6, -2, 7, -2, -2, 0,
    -- layer=1 filter=247 channel=90
    7, -11, -7, -11, -5, -7, -10, -2, -6,
    -- layer=1 filter=247 channel=91
    6, -4, 6, -6, 7, -6, -8, -3, 7,
    -- layer=1 filter=247 channel=92
    3, 1, 0, 6, -6, -12, -6, -5, 0,
    -- layer=1 filter=247 channel=93
    -3, 5, 1, -5, 4, 0, 0, -3, 1,
    -- layer=1 filter=247 channel=94
    -9, 7, 7, -5, 1, -10, -9, -6, 2,
    -- layer=1 filter=247 channel=95
    5, 1, -12, 2, 2, -4, 5, 1, 5,
    -- layer=1 filter=247 channel=96
    4, 8, 0, 0, -7, 1, -4, 1, -10,
    -- layer=1 filter=247 channel=97
    0, -3, -1, 5, 4, -12, 2, 2, 4,
    -- layer=1 filter=247 channel=98
    2, -10, 2, -10, 4, -5, -1, 0, -2,
    -- layer=1 filter=247 channel=99
    -7, 5, 2, -6, -5, 6, 1, -1, 0,
    -- layer=1 filter=247 channel=100
    3, -4, 7, 4, -4, -9, 7, -4, -1,
    -- layer=1 filter=247 channel=101
    -11, 0, 3, 0, 0, 6, 5, -10, 8,
    -- layer=1 filter=247 channel=102
    -7, -7, -7, 7, -1, 6, -12, -3, 6,
    -- layer=1 filter=247 channel=103
    2, -3, 0, 1, 7, -3, 5, 3, -9,
    -- layer=1 filter=247 channel=104
    -12, 0, -6, 6, -4, -4, 3, -6, -9,
    -- layer=1 filter=247 channel=105
    0, -8, 3, 0, 0, -6, -8, -3, -7,
    -- layer=1 filter=247 channel=106
    -7, -3, -7, -9, 5, 5, 0, 4, 1,
    -- layer=1 filter=247 channel=107
    4, 9, 9, 6, 5, 4, -5, -3, 7,
    -- layer=1 filter=247 channel=108
    -6, 4, 11, -15, -6, 3, 4, -7, -6,
    -- layer=1 filter=247 channel=109
    -5, -11, 6, 9, 8, 7, 1, 9, -8,
    -- layer=1 filter=247 channel=110
    -1, 6, 5, -8, 0, -9, -7, -3, 7,
    -- layer=1 filter=247 channel=111
    -1, -5, 0, -3, 0, -12, 2, 2, 0,
    -- layer=1 filter=247 channel=112
    4, 3, -4, -7, 7, 6, 8, 4, 0,
    -- layer=1 filter=247 channel=113
    0, 9, -7, -4, -6, -9, 0, 0, -2,
    -- layer=1 filter=247 channel=114
    4, 1, 0, -6, 2, -16, -5, -15, 3,
    -- layer=1 filter=247 channel=115
    -10, -7, 4, 2, 3, -4, -7, 0, -6,
    -- layer=1 filter=247 channel=116
    -7, 5, -6, -5, -7, 0, 10, -2, -3,
    -- layer=1 filter=247 channel=117
    1, 7, 0, -3, 6, 2, 2, 0, -1,
    -- layer=1 filter=247 channel=118
    7, 2, 0, 0, -4, -2, 0, -1, -2,
    -- layer=1 filter=247 channel=119
    -9, -11, 0, -8, -6, 9, 8, 6, 4,
    -- layer=1 filter=247 channel=120
    0, 8, -11, -2, -3, -3, 6, 6, -8,
    -- layer=1 filter=247 channel=121
    0, -7, -2, -5, 4, -8, -13, -6, 0,
    -- layer=1 filter=247 channel=122
    -4, 8, 7, -6, 1, 4, -8, 3, 0,
    -- layer=1 filter=247 channel=123
    -8, 4, 0, 0, -9, -10, 4, 3, 0,
    -- layer=1 filter=247 channel=124
    0, -2, 5, -6, 4, 6, 1, 4, -3,
    -- layer=1 filter=247 channel=125
    -3, -1, -3, -15, 9, 3, 8, -6, 1,
    -- layer=1 filter=247 channel=126
    -9, 7, -10, -1, -11, 7, 3, -7, 7,
    -- layer=1 filter=247 channel=127
    4, 3, 1, 0, -3, -12, -10, -4, -11,
    -- layer=1 filter=248 channel=0
    -3, 3, 3, -9, -5, 2, 7, -9, 0,
    -- layer=1 filter=248 channel=1
    -2, -6, 0, -2, -2, 4, 8, -6, -1,
    -- layer=1 filter=248 channel=2
    -10, -16, 5, -1, -12, -4, -8, -7, 7,
    -- layer=1 filter=248 channel=3
    -1, -3, 4, -3, 2, 8, 1, -4, -8,
    -- layer=1 filter=248 channel=4
    -5, -1, -3, 8, -4, -5, -4, -2, -2,
    -- layer=1 filter=248 channel=5
    -8, 0, -4, -15, -6, -7, 3, -4, -16,
    -- layer=1 filter=248 channel=6
    -4, -5, 8, 6, -8, 4, -6, 10, -2,
    -- layer=1 filter=248 channel=7
    8, -10, -2, 0, -16, 1, 2, 0, 1,
    -- layer=1 filter=248 channel=8
    6, 1, -9, -10, -3, 0, 4, -10, 7,
    -- layer=1 filter=248 channel=9
    -3, -6, 3, 5, -4, 0, -3, 11, 6,
    -- layer=1 filter=248 channel=10
    -5, -7, 4, -1, -7, -8, -2, -6, -19,
    -- layer=1 filter=248 channel=11
    1, -6, -1, 0, 2, 3, -8, 7, -4,
    -- layer=1 filter=248 channel=12
    -3, -5, -4, -6, -2, 3, -8, 3, 0,
    -- layer=1 filter=248 channel=13
    -2, -8, 0, -5, 0, 1, 5, -1, -6,
    -- layer=1 filter=248 channel=14
    -1, -3, -14, -2, -13, -6, -12, -4, -11,
    -- layer=1 filter=248 channel=15
    -6, 0, -3, -14, -1, 7, -11, 5, -2,
    -- layer=1 filter=248 channel=16
    -9, -7, 9, 1, 0, 0, 2, -12, -10,
    -- layer=1 filter=248 channel=17
    4, -6, 2, 0, -3, 8, 8, 1, -5,
    -- layer=1 filter=248 channel=18
    -11, -1, -3, 3, -8, -3, -14, -15, 10,
    -- layer=1 filter=248 channel=19
    -2, -5, 8, -5, -1, -5, -3, -11, -7,
    -- layer=1 filter=248 channel=20
    8, -10, -9, -12, -10, 3, 0, -8, -6,
    -- layer=1 filter=248 channel=21
    -6, -8, -7, -9, -15, 0, 4, 6, 3,
    -- layer=1 filter=248 channel=22
    -8, -7, 0, -3, -3, 3, 0, -4, 2,
    -- layer=1 filter=248 channel=23
    1, 6, -9, -1, 2, -10, -5, -5, -12,
    -- layer=1 filter=248 channel=24
    -12, -11, 0, -3, -11, -1, 6, 7, -4,
    -- layer=1 filter=248 channel=25
    -11, -5, 7, 3, -3, -12, 3, -1, 0,
    -- layer=1 filter=248 channel=26
    1, -3, -10, 0, -8, 1, 0, 1, 0,
    -- layer=1 filter=248 channel=27
    -13, -19, -21, -11, -9, -9, -4, -5, 6,
    -- layer=1 filter=248 channel=28
    0, 0, -4, 1, 4, -11, -3, -11, 1,
    -- layer=1 filter=248 channel=29
    -1, -6, 0, 5, 2, -2, 7, -6, -2,
    -- layer=1 filter=248 channel=30
    -12, -5, 2, 4, 0, -7, 0, -19, -7,
    -- layer=1 filter=248 channel=31
    -13, -7, -9, 6, 1, 1, -5, -12, 2,
    -- layer=1 filter=248 channel=32
    -12, -2, -5, -6, 2, 4, -3, 0, 2,
    -- layer=1 filter=248 channel=33
    -2, -2, -5, 5, 5, 2, 0, -1, -1,
    -- layer=1 filter=248 channel=34
    1, 8, 3, 8, 6, 5, 2, -11, 5,
    -- layer=1 filter=248 channel=35
    -5, 0, 5, -9, 7, -4, -3, -8, -1,
    -- layer=1 filter=248 channel=36
    6, 6, -2, -5, -5, -10, 2, 3, 1,
    -- layer=1 filter=248 channel=37
    -4, 2, -11, 4, 1, 6, 4, -13, 1,
    -- layer=1 filter=248 channel=38
    -11, 5, -6, -1, -2, 8, 5, 10, 2,
    -- layer=1 filter=248 channel=39
    -9, 0, 3, -5, 3, -10, 2, 4, 6,
    -- layer=1 filter=248 channel=40
    3, -10, 10, -5, -1, 5, 4, -8, -6,
    -- layer=1 filter=248 channel=41
    -4, 8, -9, 4, 1, 0, 0, -3, 0,
    -- layer=1 filter=248 channel=42
    -1, -8, 0, 0, -1, -5, 3, 5, 9,
    -- layer=1 filter=248 channel=43
    -1, 4, 0, -9, 1, 0, 8, 1, 3,
    -- layer=1 filter=248 channel=44
    0, -3, -3, -7, -10, -5, 1, -9, 2,
    -- layer=1 filter=248 channel=45
    -13, 2, 6, -8, -13, -10, -6, -12, -5,
    -- layer=1 filter=248 channel=46
    1, 0, -4, 8, 10, 0, 0, -5, -7,
    -- layer=1 filter=248 channel=47
    3, -3, 3, -2, -1, -5, -8, -9, 0,
    -- layer=1 filter=248 channel=48
    8, 0, 5, 8, -3, -2, -11, -2, -5,
    -- layer=1 filter=248 channel=49
    3, -7, 8, -11, 4, -7, -6, -9, 7,
    -- layer=1 filter=248 channel=50
    -3, 0, 0, -4, -9, -3, 0, 0, 7,
    -- layer=1 filter=248 channel=51
    -7, -8, -6, -6, 1, -3, -2, -3, 0,
    -- layer=1 filter=248 channel=52
    9, 8, -11, 9, 3, -12, 5, -6, 8,
    -- layer=1 filter=248 channel=53
    1, 6, 0, 1, -6, 0, -3, 7, -9,
    -- layer=1 filter=248 channel=54
    -7, 3, 1, -6, 1, -8, -8, 0, -12,
    -- layer=1 filter=248 channel=55
    -6, -15, -7, -13, 0, -11, -6, 0, -6,
    -- layer=1 filter=248 channel=56
    -11, 0, -3, 3, 0, 3, -1, 0, -4,
    -- layer=1 filter=248 channel=57
    2, -1, -10, -3, -1, 2, 4, 1, 0,
    -- layer=1 filter=248 channel=58
    3, -14, 1, -8, 5, -4, 0, -3, 1,
    -- layer=1 filter=248 channel=59
    2, 1, -10, 4, -8, -6, 6, -4, 1,
    -- layer=1 filter=248 channel=60
    -8, -6, -10, 6, 1, -7, -4, -6, 2,
    -- layer=1 filter=248 channel=61
    -2, -3, 8, 6, -6, 2, -10, 4, 7,
    -- layer=1 filter=248 channel=62
    -4, -6, 4, 2, 8, 0, 3, -13, -11,
    -- layer=1 filter=248 channel=63
    -7, 5, 0, 4, -1, 3, 8, -9, 1,
    -- layer=1 filter=248 channel=64
    -6, 4, 0, 6, -9, 7, 6, -3, -6,
    -- layer=1 filter=248 channel=65
    8, -2, -11, -2, 6, -1, 6, 3, -10,
    -- layer=1 filter=248 channel=66
    6, -11, -2, -11, 0, -1, -11, 7, 0,
    -- layer=1 filter=248 channel=67
    7, -5, -5, -5, -4, -2, 1, 1, 4,
    -- layer=1 filter=248 channel=68
    -9, -2, -7, -12, -2, -12, -11, 11, 4,
    -- layer=1 filter=248 channel=69
    0, -12, 3, -11, 2, 6, -5, -6, 0,
    -- layer=1 filter=248 channel=70
    1, -13, -8, -3, 5, 4, -1, -8, 7,
    -- layer=1 filter=248 channel=71
    -2, 1, -2, -4, 2, 3, 0, -4, -9,
    -- layer=1 filter=248 channel=72
    1, 0, 6, -10, -7, 8, 3, -5, -2,
    -- layer=1 filter=248 channel=73
    7, -3, 3, 7, 4, -1, -4, 1, 3,
    -- layer=1 filter=248 channel=74
    -2, 7, 2, 2, 6, -8, 7, -7, 9,
    -- layer=1 filter=248 channel=75
    5, 1, -5, 4, 3, 6, -21, 0, 6,
    -- layer=1 filter=248 channel=76
    -1, -7, -8, 4, 6, 9, -2, -5, -4,
    -- layer=1 filter=248 channel=77
    6, -7, -3, 5, -5, 0, -2, -4, -11,
    -- layer=1 filter=248 channel=78
    6, -2, -9, 1, -11, -8, -5, 9, 5,
    -- layer=1 filter=248 channel=79
    -1, -10, -9, 2, -2, -1, -9, -15, -1,
    -- layer=1 filter=248 channel=80
    3, 0, -5, -9, 0, 6, -5, 6, -9,
    -- layer=1 filter=248 channel=81
    0, -7, 4, -10, 2, 4, -8, -9, -6,
    -- layer=1 filter=248 channel=82
    0, -6, -11, -5, 7, 3, -5, -5, -5,
    -- layer=1 filter=248 channel=83
    -4, 8, 7, 1, -11, -11, 7, -7, 9,
    -- layer=1 filter=248 channel=84
    -4, -4, -1, -7, -9, -2, -5, -6, 0,
    -- layer=1 filter=248 channel=85
    -1, 3, 8, -3, -4, -4, -5, -2, 4,
    -- layer=1 filter=248 channel=86
    4, 4, 4, -13, -14, -9, -12, 5, -9,
    -- layer=1 filter=248 channel=87
    3, -4, 7, -1, -6, -3, -7, -4, -11,
    -- layer=1 filter=248 channel=88
    5, -11, -7, -3, -5, -1, -10, 4, 6,
    -- layer=1 filter=248 channel=89
    0, -1, -5, -2, -5, -8, -13, 6, -7,
    -- layer=1 filter=248 channel=90
    6, -9, -5, -1, 6, 2, -4, 6, -6,
    -- layer=1 filter=248 channel=91
    -1, -2, -11, -10, 0, -5, -14, 0, 4,
    -- layer=1 filter=248 channel=92
    -7, 7, -4, -1, 0, 8, -2, -8, 4,
    -- layer=1 filter=248 channel=93
    0, -2, 6, 0, -12, 4, 0, -13, 3,
    -- layer=1 filter=248 channel=94
    -10, 0, -9, -6, -11, -4, 1, 2, -11,
    -- layer=1 filter=248 channel=95
    -3, 5, 6, 11, 2, 10, -12, -8, 10,
    -- layer=1 filter=248 channel=96
    -4, -2, 8, -10, 0, 6, 3, 5, 2,
    -- layer=1 filter=248 channel=97
    -3, 8, 6, -1, 6, 0, 8, -10, -4,
    -- layer=1 filter=248 channel=98
    -9, 0, -7, 0, 0, 1, -2, -1, 1,
    -- layer=1 filter=248 channel=99
    -6, 8, -11, -11, -5, 6, -8, -4, -7,
    -- layer=1 filter=248 channel=100
    1, 0, 5, 6, 4, -1, -11, -5, -7,
    -- layer=1 filter=248 channel=101
    -3, 5, -5, 8, -5, 7, 7, -9, 5,
    -- layer=1 filter=248 channel=102
    7, 6, 7, -2, -3, 2, -4, -10, 3,
    -- layer=1 filter=248 channel=103
    -12, -3, -5, -1, -5, -3, -6, -5, -8,
    -- layer=1 filter=248 channel=104
    7, 1, -7, -11, -7, -6, -2, 3, -8,
    -- layer=1 filter=248 channel=105
    -6, 0, -12, 2, 2, -7, -5, 8, -2,
    -- layer=1 filter=248 channel=106
    -5, -4, -11, -16, 2, 6, 2, 6, -7,
    -- layer=1 filter=248 channel=107
    6, 4, 1, 4, 2, -7, -6, 4, 6,
    -- layer=1 filter=248 channel=108
    -21, 3, -11, -10, -1, -2, -1, 9, -10,
    -- layer=1 filter=248 channel=109
    -2, 7, 0, 1, 8, -5, -3, -4, 4,
    -- layer=1 filter=248 channel=110
    0, 5, -5, -4, -9, -2, -10, -1, 8,
    -- layer=1 filter=248 channel=111
    -8, -14, -3, -8, -6, 2, -1, -13, 10,
    -- layer=1 filter=248 channel=112
    -4, 6, 4, 1, -11, -6, -7, -6, 0,
    -- layer=1 filter=248 channel=113
    0, 2, -6, 0, 7, -2, 7, -1, -2,
    -- layer=1 filter=248 channel=114
    -12, -15, -4, -11, -1, 4, 13, -12, -3,
    -- layer=1 filter=248 channel=115
    6, -6, 2, -1, 1, -6, -12, 1, 6,
    -- layer=1 filter=248 channel=116
    -2, 9, -9, 1, -1, 6, 2, 5, 11,
    -- layer=1 filter=248 channel=117
    0, -13, -2, -1, 3, -9, -10, 0, 0,
    -- layer=1 filter=248 channel=118
    1, 7, -8, 4, 5, 7, 0, 4, 3,
    -- layer=1 filter=248 channel=119
    -6, -4, -6, -11, 1, 2, 3, 10, 0,
    -- layer=1 filter=248 channel=120
    -9, 0, 2, -3, -3, -7, -2, -5, -2,
    -- layer=1 filter=248 channel=121
    -12, 3, -16, 3, -11, -11, -4, -6, -12,
    -- layer=1 filter=248 channel=122
    -9, -3, -4, -2, 9, -9, 10, 0, -10,
    -- layer=1 filter=248 channel=123
    -6, -2, -11, 0, -10, -7, -9, 8, 2,
    -- layer=1 filter=248 channel=124
    6, -5, 7, -7, 4, 4, 9, -2, 5,
    -- layer=1 filter=248 channel=125
    2, 2, 5, 5, 4, 6, 1, 1, 0,
    -- layer=1 filter=248 channel=126
    -4, -5, -8, 5, -2, -10, 0, -4, -6,
    -- layer=1 filter=248 channel=127
    6, 9, 3, -6, 4, 3, -6, -6, 8,
    -- layer=1 filter=249 channel=0
    -4, -9, 3, -3, -8, -3, -6, -2, 1,
    -- layer=1 filter=249 channel=1
    -11, 3, -12, -5, 7, -6, -12, -8, -2,
    -- layer=1 filter=249 channel=2
    7, -11, 6, 11, 0, 0, -10, -10, -11,
    -- layer=1 filter=249 channel=3
    0, -4, 6, 5, 3, 11, -2, 3, -5,
    -- layer=1 filter=249 channel=4
    -10, -11, -2, -4, 2, -5, -12, -2, -7,
    -- layer=1 filter=249 channel=5
    0, 6, 1, 6, 8, 3, 7, 1, 10,
    -- layer=1 filter=249 channel=6
    -8, -3, 9, 0, -7, -2, -3, 6, -6,
    -- layer=1 filter=249 channel=7
    -2, 2, -10, -1, -6, -8, -6, -8, 4,
    -- layer=1 filter=249 channel=8
    1, 7, 1, 2, -9, 4, 2, 3, -4,
    -- layer=1 filter=249 channel=9
    1, -9, 0, 10, 1, 4, -2, 1, 6,
    -- layer=1 filter=249 channel=10
    7, -7, 7, -10, 6, 5, -8, -2, -5,
    -- layer=1 filter=249 channel=11
    -4, 0, 4, -9, -10, -2, -2, -10, 1,
    -- layer=1 filter=249 channel=12
    -3, 6, 2, -4, 5, 9, -9, -2, -8,
    -- layer=1 filter=249 channel=13
    0, 0, -8, 2, -2, 8, 1, -7, -8,
    -- layer=1 filter=249 channel=14
    0, -5, -2, 5, 6, -10, 0, 0, -6,
    -- layer=1 filter=249 channel=15
    7, 5, 8, -9, -4, 0, 1, 4, -1,
    -- layer=1 filter=249 channel=16
    2, 6, 5, -7, -2, -6, 1, -1, -8,
    -- layer=1 filter=249 channel=17
    -11, -2, -2, 0, -6, -3, 0, -11, 2,
    -- layer=1 filter=249 channel=18
    -8, -9, 0, -8, -11, -11, 7, -6, -7,
    -- layer=1 filter=249 channel=19
    -11, -3, -6, -6, -6, -2, -6, -12, 5,
    -- layer=1 filter=249 channel=20
    2, -1, 2, -2, 0, 3, -4, -7, -8,
    -- layer=1 filter=249 channel=21
    -7, 2, -1, -6, 7, -5, -1, 10, -6,
    -- layer=1 filter=249 channel=22
    -5, -10, 3, -2, -6, 0, -3, 0, -11,
    -- layer=1 filter=249 channel=23
    10, -7, -8, -9, -8, -5, -9, 6, 2,
    -- layer=1 filter=249 channel=24
    -6, -4, 0, 4, 0, 6, -4, 3, -4,
    -- layer=1 filter=249 channel=25
    -8, 7, 7, 1, -11, 4, -8, 0, 8,
    -- layer=1 filter=249 channel=26
    -9, -4, 6, 5, 2, 3, -6, -1, 6,
    -- layer=1 filter=249 channel=27
    -10, -4, 5, 5, -1, -10, -7, 2, 3,
    -- layer=1 filter=249 channel=28
    0, 3, -2, -3, 2, -10, -13, 0, 3,
    -- layer=1 filter=249 channel=29
    -10, 5, -11, 0, 3, -4, 3, 9, 0,
    -- layer=1 filter=249 channel=30
    -5, -6, 5, -13, 1, -8, 2, 5, 6,
    -- layer=1 filter=249 channel=31
    -10, -10, -4, -7, -3, -6, -6, -3, 7,
    -- layer=1 filter=249 channel=32
    7, -6, -2, 5, -11, -11, -3, -10, 0,
    -- layer=1 filter=249 channel=33
    -6, -1, 0, 10, -9, 0, -8, 8, -5,
    -- layer=1 filter=249 channel=34
    -10, 5, -8, -10, 0, -6, -10, -3, -11,
    -- layer=1 filter=249 channel=35
    0, 3, -5, 7, -2, 0, -3, -1, 2,
    -- layer=1 filter=249 channel=36
    3, -5, 6, -6, -1, 6, -3, -8, 4,
    -- layer=1 filter=249 channel=37
    -9, 5, 0, 5, -5, -8, -1, 0, -7,
    -- layer=1 filter=249 channel=38
    0, -9, 1, -2, 3, -8, -7, 0, 9,
    -- layer=1 filter=249 channel=39
    -1, 4, -5, 2, -9, -10, -11, -7, 8,
    -- layer=1 filter=249 channel=40
    -9, 0, 6, -11, 8, -3, 5, 1, 8,
    -- layer=1 filter=249 channel=41
    6, 7, -2, -5, 0, -7, 0, -2, 2,
    -- layer=1 filter=249 channel=42
    7, -6, -6, -6, 2, 0, -3, -10, -9,
    -- layer=1 filter=249 channel=43
    -4, 0, -4, -9, 3, -5, 3, 5, 1,
    -- layer=1 filter=249 channel=44
    -9, 0, -9, 0, 0, -10, 9, 5, 5,
    -- layer=1 filter=249 channel=45
    4, 0, 1, -9, 5, -9, -7, 3, 5,
    -- layer=1 filter=249 channel=46
    0, 4, -4, -1, 2, 2, -4, 1, -6,
    -- layer=1 filter=249 channel=47
    -3, -9, -8, -9, -4, -6, 8, 5, -8,
    -- layer=1 filter=249 channel=48
    1, 4, -8, 6, 2, 4, 1, 1, -11,
    -- layer=1 filter=249 channel=49
    3, -7, -4, 7, 1, 0, 6, -5, -10,
    -- layer=1 filter=249 channel=50
    5, -1, -8, -6, -10, 1, -6, 2, -7,
    -- layer=1 filter=249 channel=51
    -8, -9, 5, -1, 3, 5, 0, 4, -3,
    -- layer=1 filter=249 channel=52
    -5, -2, 5, 1, -8, 5, 0, 0, -9,
    -- layer=1 filter=249 channel=53
    7, -6, 9, -1, -8, 1, 8, -4, -4,
    -- layer=1 filter=249 channel=54
    -7, 3, 6, 0, -2, -5, 6, 3, -4,
    -- layer=1 filter=249 channel=55
    -10, -3, 0, 1, 1, -9, -9, -6, -6,
    -- layer=1 filter=249 channel=56
    0, -1, 3, -2, 1, -2, -1, 11, 0,
    -- layer=1 filter=249 channel=57
    2, -6, 8, -7, 6, -4, 5, -9, -7,
    -- layer=1 filter=249 channel=58
    -7, 0, -2, -5, 0, -6, -12, 0, 6,
    -- layer=1 filter=249 channel=59
    5, -4, 4, 5, 2, 9, 6, -9, -2,
    -- layer=1 filter=249 channel=60
    4, 2, 0, -10, -9, -6, -7, -1, 2,
    -- layer=1 filter=249 channel=61
    -1, 3, 7, -8, -1, -3, -2, -3, 7,
    -- layer=1 filter=249 channel=62
    -3, 1, 3, 5, 6, -12, 7, -3, 0,
    -- layer=1 filter=249 channel=63
    3, 6, -7, -12, 5, -12, 2, -4, -7,
    -- layer=1 filter=249 channel=64
    -6, 1, -6, -9, -3, 4, -3, -2, -9,
    -- layer=1 filter=249 channel=65
    -8, 2, -12, -6, -7, 6, 2, -6, 6,
    -- layer=1 filter=249 channel=66
    0, -1, 6, 6, 1, -12, 4, -7, -3,
    -- layer=1 filter=249 channel=67
    -1, 3, 9, -3, 3, 0, 7, -7, 5,
    -- layer=1 filter=249 channel=68
    1, -6, -6, 3, -12, 0, 0, -1, 0,
    -- layer=1 filter=249 channel=69
    -12, 9, 1, 4, 2, -2, -1, -1, 7,
    -- layer=1 filter=249 channel=70
    -2, -2, -6, 0, -5, 1, 5, 3, -4,
    -- layer=1 filter=249 channel=71
    2, -4, -4, 6, -7, -13, 6, -6, 5,
    -- layer=1 filter=249 channel=72
    -1, 2, -4, 5, 0, 3, -9, -7, 1,
    -- layer=1 filter=249 channel=73
    -5, -7, -9, -4, 0, -11, -5, -7, -1,
    -- layer=1 filter=249 channel=74
    -7, 1, -8, 1, 7, 0, -2, 0, 5,
    -- layer=1 filter=249 channel=75
    -2, 10, 5, -4, -7, -5, 1, 3, 3,
    -- layer=1 filter=249 channel=76
    -8, 5, 7, -3, 1, -2, -9, 5, -5,
    -- layer=1 filter=249 channel=77
    0, 6, -6, -1, -10, 0, 8, -7, -2,
    -- layer=1 filter=249 channel=78
    -10, -1, 3, 5, 5, 3, 5, 6, -5,
    -- layer=1 filter=249 channel=79
    -10, -12, 7, 4, 3, -4, 3, 6, -5,
    -- layer=1 filter=249 channel=80
    -1, -4, 7, -10, -12, -4, 6, 2, -2,
    -- layer=1 filter=249 channel=81
    -4, 1, 1, -9, -1, 4, -7, -12, 6,
    -- layer=1 filter=249 channel=82
    -8, 0, 7, 2, 0, -2, -2, 6, -2,
    -- layer=1 filter=249 channel=83
    -3, -9, -3, 6, -2, -7, -8, -3, 7,
    -- layer=1 filter=249 channel=84
    -10, 4, 0, -7, -6, -11, -2, -1, -8,
    -- layer=1 filter=249 channel=85
    -5, -6, 1, -11, 4, 7, 8, -7, -3,
    -- layer=1 filter=249 channel=86
    -2, 5, -7, -10, -12, 8, -10, -14, -8,
    -- layer=1 filter=249 channel=87
    4, -9, 8, -8, -10, -2, -8, -1, -9,
    -- layer=1 filter=249 channel=88
    -6, -1, 4, 10, -9, 7, 1, 0, 7,
    -- layer=1 filter=249 channel=89
    -2, -6, -1, 4, 8, -1, 9, 5, 2,
    -- layer=1 filter=249 channel=90
    -7, 2, -1, -7, 0, 2, 2, -1, 1,
    -- layer=1 filter=249 channel=91
    6, -7, -5, -10, 0, 0, 7, 4, -8,
    -- layer=1 filter=249 channel=92
    -5, 5, 6, 3, 5, 4, 1, -5, -4,
    -- layer=1 filter=249 channel=93
    -7, 4, 5, -9, -9, 8, 1, 7, -4,
    -- layer=1 filter=249 channel=94
    -12, 5, -3, -3, 5, 1, 5, -10, 0,
    -- layer=1 filter=249 channel=95
    10, -8, 4, 3, 2, -6, 9, -5, -4,
    -- layer=1 filter=249 channel=96
    0, -1, 8, -1, -10, -1, -12, -7, -7,
    -- layer=1 filter=249 channel=97
    -3, -9, -12, 0, 8, -4, -7, -11, 1,
    -- layer=1 filter=249 channel=98
    5, -1, -6, 2, -3, -9, 1, -12, -3,
    -- layer=1 filter=249 channel=99
    4, 8, 8, 7, 6, 5, 6, -8, -2,
    -- layer=1 filter=249 channel=100
    -7, -3, 1, -8, -5, 3, -10, -6, -4,
    -- layer=1 filter=249 channel=101
    2, 1, -7, 5, 1, 0, 0, 0, 7,
    -- layer=1 filter=249 channel=102
    -4, -3, -3, 5, -2, -12, -2, -5, -4,
    -- layer=1 filter=249 channel=103
    6, 5, -1, 5, -5, -4, 1, -8, 8,
    -- layer=1 filter=249 channel=104
    -6, 8, -8, 0, 7, 1, -9, -5, -5,
    -- layer=1 filter=249 channel=105
    -9, -2, 2, 3, -9, -5, -6, -11, 1,
    -- layer=1 filter=249 channel=106
    -5, -7, -7, 2, 1, 3, 0, -1, -10,
    -- layer=1 filter=249 channel=107
    7, 0, 7, -8, -6, -6, 7, 11, -6,
    -- layer=1 filter=249 channel=108
    -1, -13, -5, -2, -1, 10, 0, -1, 6,
    -- layer=1 filter=249 channel=109
    3, 9, -9, -8, -6, 10, 6, -3, 6,
    -- layer=1 filter=249 channel=110
    6, -2, -8, 0, 2, 7, -3, -8, -7,
    -- layer=1 filter=249 channel=111
    4, 0, -7, -13, 4, -3, -9, -6, -9,
    -- layer=1 filter=249 channel=112
    -7, -2, -4, 7, -9, 5, 0, 5, 0,
    -- layer=1 filter=249 channel=113
    -2, -12, 0, -10, -3, -5, -5, -1, -5,
    -- layer=1 filter=249 channel=114
    -1, -6, 4, 1, 2, 1, -7, 8, 8,
    -- layer=1 filter=249 channel=115
    3, 4, -11, 3, -3, -8, 4, 3, -4,
    -- layer=1 filter=249 channel=116
    -4, 0, -4, 3, 9, 2, -2, 0, -9,
    -- layer=1 filter=249 channel=117
    2, -6, -3, -5, -3, -8, 4, -8, 6,
    -- layer=1 filter=249 channel=118
    -3, -1, 2, 8, 4, -6, -2, -9, 7,
    -- layer=1 filter=249 channel=119
    -1, -1, 2, -8, -6, 0, 5, -11, -2,
    -- layer=1 filter=249 channel=120
    -6, -3, 0, -1, 0, 2, 6, -12, -8,
    -- layer=1 filter=249 channel=121
    7, 3, -9, -2, -10, 0, -4, 3, -3,
    -- layer=1 filter=249 channel=122
    3, -5, -8, 9, 8, -5, 5, 1, 6,
    -- layer=1 filter=249 channel=123
    -7, -2, -4, 6, 6, 7, -4, 0, 5,
    -- layer=1 filter=249 channel=124
    -3, -10, -1, -4, -3, -11, -1, 2, 7,
    -- layer=1 filter=249 channel=125
    -8, -10, 9, 6, -8, -9, 0, 5, -6,
    -- layer=1 filter=249 channel=126
    4, -3, -4, 3, -8, 7, 0, -11, -11,
    -- layer=1 filter=249 channel=127
    -8, 3, 6, -4, -5, -10, -5, 10, 4,
    -- layer=1 filter=250 channel=0
    -12, -5, -14, -7, -4, -11, -2, -23, -24,
    -- layer=1 filter=250 channel=1
    -50, -49, -48, 16, -19, -49, -3, 12, -22,
    -- layer=1 filter=250 channel=2
    41, 26, -25, 41, 8, -11, 35, 3, -14,
    -- layer=1 filter=250 channel=3
    6, -5, -3, -2, -16, 3, 5, -2, 6,
    -- layer=1 filter=250 channel=4
    -6, 0, 2, -10, 5, -19, -8, -2, -7,
    -- layer=1 filter=250 channel=5
    -36, -61, -87, 56, 19, -19, -24, -1, 3,
    -- layer=1 filter=250 channel=6
    1, 6, 2, -10, 22, 63, -24, 2, 25,
    -- layer=1 filter=250 channel=7
    -6, -8, -11, 26, 12, -10, 5, 13, 15,
    -- layer=1 filter=250 channel=8
    -47, -56, -48, 51, -1, -23, 16, 12, -19,
    -- layer=1 filter=250 channel=9
    3, -1, 0, -32, -33, -15, -47, -106, -27,
    -- layer=1 filter=250 channel=10
    16, 15, -22, 25, 17, -3, 13, 9, 9,
    -- layer=1 filter=250 channel=11
    4, 2, 4, 12, 38, 17, 17, 22, 13,
    -- layer=1 filter=250 channel=12
    10, -27, -23, 24, 74, 46, -3, -7, 2,
    -- layer=1 filter=250 channel=13
    -13, 3, 46, -26, -8, 28, -25, -17, 8,
    -- layer=1 filter=250 channel=14
    -7, -31, -18, 19, 39, -23, 47, -3, 7,
    -- layer=1 filter=250 channel=15
    -17, -47, -7, 67, 26, -10, 44, 55, 37,
    -- layer=1 filter=250 channel=16
    -57, -44, -51, 69, 9, 9, -6, 13, 1,
    -- layer=1 filter=250 channel=17
    13, 2, 36, -22, -42, -29, -12, -33, -34,
    -- layer=1 filter=250 channel=18
    16, 0, -18, 5, 61, 45, -22, -21, 22,
    -- layer=1 filter=250 channel=19
    -33, -94, -44, 15, -13, -3, -55, -99, 36,
    -- layer=1 filter=250 channel=20
    4, 23, 44, -12, 8, 30, -31, -3, 0,
    -- layer=1 filter=250 channel=21
    -31, -25, -28, 3, -8, -7, 28, 10, -18,
    -- layer=1 filter=250 channel=22
    -7, 17, 40, 0, 4, 11, -5, 2, 3,
    -- layer=1 filter=250 channel=23
    36, -11, -12, 73, 9, 23, 37, 57, 11,
    -- layer=1 filter=250 channel=24
    -80, -107, -35, -18, -46, -68, 51, -9, -5,
    -- layer=1 filter=250 channel=25
    -40, -8, -9, 17, -27, -5, -5, -20, -6,
    -- layer=1 filter=250 channel=26
    -25, -73, 32, 14, -42, -27, 43, 14, 2,
    -- layer=1 filter=250 channel=27
    23, 23, 9, 39, 52, 39, 9, 29, 28,
    -- layer=1 filter=250 channel=28
    -48, -5, -24, 15, -10, -41, 10, -15, -18,
    -- layer=1 filter=250 channel=29
    19, -2, -7, 1, -5, -5, -16, -35, -24,
    -- layer=1 filter=250 channel=30
    23, -18, -41, -8, 42, 37, -84, -36, -9,
    -- layer=1 filter=250 channel=31
    62, 42, 0, 33, 56, 47, -49, 35, 38,
    -- layer=1 filter=250 channel=32
    7, -74, 1, 34, -14, -15, 37, 38, -21,
    -- layer=1 filter=250 channel=33
    23, 14, 5, 9, 11, 12, 26, 0, 5,
    -- layer=1 filter=250 channel=34
    -17, -20, -26, -2, -15, 7, 6, 7, -4,
    -- layer=1 filter=250 channel=35
    -5, 8, 9, 17, 12, 13, 8, 9, 8,
    -- layer=1 filter=250 channel=36
    5, 0, 1, 14, 31, 5, 6, 17, 1,
    -- layer=1 filter=250 channel=37
    -55, -67, -37, 58, 2, -9, -5, 5, 43,
    -- layer=1 filter=250 channel=38
    0, 12, 17, -28, 23, 37, -37, -10, 13,
    -- layer=1 filter=250 channel=39
    0, 1, 7, -3, 3, 8, -14, 14, -3,
    -- layer=1 filter=250 channel=40
    53, 57, 12, -28, 71, 58, -48, 10, 24,
    -- layer=1 filter=250 channel=41
    -14, -75, 6, -9, -52, -60, 2, -26, -61,
    -- layer=1 filter=250 channel=42
    33, -2, -26, 36, 15, -2, 0, 13, -2,
    -- layer=1 filter=250 channel=43
    -56, -33, -53, 35, -37, -12, 9, 12, -3,
    -- layer=1 filter=250 channel=44
    -25, -75, 19, 26, -48, -29, 47, 52, -11,
    -- layer=1 filter=250 channel=45
    -56, -43, 11, 12, 7, -3, 29, 40, 19,
    -- layer=1 filter=250 channel=46
    -8, -38, -63, 60, 50, 36, -30, -3, 60,
    -- layer=1 filter=250 channel=47
    29, -18, -27, 58, 28, -3, 12, 22, 2,
    -- layer=1 filter=250 channel=48
    0, 0, -5, -22, -5, -11, 3, -2, -2,
    -- layer=1 filter=250 channel=49
    15, 18, -1, 10, 13, 0, 4, -4, 11,
    -- layer=1 filter=250 channel=50
    9, 1, -7, -3, -13, 5, -5, -4, -11,
    -- layer=1 filter=250 channel=51
    7, 9, 9, -11, 21, 13, -6, 3, 1,
    -- layer=1 filter=250 channel=52
    -15, -15, -15, 9, -26, -2, -7, -1, -3,
    -- layer=1 filter=250 channel=53
    8, -16, 1, 0, 11, 5, 16, 27, 16,
    -- layer=1 filter=250 channel=54
    -36, -39, -24, 44, -41, 0, -17, -36, 6,
    -- layer=1 filter=250 channel=55
    13, -19, -6, 39, 26, -5, 27, 51, 0,
    -- layer=1 filter=250 channel=56
    -7, -3, 7, 9, -3, 12, 9, 6, 10,
    -- layer=1 filter=250 channel=57
    43, 57, 27, 21, 40, 15, -13, 8, 26,
    -- layer=1 filter=250 channel=58
    29, -21, 15, 23, 25, 0, 14, 27, 17,
    -- layer=1 filter=250 channel=59
    -6, 5, 8, -4, -19, 5, -6, -12, -12,
    -- layer=1 filter=250 channel=60
    3, -3, -5, 2, 1, 3, 2, -11, 10,
    -- layer=1 filter=250 channel=61
    13, -3, 12, 0, -1, -9, 3, 9, -15,
    -- layer=1 filter=250 channel=62
    -65, -56, -29, 48, -14, -27, -1, -11, -1,
    -- layer=1 filter=250 channel=63
    -15, -9, -16, 5, 14, -7, 7, 0, -24,
    -- layer=1 filter=250 channel=64
    3, -5, 15, -19, -6, 1, -13, 3, -1,
    -- layer=1 filter=250 channel=65
    -23, 0, -11, -2, 3, 14, -2, -11, -21,
    -- layer=1 filter=250 channel=66
    -4, -4, -8, 4, 6, -12, 10, 5, -22,
    -- layer=1 filter=250 channel=67
    2, -22, -16, -37, -1, -19, -31, -14, -28,
    -- layer=1 filter=250 channel=68
    -55, -65, 22, 17, -72, -22, 61, 47, 5,
    -- layer=1 filter=250 channel=69
    -52, -100, -27, 38, 44, -14, 17, 31, 42,
    -- layer=1 filter=250 channel=70
    34, 1, -42, 5, 12, 14, -14, 54, 33,
    -- layer=1 filter=250 channel=71
    -53, -68, -79, 15, -34, -33, 22, 1, -6,
    -- layer=1 filter=250 channel=72
    0, -33, -44, -18, 10, 0, -97, -46, -24,
    -- layer=1 filter=250 channel=73
    0, -9, 6, 10, 6, 0, 3, -3, 0,
    -- layer=1 filter=250 channel=74
    -20, 14, 17, -14, -6, 35, 4, -5, 25,
    -- layer=1 filter=250 channel=75
    19, -43, -37, 35, 62, 35, -70, -9, -34,
    -- layer=1 filter=250 channel=76
    -30, -37, 7, 0, -23, 12, 0, -13, -30,
    -- layer=1 filter=250 channel=77
    -54, -59, -31, -28, -46, -46, 37, 0, -28,
    -- layer=1 filter=250 channel=78
    24, 2, -13, 5, -8, -4, 15, -29, 4,
    -- layer=1 filter=250 channel=79
    -55, -47, -36, 50, 12, -17, 0, 0, 16,
    -- layer=1 filter=250 channel=80
    17, 2, -7, 12, -2, 19, 3, 23, 11,
    -- layer=1 filter=250 channel=81
    -73, -103, -74, -1, -72, -68, 64, 6, -5,
    -- layer=1 filter=250 channel=82
    -21, 0, 5, -7, -8, 10, 22, 4, 6,
    -- layer=1 filter=250 channel=83
    -31, -50, 19, 16, 2, -42, 37, 53, 25,
    -- layer=1 filter=250 channel=84
    -9, -10, -10, 4, 27, 36, -17, -49, -29,
    -- layer=1 filter=250 channel=85
    2, -11, 8, 18, 17, -39, 1, 14, 18,
    -- layer=1 filter=250 channel=86
    17, 21, 5, 30, 19, 7, -36, -1, -22,
    -- layer=1 filter=250 channel=87
    32, -35, -18, 23, -12, 1, -72, -61, 80,
    -- layer=1 filter=250 channel=88
    5, 12, -16, 10, 7, -10, 3, 0, -3,
    -- layer=1 filter=250 channel=89
    -26, -23, -14, -7, -15, 11, 21, 17, -18,
    -- layer=1 filter=250 channel=90
    -38, -86, 38, 9, -62, -20, 67, 45, 32,
    -- layer=1 filter=250 channel=91
    19, 23, 27, -32, 26, 47, -50, -22, 8,
    -- layer=1 filter=250 channel=92
    -27, -38, 30, 32, 0, 6, 62, 38, -1,
    -- layer=1 filter=250 channel=93
    -29, -40, -12, -13, -46, -47, 21, -2, -28,
    -- layer=1 filter=250 channel=94
    -13, 1, -13, 6, 4, 8, -17, -47, -30,
    -- layer=1 filter=250 channel=95
    -14, -27, -46, 17, 38, 38, -58, -31, -33,
    -- layer=1 filter=250 channel=96
    11, 1, -13, 2, -4, -15, 9, 3, -10,
    -- layer=1 filter=250 channel=97
    -37, -18, -13, -16, -57, -29, 26, -15, -31,
    -- layer=1 filter=250 channel=98
    -41, -23, -4, 28, -14, -35, 12, 14, 2,
    -- layer=1 filter=250 channel=99
    26, 28, 3, 33, 2, -17, 69, 19, 51,
    -- layer=1 filter=250 channel=100
    1, 5, 8, 22, 33, 8, -11, 1, 1,
    -- layer=1 filter=250 channel=101
    5, 22, 25, -20, 19, 17, -31, -10, 3,
    -- layer=1 filter=250 channel=102
    -18, 5, -12, -13, 12, 8, -55, -72, -52,
    -- layer=1 filter=250 channel=103
    26, 26, 29, 24, 33, 50, -1, 18, 20,
    -- layer=1 filter=250 channel=104
    47, 10, 9, 40, 8, 0, -4, 22, -14,
    -- layer=1 filter=250 channel=105
    -23, 0, -22, -23, -20, -29, 15, -26, -29,
    -- layer=1 filter=250 channel=106
    1, -7, 23, -15, -1, 20, 11, 12, 8,
    -- layer=1 filter=250 channel=107
    -4, -11, -16, -6, 2, -10, 3, 14, 9,
    -- layer=1 filter=250 channel=108
    -5, -93, 17, 35, -1, -43, 56, 72, 3,
    -- layer=1 filter=250 channel=109
    -5, 5, 10, 5, 4, 3, -3, 7, -3,
    -- layer=1 filter=250 channel=110
    3, 0, 6, -1, 11, -2, 6, -15, 5,
    -- layer=1 filter=250 channel=111
    16, -8, -39, -4, 52, 23, -47, -53, 18,
    -- layer=1 filter=250 channel=112
    -12, -41, -38, 10, 32, 9, -18, 10, 21,
    -- layer=1 filter=250 channel=113
    0, 20, -6, 31, 33, 25, -2, 53, 4,
    -- layer=1 filter=250 channel=114
    -5, -9, -7, 71, 51, 27, 3, 38, 18,
    -- layer=1 filter=250 channel=115
    29, 33, 11, 7, 26, 3, -27, -18, 5,
    -- layer=1 filter=250 channel=116
    -1, -3, 6, 9, -11, -7, 6, -7, 8,
    -- layer=1 filter=250 channel=117
    19, -13, -14, 22, 73, 39, 18, 17, 98,
    -- layer=1 filter=250 channel=118
    14, 13, -15, -15, 10, 47, -30, -38, 2,
    -- layer=1 filter=250 channel=119
    -28, -115, 15, 20, -56, -42, 65, 33, -7,
    -- layer=1 filter=250 channel=120
    -11, -1, 0, 10, -12, -23, 4, -15, 0,
    -- layer=1 filter=250 channel=121
    29, -5, -30, 33, 69, 11, -69, -20, 1,
    -- layer=1 filter=250 channel=122
    2, -6, 0, -2, -2, -4, 7, -5, 9,
    -- layer=1 filter=250 channel=123
    11, -23, -13, 35, 53, 5, -19, 37, 31,
    -- layer=1 filter=250 channel=124
    -1, -1, -2, 18, -3, -2, 0, 3, 0,
    -- layer=1 filter=250 channel=125
    37, 33, 0, -25, 32, -14, -24, 25, 51,
    -- layer=1 filter=250 channel=126
    -42, -63, -14, 17, -22, -71, 59, 51, 14,
    -- layer=1 filter=250 channel=127
    23, 9, -18, 19, 42, 51, -48, -25, 10,
    -- layer=1 filter=251 channel=0
    -7, 4, 4, -1, 2, -5, 4, -1, 7,
    -- layer=1 filter=251 channel=1
    3, -3, 6, -3, -7, 0, -9, 1, 6,
    -- layer=1 filter=251 channel=2
    -7, 7, 5, 5, 5, -9, -1, -8, -12,
    -- layer=1 filter=251 channel=3
    -7, 8, 8, 9, 0, -6, 0, 10, 1,
    -- layer=1 filter=251 channel=4
    2, 6, 1, 5, -5, -11, -9, 7, 0,
    -- layer=1 filter=251 channel=5
    -2, -11, -3, -1, -10, -3, 6, -6, -9,
    -- layer=1 filter=251 channel=6
    7, -4, 8, 6, 2, 8, 2, 8, 5,
    -- layer=1 filter=251 channel=7
    1, -8, 7, -8, -4, 6, -2, -5, 9,
    -- layer=1 filter=251 channel=8
    -4, 8, -8, -8, -8, 4, 1, -2, -7,
    -- layer=1 filter=251 channel=9
    -3, -2, 4, -4, -9, 7, 5, -10, 7,
    -- layer=1 filter=251 channel=10
    -6, 0, -6, 10, -3, -3, 0, 7, -2,
    -- layer=1 filter=251 channel=11
    0, -13, -5, 2, -1, -11, -12, 0, 9,
    -- layer=1 filter=251 channel=12
    -5, 7, -5, -9, -7, -1, 1, 7, 0,
    -- layer=1 filter=251 channel=13
    -9, 2, 3, -2, -6, 4, 2, -3, 3,
    -- layer=1 filter=251 channel=14
    -9, 7, -8, 2, 0, -1, 1, -5, -4,
    -- layer=1 filter=251 channel=15
    7, -11, -11, -8, 2, -3, -7, 6, 3,
    -- layer=1 filter=251 channel=16
    -3, -7, -11, 4, 2, 6, -10, 3, 1,
    -- layer=1 filter=251 channel=17
    4, -10, -10, -9, -5, -10, -8, -9, -1,
    -- layer=1 filter=251 channel=18
    -10, -4, -1, 7, 7, 1, -7, -1, -5,
    -- layer=1 filter=251 channel=19
    -4, -6, -4, -5, 1, 4, 3, -4, 0,
    -- layer=1 filter=251 channel=20
    -4, -8, 2, 7, 4, 6, 8, -5, -11,
    -- layer=1 filter=251 channel=21
    -8, -11, 6, -11, -1, -1, 8, -6, 4,
    -- layer=1 filter=251 channel=22
    -10, 1, 2, 3, 0, 6, 1, 8, -1,
    -- layer=1 filter=251 channel=23
    0, 2, 2, 0, 4, -3, 1, 5, -1,
    -- layer=1 filter=251 channel=24
    -5, -9, -2, -11, 1, 1, 5, -7, 6,
    -- layer=1 filter=251 channel=25
    -5, 2, -6, -10, -1, -6, 9, -8, -1,
    -- layer=1 filter=251 channel=26
    0, 9, -10, -9, 5, -10, 0, -7, 4,
    -- layer=1 filter=251 channel=27
    -4, -5, 9, -2, -9, -3, 2, 8, -1,
    -- layer=1 filter=251 channel=28
    5, -2, -7, 5, -1, 3, -7, -10, 7,
    -- layer=1 filter=251 channel=29
    5, 6, 5, -8, 0, 1, -4, -9, -4,
    -- layer=1 filter=251 channel=30
    -2, -12, -7, 4, 4, 0, -1, 10, -7,
    -- layer=1 filter=251 channel=31
    2, 3, 5, -6, 1, 1, 0, -11, -6,
    -- layer=1 filter=251 channel=32
    -12, -9, -8, -11, 0, 6, 4, -3, -4,
    -- layer=1 filter=251 channel=33
    8, 8, -8, -1, 8, -1, 0, 4, 4,
    -- layer=1 filter=251 channel=34
    -6, 3, -9, -9, 7, 9, 4, -10, -12,
    -- layer=1 filter=251 channel=35
    -6, 6, 4, 5, 10, -6, 0, 3, 0,
    -- layer=1 filter=251 channel=36
    8, -7, -8, 4, 3, -10, -7, 0, 2,
    -- layer=1 filter=251 channel=37
    8, -9, -10, -3, 4, 10, -4, -3, 9,
    -- layer=1 filter=251 channel=38
    5, 0, -4, -3, -3, 1, -1, -7, 1,
    -- layer=1 filter=251 channel=39
    3, -4, 2, -5, -5, 8, 3, 7, 2,
    -- layer=1 filter=251 channel=40
    0, -14, -4, 10, 9, -9, -10, 6, 0,
    -- layer=1 filter=251 channel=41
    -3, 6, -1, -10, 0, 5, 2, -1, 0,
    -- layer=1 filter=251 channel=42
    1, -4, -9, 7, -4, 3, -10, -3, 0,
    -- layer=1 filter=251 channel=43
    2, 7, -6, -11, 0, -7, -11, 8, -9,
    -- layer=1 filter=251 channel=44
    -3, -7, -11, 7, 0, 5, -8, 3, -6,
    -- layer=1 filter=251 channel=45
    7, -5, 6, -1, -10, -10, 0, 2, -12,
    -- layer=1 filter=251 channel=46
    -4, -4, 4, 10, 2, 0, 6, -2, 0,
    -- layer=1 filter=251 channel=47
    3, -7, 8, -2, -2, 1, 8, 4, 2,
    -- layer=1 filter=251 channel=48
    -3, -6, 1, 9, 0, -2, 8, -9, -10,
    -- layer=1 filter=251 channel=49
    0, -5, 6, -6, 0, 1, -6, -1, 7,
    -- layer=1 filter=251 channel=50
    0, -5, -8, -9, -5, -5, 0, 5, -10,
    -- layer=1 filter=251 channel=51
    9, -6, 4, 6, 1, -5, -11, 5, -1,
    -- layer=1 filter=251 channel=52
    -5, 8, -10, 6, -5, -2, -9, -1, -9,
    -- layer=1 filter=251 channel=53
    3, 3, -2, -9, -7, -9, -7, -8, -5,
    -- layer=1 filter=251 channel=54
    -11, 5, -5, -5, -8, 5, -7, -11, -2,
    -- layer=1 filter=251 channel=55
    -5, -3, -3, -6, -10, -6, -5, 7, -7,
    -- layer=1 filter=251 channel=56
    9, -1, -2, -4, 2, 8, 7, -5, 0,
    -- layer=1 filter=251 channel=57
    -11, 3, 9, -1, -11, -1, 0, 0, -10,
    -- layer=1 filter=251 channel=58
    1, 0, -6, 7, 0, -1, -2, -3, -5,
    -- layer=1 filter=251 channel=59
    -3, 4, -10, 6, -5, -7, 4, -12, -4,
    -- layer=1 filter=251 channel=60
    -10, 4, -6, -4, 9, 9, -3, 3, -7,
    -- layer=1 filter=251 channel=61
    -1, -6, 9, 9, 8, 9, -9, -8, -6,
    -- layer=1 filter=251 channel=62
    9, -11, 5, -4, 0, 0, -2, 8, -4,
    -- layer=1 filter=251 channel=63
    0, -11, 1, -2, 7, -6, -9, -7, -6,
    -- layer=1 filter=251 channel=64
    3, -9, 6, -10, -6, 3, -3, -5, -3,
    -- layer=1 filter=251 channel=65
    3, 4, -8, -3, -10, -7, -11, 4, -10,
    -- layer=1 filter=251 channel=66
    -10, 7, -11, -9, 2, -8, 3, -9, 2,
    -- layer=1 filter=251 channel=67
    0, 8, 9, 0, 1, 7, -2, 0, 6,
    -- layer=1 filter=251 channel=68
    2, -4, -1, 2, -2, 2, -4, -5, 0,
    -- layer=1 filter=251 channel=69
    -8, -4, 3, 3, 3, -9, 4, 3, -4,
    -- layer=1 filter=251 channel=70
    1, 0, -3, -11, 6, -6, 0, 0, -3,
    -- layer=1 filter=251 channel=71
    2, -5, 1, -11, 0, 8, -9, 1, -3,
    -- layer=1 filter=251 channel=72
    -3, -10, 4, -9, -9, -5, -2, 0, -5,
    -- layer=1 filter=251 channel=73
    -2, 1, -4, 1, -8, 2, -7, 4, -7,
    -- layer=1 filter=251 channel=74
    -4, -6, 6, 4, 0, 2, -8, -2, 2,
    -- layer=1 filter=251 channel=75
    -1, 0, -3, 6, 0, -7, 3, 0, -8,
    -- layer=1 filter=251 channel=76
    1, -8, 0, 6, -1, 0, -12, -6, -6,
    -- layer=1 filter=251 channel=77
    2, -5, 5, -9, -5, 6, -7, 7, 1,
    -- layer=1 filter=251 channel=78
    2, -8, -7, 4, -1, 1, -1, -1, -6,
    -- layer=1 filter=251 channel=79
    5, -10, -6, 4, -10, 0, -4, 4, 2,
    -- layer=1 filter=251 channel=80
    4, -5, 0, 7, -3, -5, 5, 10, 0,
    -- layer=1 filter=251 channel=81
    6, 6, -4, -12, 5, 11, 5, -11, 4,
    -- layer=1 filter=251 channel=82
    -10, 6, -9, -8, -6, 6, -11, -2, 3,
    -- layer=1 filter=251 channel=83
    0, 0, -6, 5, -6, 0, 0, 8, -1,
    -- layer=1 filter=251 channel=84
    5, 6, -3, 7, -9, 1, -6, 2, -6,
    -- layer=1 filter=251 channel=85
    -1, -4, 0, 5, -6, 0, -3, -7, 3,
    -- layer=1 filter=251 channel=86
    4, -9, -4, 8, -6, -4, 5, 5, 0,
    -- layer=1 filter=251 channel=87
    6, 4, 0, -6, 8, -8, -11, 0, 0,
    -- layer=1 filter=251 channel=88
    0, -4, 7, 6, 8, 1, -2, 6, -6,
    -- layer=1 filter=251 channel=89
    -8, 1, -10, -6, 4, 2, -7, -7, -9,
    -- layer=1 filter=251 channel=90
    2, -9, 1, -6, -10, -11, 6, 6, -5,
    -- layer=1 filter=251 channel=91
    -3, -12, 5, -6, 0, 2, -1, -9, -6,
    -- layer=1 filter=251 channel=92
    7, 0, -1, 5, -3, 7, -7, -7, 8,
    -- layer=1 filter=251 channel=93
    -4, 0, 1, 3, -2, -8, -3, -3, 7,
    -- layer=1 filter=251 channel=94
    6, -4, -4, -4, 0, 0, -11, -1, -10,
    -- layer=1 filter=251 channel=95
    -12, -2, -1, -11, -2, -3, 7, -5, -1,
    -- layer=1 filter=251 channel=96
    2, 0, -2, -6, 2, -1, -11, 2, -5,
    -- layer=1 filter=251 channel=97
    -5, 1, 0, 6, 4, -6, -6, -9, -3,
    -- layer=1 filter=251 channel=98
    0, 1, 5, -11, 0, 3, -7, 0, 7,
    -- layer=1 filter=251 channel=99
    4, -4, -9, -3, -5, -10, -7, 7, -9,
    -- layer=1 filter=251 channel=100
    5, 6, 0, -4, -6, -11, -6, 5, 8,
    -- layer=1 filter=251 channel=101
    -1, 0, -1, 0, -5, -5, 6, -2, -8,
    -- layer=1 filter=251 channel=102
    -10, 8, 2, 7, -3, -11, -7, -1, -6,
    -- layer=1 filter=251 channel=103
    -2, 8, 4, 3, 4, -3, -1, -11, -6,
    -- layer=1 filter=251 channel=104
    -3, 8, 7, 0, -5, 3, 1, 9, -5,
    -- layer=1 filter=251 channel=105
    0, 0, 6, 2, 3, -8, -10, -8, 1,
    -- layer=1 filter=251 channel=106
    -8, -11, -11, -1, 5, -10, -5, 3, -4,
    -- layer=1 filter=251 channel=107
    7, -2, 1, -8, 4, -6, -3, 3, 7,
    -- layer=1 filter=251 channel=108
    5, -10, 0, 2, 0, 8, 1, -3, -2,
    -- layer=1 filter=251 channel=109
    4, 8, -8, 1, -6, -10, 1, 0, 4,
    -- layer=1 filter=251 channel=110
    -9, -1, -7, -6, 6, 2, 0, -11, 8,
    -- layer=1 filter=251 channel=111
    -11, 0, 1, -6, -6, -2, -6, 2, -5,
    -- layer=1 filter=251 channel=112
    -5, -5, -4, 2, -11, -6, 7, 6, -1,
    -- layer=1 filter=251 channel=113
    -1, -9, -11, 5, -4, -11, 5, -3, 7,
    -- layer=1 filter=251 channel=114
    -2, 0, -4, 5, -10, -9, 2, -1, 6,
    -- layer=1 filter=251 channel=115
    7, 2, -6, 3, -10, 5, 0, -4, -8,
    -- layer=1 filter=251 channel=116
    3, -3, -1, 5, -7, 5, 9, -3, -6,
    -- layer=1 filter=251 channel=117
    4, 1, -13, -1, 3, 3, 6, 10, 0,
    -- layer=1 filter=251 channel=118
    5, 6, 2, -9, 7, 8, -2, 7, 0,
    -- layer=1 filter=251 channel=119
    2, -6, 8, 4, 3, -8, -7, 5, -11,
    -- layer=1 filter=251 channel=120
    8, 6, -8, -1, 3, 7, -2, 4, -10,
    -- layer=1 filter=251 channel=121
    -3, 2, -5, -1, 8, 8, -7, -7, 1,
    -- layer=1 filter=251 channel=122
    9, -5, -4, 0, -2, 8, 2, -9, 9,
    -- layer=1 filter=251 channel=123
    7, -9, 2, -3, -4, -5, -10, -12, -1,
    -- layer=1 filter=251 channel=124
    7, -9, -4, 4, -4, -5, -1, 4, 6,
    -- layer=1 filter=251 channel=125
    -4, 8, -5, -5, 3, -7, -7, 0, 9,
    -- layer=1 filter=251 channel=126
    -3, 3, 7, -2, 7, 9, 8, 8, 3,
    -- layer=1 filter=251 channel=127
    -12, 2, -2, -10, -1, -1, -4, -3, 2,
    -- layer=1 filter=252 channel=0
    -26, -8, -12, -18, -37, -9, -20, -27, -10,
    -- layer=1 filter=252 channel=1
    7, -10, 9, -35, -17, -40, 6, 11, 4,
    -- layer=1 filter=252 channel=2
    2, 30, 0, 12, 11, 16, 22, 17, 7,
    -- layer=1 filter=252 channel=3
    0, -2, 0, -8, 0, 11, 5, 13, 0,
    -- layer=1 filter=252 channel=4
    6, 5, 6, 1, -1, 0, -5, 0, -1,
    -- layer=1 filter=252 channel=5
    -52, -41, -37, -128, -127, -103, 55, 61, 37,
    -- layer=1 filter=252 channel=6
    -4, -6, -7, 30, 33, 22, 38, 46, 30,
    -- layer=1 filter=252 channel=7
    -33, -2, 33, -39, 9, 0, -21, 1, 4,
    -- layer=1 filter=252 channel=8
    21, 21, 36, -68, -56, -61, 9, 6, -25,
    -- layer=1 filter=252 channel=9
    -12, -9, 5, 26, 7, 24, 14, -36, 18,
    -- layer=1 filter=252 channel=10
    -29, -22, 16, -29, -5, -1, 11, 24, 10,
    -- layer=1 filter=252 channel=11
    -10, -13, 10, -20, -56, -11, -12, -26, 2,
    -- layer=1 filter=252 channel=12
    -18, -10, -18, 26, 21, 22, -14, 5, -8,
    -- layer=1 filter=252 channel=13
    0, 6, -8, 18, 33, 16, 4, 12, 8,
    -- layer=1 filter=252 channel=14
    -15, -22, 9, -66, -39, -15, -29, -20, -34,
    -- layer=1 filter=252 channel=15
    -52, -45, -47, -69, -73, -58, -20, 1, 35,
    -- layer=1 filter=252 channel=16
    2, 19, 16, -71, -71, -69, 0, -20, -20,
    -- layer=1 filter=252 channel=17
    -2, -27, 10, -21, -19, -12, -42, -44, -47,
    -- layer=1 filter=252 channel=18
    -2, 25, 27, -14, -35, -26, -8, 0, -8,
    -- layer=1 filter=252 channel=19
    -53, -15, -29, -25, -25, -16, 10, -24, 4,
    -- layer=1 filter=252 channel=20
    -1, 9, 4, 28, 29, 21, 19, 13, 0,
    -- layer=1 filter=252 channel=21
    -3, -3, 4, 13, 24, 2, 13, 14, 7,
    -- layer=1 filter=252 channel=22
    -3, 10, -10, 11, 25, 20, 4, -1, -23,
    -- layer=1 filter=252 channel=23
    -4, 7, -27, -57, -64, 0, -36, -62, 0,
    -- layer=1 filter=252 channel=24
    -6, 17, -1, -10, -27, -4, -6, -13, -12,
    -- layer=1 filter=252 channel=25
    -33, -21, 3, -51, -19, -3, -9, -7, 6,
    -- layer=1 filter=252 channel=26
    -6, 16, 17, 2, 3, 11, -5, 1, -4,
    -- layer=1 filter=252 channel=27
    -2, -4, 0, -12, -10, -30, 10, -11, -14,
    -- layer=1 filter=252 channel=28
    -5, 35, 35, -23, 33, 16, -41, 8, 4,
    -- layer=1 filter=252 channel=29
    -39, -39, -37, -23, -19, -11, -25, -5, -12,
    -- layer=1 filter=252 channel=30
    -13, 3, 22, -15, -16, -6, 14, 10, -2,
    -- layer=1 filter=252 channel=31
    20, 9, 2, 16, 20, 18, 38, 41, 20,
    -- layer=1 filter=252 channel=32
    -44, -6, 8, -22, -13, 8, 0, -8, 14,
    -- layer=1 filter=252 channel=33
    -27, -29, -4, -12, -5, -18, 6, -15, -7,
    -- layer=1 filter=252 channel=34
    -56, -63, -53, -38, -49, -45, -37, -31, -29,
    -- layer=1 filter=252 channel=35
    0, 7, 23, -21, -6, -4, 16, 13, 32,
    -- layer=1 filter=252 channel=36
    6, 8, 14, -24, -51, -19, 1, -25, 14,
    -- layer=1 filter=252 channel=37
    -66, -48, -25, -141, -128, -82, 56, 54, 61,
    -- layer=1 filter=252 channel=38
    -11, 4, -13, 16, 36, 21, 24, 30, 19,
    -- layer=1 filter=252 channel=39
    2, 14, 5, -11, -23, -8, -8, -10, -23,
    -- layer=1 filter=252 channel=40
    26, 26, 16, 47, 48, 39, 54, 53, 44,
    -- layer=1 filter=252 channel=41
    -29, 9, 18, -16, -42, -10, -29, -52, 14,
    -- layer=1 filter=252 channel=42
    13, 5, 9, 34, 21, 31, 30, 7, 12,
    -- layer=1 filter=252 channel=43
    0, 13, 15, -43, -61, -70, -22, -11, -51,
    -- layer=1 filter=252 channel=44
    -35, 10, 23, -22, -19, 6, -4, -9, 2,
    -- layer=1 filter=252 channel=45
    -16, -1, -1, -10, -13, -2, 13, 21, 0,
    -- layer=1 filter=252 channel=46
    -56, -57, -18, -41, -31, -27, 39, 33, 42,
    -- layer=1 filter=252 channel=47
    -45, -8, -7, -50, -14, 50, 10, 20, 62,
    -- layer=1 filter=252 channel=48
    1, -6, -10, 14, 12, 4, -14, 13, -8,
    -- layer=1 filter=252 channel=49
    -2, -20, -18, 19, 10, 11, 37, 20, 20,
    -- layer=1 filter=252 channel=50
    -8, -8, -24, 6, 17, 16, -10, -31, -24,
    -- layer=1 filter=252 channel=51
    -7, 10, -6, 12, 28, 2, 22, 31, 18,
    -- layer=1 filter=252 channel=52
    2, 0, 0, 1, -16, -22, -28, -6, -2,
    -- layer=1 filter=252 channel=53
    14, 2, -12, 0, 1, -18, -4, 1, 2,
    -- layer=1 filter=252 channel=54
    -51, -68, -19, -64, -67, -34, 17, 8, 15,
    -- layer=1 filter=252 channel=55
    12, 2, 34, -44, -50, -15, -25, -26, -6,
    -- layer=1 filter=252 channel=56
    -8, 0, 0, -5, 1, 4, -1, 1, -6,
    -- layer=1 filter=252 channel=57
    -2, 14, 22, -5, 33, 24, 18, 40, 40,
    -- layer=1 filter=252 channel=58
    -16, -29, -17, -63, -27, -24, 29, 9, 0,
    -- layer=1 filter=252 channel=59
    -10, 0, -2, -14, -2, -5, -16, -10, -11,
    -- layer=1 filter=252 channel=60
    0, -2, -14, -6, 11, 0, 8, -6, -3,
    -- layer=1 filter=252 channel=61
    -4, 15, 0, 6, -4, -7, 16, -4, 3,
    -- layer=1 filter=252 channel=62
    -1, -2, -1, -100, -94, -62, -10, -23, -33,
    -- layer=1 filter=252 channel=63
    -21, 3, 7, -46, -59, -44, -23, -54, -15,
    -- layer=1 filter=252 channel=64
    -11, -14, -5, -18, 1, -12, -20, 0, -14,
    -- layer=1 filter=252 channel=65
    -3, 21, 10, 7, 25, 3, -7, 0, -7,
    -- layer=1 filter=252 channel=66
    -1, -24, 0, -40, -43, -20, -2, -6, -17,
    -- layer=1 filter=252 channel=67
    -7, -18, -8, 23, 56, 9, 6, 12, 8,
    -- layer=1 filter=252 channel=68
    -37, 0, 10, -13, -36, 3, -18, -8, 3,
    -- layer=1 filter=252 channel=69
    2, 14, 9, -61, -79, -50, -1, 1, 20,
    -- layer=1 filter=252 channel=70
    2, -45, -9, 8, 12, 24, 55, 52, 26,
    -- layer=1 filter=252 channel=71
    -9, -20, -9, -16, -20, -39, -14, -23, -24,
    -- layer=1 filter=252 channel=72
    -1, 12, 18, 11, -17, 11, -10, -32, -26,
    -- layer=1 filter=252 channel=73
    -12, -9, -12, -6, 0, 0, -12, -14, -10,
    -- layer=1 filter=252 channel=74
    9, -1, 32, 5, 5, 8, 19, 20, 21,
    -- layer=1 filter=252 channel=75
    -3, -13, 21, -11, -27, 2, -32, -19, -34,
    -- layer=1 filter=252 channel=76
    -6, 16, 24, 4, -20, 1, -15, -25, -18,
    -- layer=1 filter=252 channel=77
    -15, 6, -1, -20, -5, -1, -4, 2, -1,
    -- layer=1 filter=252 channel=78
    -8, 9, 19, -11, 17, 5, -3, 21, 14,
    -- layer=1 filter=252 channel=79
    10, 17, 8, -55, -61, -38, -4, -12, -34,
    -- layer=1 filter=252 channel=80
    -11, -9, -4, -28, -8, -21, 0, -27, -7,
    -- layer=1 filter=252 channel=81
    3, 32, 27, -26, -45, -15, -33, -44, -33,
    -- layer=1 filter=252 channel=82
    -5, 6, -7, 14, 24, 10, 8, 5, 6,
    -- layer=1 filter=252 channel=83
    -2, 14, -2, -32, -59, -8, -29, -17, -28,
    -- layer=1 filter=252 channel=84
    16, 18, 35, 0, -9, 6, -5, -6, -7,
    -- layer=1 filter=252 channel=85
    -28, -15, -35, -51, -29, 0, -6, -21, 5,
    -- layer=1 filter=252 channel=86
    4, 0, 9, -10, -32, -7, 3, -20, -9,
    -- layer=1 filter=252 channel=87
    11, 5, 15, 1, 12, 21, 78, 13, 58,
    -- layer=1 filter=252 channel=88
    1, -8, -23, 12, 14, -12, 6, 17, -16,
    -- layer=1 filter=252 channel=89
    1, 13, 3, 7, 23, 0, 9, 4, 2,
    -- layer=1 filter=252 channel=90
    -48, -10, 0, -67, -51, 1, -30, -46, 5,
    -- layer=1 filter=252 channel=91
    -5, 17, 13, 31, 35, 32, 22, 38, 29,
    -- layer=1 filter=252 channel=92
    -17, 7, 8, -34, -66, 0, -50, -51, 22,
    -- layer=1 filter=252 channel=93
    1, -2, -2, -9, -11, -20, -6, -12, -25,
    -- layer=1 filter=252 channel=94
    7, 0, 27, -11, -8, 0, -35, -17, 4,
    -- layer=1 filter=252 channel=95
    2, -6, 29, -24, -32, -23, -9, -3, -4,
    -- layer=1 filter=252 channel=96
    -25, -24, -17, -19, -15, -25, -14, -3, -17,
    -- layer=1 filter=252 channel=97
    13, 4, 14, -16, -19, -11, -45, -42, -20,
    -- layer=1 filter=252 channel=98
    8, 13, 15, -34, -31, -21, -18, -28, -46,
    -- layer=1 filter=252 channel=99
    -23, -4, 28, -6, 3, -21, -1, -2, 21,
    -- layer=1 filter=252 channel=100
    -19, -5, 0, -42, -46, -17, -14, -35, -18,
    -- layer=1 filter=252 channel=101
    4, 8, -5, 23, 20, 28, 26, 30, 10,
    -- layer=1 filter=252 channel=102
    0, -5, 10, -2, 8, 9, -24, -24, -10,
    -- layer=1 filter=252 channel=103
    -17, -26, -9, -34, -29, -37, -13, -21, -20,
    -- layer=1 filter=252 channel=104
    11, 17, -7, -30, -22, -10, -17, -18, -5,
    -- layer=1 filter=252 channel=105
    -11, -2, 8, -21, -35, -21, -37, -45, -11,
    -- layer=1 filter=252 channel=106
    -5, -5, -9, 32, 18, 27, 29, 26, 20,
    -- layer=1 filter=252 channel=107
    -1, 9, 10, 8, -8, 12, -4, 16, -6,
    -- layer=1 filter=252 channel=108
    -17, 0, -3, -20, -37, -8, -17, -17, -14,
    -- layer=1 filter=252 channel=109
    4, 1, 7, -3, -3, 9, -8, -10, 8,
    -- layer=1 filter=252 channel=110
    -1, 9, 0, 2, 10, 0, -9, -8, 5,
    -- layer=1 filter=252 channel=111
    -1, 15, 32, -13, -19, -6, 12, 4, -1,
    -- layer=1 filter=252 channel=112
    -22, -4, 36, -30, -66, -27, -25, -10, -4,
    -- layer=1 filter=252 channel=113
    -38, -59, -42, -6, -7, -30, 29, 28, 0,
    -- layer=1 filter=252 channel=114
    11, 22, 20, -47, -54, -48, 33, 61, 33,
    -- layer=1 filter=252 channel=115
    9, 13, 31, -21, -14, -12, -5, -32, -15,
    -- layer=1 filter=252 channel=116
    -3, -6, -5, -3, -5, 8, -1, 0, 3,
    -- layer=1 filter=252 channel=117
    -14, 3, 21, -28, -60, -46, -31, -35, -56,
    -- layer=1 filter=252 channel=118
    3, 23, 37, 3, 0, 11, 30, 41, 30,
    -- layer=1 filter=252 channel=119
    -65, -16, -8, -46, -44, -8, -46, -28, -15,
    -- layer=1 filter=252 channel=120
    -14, -7, -4, 0, 15, 2, 3, 6, 3,
    -- layer=1 filter=252 channel=121
    27, -7, 29, -30, -21, -18, -9, -43, -11,
    -- layer=1 filter=252 channel=122
    -2, -6, -8, -6, 3, -9, 0, -3, -3,
    -- layer=1 filter=252 channel=123
    15, -26, 14, -60, -69, -28, -9, -36, -36,
    -- layer=1 filter=252 channel=124
    -9, -7, 9, -12, 2, -10, 1, -8, -2,
    -- layer=1 filter=252 channel=125
    -30, -47, -50, -10, 15, -11, 57, 43, 35,
    -- layer=1 filter=252 channel=126
    -14, -9, 16, -73, -62, -33, -45, -36, -45,
    -- layer=1 filter=252 channel=127
    18, 27, 44, -10, -18, 6, 15, 27, 11,
    -- layer=1 filter=253 channel=0
    17, 11, 0, 3, 4, -1, 8, 0, -5,
    -- layer=1 filter=253 channel=1
    6, 8, 38, -20, -22, 11, -4, -12, -12,
    -- layer=1 filter=253 channel=2
    17, 26, -13, 14, 37, 24, 20, 32, 22,
    -- layer=1 filter=253 channel=3
    4, 9, 0, -5, -7, 9, 1, 11, -9,
    -- layer=1 filter=253 channel=4
    -3, 0, 1, 4, 1, 8, 6, -3, 3,
    -- layer=1 filter=253 channel=5
    -12, -4, -3, -45, -41, -4, -40, -46, -48,
    -- layer=1 filter=253 channel=6
    -11, 2, 23, 12, 15, 22, 30, 39, 10,
    -- layer=1 filter=253 channel=7
    4, 42, 65, -1, 51, 21, 19, 50, 5,
    -- layer=1 filter=253 channel=8
    15, 14, 41, -8, -24, -13, -20, -47, -41,
    -- layer=1 filter=253 channel=9
    -32, -13, -42, -26, 3, -24, -25, 1, -24,
    -- layer=1 filter=253 channel=10
    -20, 27, 46, -9, 16, 17, 1, 30, 1,
    -- layer=1 filter=253 channel=11
    35, 15, 7, 28, 1, -17, 13, -7, 2,
    -- layer=1 filter=253 channel=12
    39, -15, 46, 8, -27, 77, -8, -4, -7,
    -- layer=1 filter=253 channel=13
    6, 24, 12, 10, 22, 14, 3, 17, 6,
    -- layer=1 filter=253 channel=14
    -28, 7, 55, -40, -24, -7, -33, -17, -38,
    -- layer=1 filter=253 channel=15
    -20, 28, -40, -15, -22, 0, -37, 7, -17,
    -- layer=1 filter=253 channel=16
    -18, -27, -2, -34, -37, -9, -26, -50, -46,
    -- layer=1 filter=253 channel=17
    23, 7, 20, 26, 29, 9, 20, 11, 21,
    -- layer=1 filter=253 channel=18
    9, -13, 34, -35, -37, -27, 11, -6, -18,
    -- layer=1 filter=253 channel=19
    -56, -61, -64, -79, -34, -50, -39, -48, -46,
    -- layer=1 filter=253 channel=20
    1, 12, 7, 16, 17, 6, 12, 19, 18,
    -- layer=1 filter=253 channel=21
    -11, -16, 8, -27, -22, -8, -18, 0, -21,
    -- layer=1 filter=253 channel=22
    -1, 22, 39, 7, 7, 25, 11, 32, 11,
    -- layer=1 filter=253 channel=23
    -24, -16, -15, 28, 24, 0, 21, 55, 7,
    -- layer=1 filter=253 channel=24
    -12, -18, -19, -43, -7, -38, -35, -45, -29,
    -- layer=1 filter=253 channel=25
    -19, -3, 28, 0, 3, 3, 5, 10, -23,
    -- layer=1 filter=253 channel=26
    13, 38, 8, 21, 36, 0, 31, 26, -7,
    -- layer=1 filter=253 channel=27
    52, 38, 13, 38, 28, -1, 18, -2, -13,
    -- layer=1 filter=253 channel=28
    -43, 10, 32, -14, 23, 15, -1, 35, 4,
    -- layer=1 filter=253 channel=29
    29, -2, -17, 20, -10, -19, 0, -10, -32,
    -- layer=1 filter=253 channel=30
    -14, -56, -2, -68, -57, -51, -21, -42, -21,
    -- layer=1 filter=253 channel=31
    -15, -7, 18, -28, -19, -9, 9, 21, 2,
    -- layer=1 filter=253 channel=32
    5, 8, 8, 0, 29, 18, 27, 35, -1,
    -- layer=1 filter=253 channel=33
    0, -14, 3, 8, -16, -5, 32, 26, 34,
    -- layer=1 filter=253 channel=34
    -58, -35, -36, -54, -57, -54, -26, -18, -33,
    -- layer=1 filter=253 channel=35
    -4, 2, 4, -2, -12, -9, -16, -8, -20,
    -- layer=1 filter=253 channel=36
    48, 17, 3, 34, 4, 5, 29, 14, 2,
    -- layer=1 filter=253 channel=37
    -41, -38, -19, -61, -48, 6, -62, -58, -43,
    -- layer=1 filter=253 channel=38
    0, 2, 12, -2, 22, 1, 13, 6, 17,
    -- layer=1 filter=253 channel=39
    28, 3, 8, 31, 5, 12, 21, 6, 10,
    -- layer=1 filter=253 channel=40
    -16, -2, 34, 17, 19, 31, 29, 40, 30,
    -- layer=1 filter=253 channel=41
    -14, -28, -16, -16, -18, -35, -7, 0, -45,
    -- layer=1 filter=253 channel=42
    54, 15, 20, 56, 26, 35, 41, 29, 23,
    -- layer=1 filter=253 channel=43
    1, -20, 29, -35, -46, -24, -33, -41, -76,
    -- layer=1 filter=253 channel=44
    35, 46, 22, 24, 40, 15, 46, 26, -5,
    -- layer=1 filter=253 channel=45
    -3, 12, -15, 7, -5, 9, 3, -9, -22,
    -- layer=1 filter=253 channel=46
    -64, -85, -72, -63, -12, 22, -13, -19, 26,
    -- layer=1 filter=253 channel=47
    -50, 0, -20, -17, 32, 7, 0, 58, 2,
    -- layer=1 filter=253 channel=48
    -8, -3, -7, -3, -1, -2, 0, 5, -3,
    -- layer=1 filter=253 channel=49
    -18, -1, -12, -7, -6, -4, 6, 12, 0,
    -- layer=1 filter=253 channel=50
    9, 12, 12, 16, 17, 10, 13, 17, 0,
    -- layer=1 filter=253 channel=51
    -19, -2, 11, -4, -8, 2, -8, 4, -5,
    -- layer=1 filter=253 channel=52
    -2, 7, -10, 1, 3, 3, 0, -1, -12,
    -- layer=1 filter=253 channel=53
    4, -11, 10, 14, -12, 7, 10, -22, 1,
    -- layer=1 filter=253 channel=54
    -37, -8, 7, -39, -5, -25, -16, -18, -60,
    -- layer=1 filter=253 channel=55
    9, -5, -25, 8, -7, -5, -1, -16, -20,
    -- layer=1 filter=253 channel=56
    10, 0, -1, -8, -9, -5, -7, 3, 1,
    -- layer=1 filter=253 channel=57
    -20, 21, 17, 0, 24, 1, 19, 31, 19,
    -- layer=1 filter=253 channel=58
    -17, 17, 11, 2, 19, -28, 45, 53, -5,
    -- layer=1 filter=253 channel=59
    -10, 0, 2, 0, 3, 5, 1, -13, -6,
    -- layer=1 filter=253 channel=60
    0, 2, -4, 0, 6, -5, 6, 5, 2,
    -- layer=1 filter=253 channel=61
    0, -8, -2, 10, -11, 0, 3, 10, -9,
    -- layer=1 filter=253 channel=62
    -17, -10, 0, -52, -38, -17, -38, -48, -64,
    -- layer=1 filter=253 channel=63
    29, 0, 4, 15, -5, -15, 0, 0, -18,
    -- layer=1 filter=253 channel=64
    12, 1, 5, -11, 8, 8, 5, 10, 6,
    -- layer=1 filter=253 channel=65
    -11, 0, -6, -1, -2, -12, -3, -2, -5,
    -- layer=1 filter=253 channel=66
    21, 8, -5, 11, -6, -12, 0, -11, -7,
    -- layer=1 filter=253 channel=67
    -41, -26, -24, -61, -46, -44, -72, -56, -65,
    -- layer=1 filter=253 channel=68
    35, 54, 34, 53, 39, 16, 59, 27, 8,
    -- layer=1 filter=253 channel=69
    0, 9, -6, -28, -13, 0, -47, -4, -19,
    -- layer=1 filter=253 channel=70
    -26, -14, -17, -24, -25, -12, -15, -19, -8,
    -- layer=1 filter=253 channel=71
    -16, -32, -34, -17, -35, -40, -41, -56, -52,
    -- layer=1 filter=253 channel=72
    35, -19, 25, -31, -19, -25, -20, -2, -18,
    -- layer=1 filter=253 channel=73
    -2, -11, 0, -5, -12, -10, -6, 3, 1,
    -- layer=1 filter=253 channel=74
    9, -6, 14, 7, -5, -24, 36, 18, -17,
    -- layer=1 filter=253 channel=75
    5, -16, 22, -61, -24, 7, -51, -32, -44,
    -- layer=1 filter=253 channel=76
    18, -2, 6, 15, 0, -16, 28, -12, -19,
    -- layer=1 filter=253 channel=77
    -5, -17, -7, -11, -4, 1, -12, -26, -3,
    -- layer=1 filter=253 channel=78
    0, 18, 6, -7, 9, -14, -4, 0, -15,
    -- layer=1 filter=253 channel=79
    -9, 8, -2, -31, -9, -14, -17, -20, -28,
    -- layer=1 filter=253 channel=80
    7, 3, 2, 14, -10, -3, 3, -3, 4,
    -- layer=1 filter=253 channel=81
    -12, -20, -15, -27, -31, -35, -36, -54, -36,
    -- layer=1 filter=253 channel=82
    -12, 0, -1, -15, -8, 2, -26, -5, -2,
    -- layer=1 filter=253 channel=83
    11, 25, -6, -6, -24, 15, 10, -13, -13,
    -- layer=1 filter=253 channel=84
    -3, -15, 26, 4, 6, -13, 44, -4, -19,
    -- layer=1 filter=253 channel=85
    -14, 0, -4, -3, 17, -14, 22, 68, -35,
    -- layer=1 filter=253 channel=86
    20, 1, 3, 23, 5, -5, 6, 1, -9,
    -- layer=1 filter=253 channel=87
    -25, -13, -43, -47, -8, -1, -18, 3, -19,
    -- layer=1 filter=253 channel=88
    -1, -6, -6, -9, -5, -4, -5, -14, -18,
    -- layer=1 filter=253 channel=89
    -23, -16, -10, -8, -11, -1, -6, -15, -18,
    -- layer=1 filter=253 channel=90
    43, 29, 25, 24, 41, 20, 38, 16, 5,
    -- layer=1 filter=253 channel=91
    -11, 3, 11, 6, 21, 20, 4, 11, 11,
    -- layer=1 filter=253 channel=92
    -23, -25, -18, 10, -45, -17, -22, -27, -34,
    -- layer=1 filter=253 channel=93
    -16, -16, -8, -19, -24, -19, -13, -20, -9,
    -- layer=1 filter=253 channel=94
    18, 21, -3, 14, 14, 0, 18, 13, -4,
    -- layer=1 filter=253 channel=95
    -7, -6, 8, -24, -27, -15, 15, -20, -40,
    -- layer=1 filter=253 channel=96
    -6, -1, -7, 5, 5, 6, -4, 0, 6,
    -- layer=1 filter=253 channel=97
    23, 3, -5, 9, -3, 5, -1, -10, -10,
    -- layer=1 filter=253 channel=98
    17, 13, 50, -29, -7, 5, -12, -21, -35,
    -- layer=1 filter=253 channel=99
    -39, -2, -3, -2, 18, 25, 15, 10, 26,
    -- layer=1 filter=253 channel=100
    23, 3, 2, 22, -5, -3, 17, -13, -1,
    -- layer=1 filter=253 channel=101
    -17, -3, 11, 11, 11, 18, 6, 4, 11,
    -- layer=1 filter=253 channel=102
    24, 10, 14, 18, 16, 14, 19, 21, 9,
    -- layer=1 filter=253 channel=103
    11, 0, 10, 1, 6, -7, 2, -13, -5,
    -- layer=1 filter=253 channel=104
    -4, 1, -31, 5, 4, -18, -8, 19, -21,
    -- layer=1 filter=253 channel=105
    2, 7, -1, 15, 1, -4, -3, -13, 4,
    -- layer=1 filter=253 channel=106
    -9, 19, 4, 12, 30, 10, 21, 35, 2,
    -- layer=1 filter=253 channel=107
    0, -6, 0, 1, -1, 13, -1, -8, 7,
    -- layer=1 filter=253 channel=108
    6, 24, 21, 30, 42, 4, 24, 47, -15,
    -- layer=1 filter=253 channel=109
    1, 6, -8, 4, -5, 4, -9, -10, 5,
    -- layer=1 filter=253 channel=110
    11, -3, 1, 6, 0, -15, -2, -9, 0,
    -- layer=1 filter=253 channel=111
    -10, -21, 8, -30, -19, -28, 1, -20, -38,
    -- layer=1 filter=253 channel=112
    -46, 4, 0, 9, -26, 0, 2, -28, -48,
    -- layer=1 filter=253 channel=113
    -27, -8, -4, -7, -27, -5, 14, 7, 11,
    -- layer=1 filter=253 channel=114
    -4, 7, -16, 20, -32, 10, -33, -57, -13,
    -- layer=1 filter=253 channel=115
    -4, 4, 3, -1, -1, 3, 0, 12, -3,
    -- layer=1 filter=253 channel=116
    6, 4, -2, 11, 7, 0, 7, 4, 7,
    -- layer=1 filter=253 channel=117
    -77, -2, -9, -56, -66, -16, -31, -43, -34,
    -- layer=1 filter=253 channel=118
    4, -15, 8, -1, -12, -22, 15, 0, -3,
    -- layer=1 filter=253 channel=119
    14, 21, 14, 19, 38, 14, 24, 19, -6,
    -- layer=1 filter=253 channel=120
    -12, -2, 20, -9, 5, -7, -13, 3, -7,
    -- layer=1 filter=253 channel=121
    16, -22, 2, -46, -21, -9, -51, -67, -29,
    -- layer=1 filter=253 channel=122
    7, -2, 10, 1, 9, 3, 5, 0, 3,
    -- layer=1 filter=253 channel=123
    34, -9, -4, -17, -16, -31, -31, -50, -30,
    -- layer=1 filter=253 channel=124
    3, -4, -6, 0, 0, -4, -2, -10, -4,
    -- layer=1 filter=253 channel=125
    -24, -22, -10, -21, -26, -29, 11, 1, -11,
    -- layer=1 filter=253 channel=126
    -14, 6, 25, -67, -36, -16, -47, -27, -13,
    -- layer=1 filter=253 channel=127
    -4, -23, 18, -23, -37, -29, -4, -14, -39,
    -- layer=1 filter=254 channel=0
    -3, -2, 4, -7, 1, 1, 0, -8, -4,
    -- layer=1 filter=254 channel=1
    -2, 4, 3, 4, 1, 1, -10, 3, -12,
    -- layer=1 filter=254 channel=2
    -16, -6, 1, -16, 0, -9, 3, -10, -14,
    -- layer=1 filter=254 channel=3
    4, 7, -7, 2, 0, 0, 8, 7, 3,
    -- layer=1 filter=254 channel=4
    7, 5, 4, -1, -6, -5, -2, 2, 6,
    -- layer=1 filter=254 channel=5
    9, -5, 2, -18, -4, -6, 0, -7, 0,
    -- layer=1 filter=254 channel=6
    1, -10, -5, 5, -13, 3, -3, 4, -5,
    -- layer=1 filter=254 channel=7
    -3, 0, -13, -4, -16, -17, 4, -5, -2,
    -- layer=1 filter=254 channel=8
    -7, 6, 2, -16, -9, -5, 1, 2, -14,
    -- layer=1 filter=254 channel=9
    -18, 8, -1, 5, 3, 3, -6, -1, -1,
    -- layer=1 filter=254 channel=10
    3, -14, -2, -10, -13, -6, 5, -4, -4,
    -- layer=1 filter=254 channel=11
    -9, -3, -7, 1, -5, -4, 3, -4, 3,
    -- layer=1 filter=254 channel=12
    -7, -6, 1, -13, -9, -7, -8, -6, -2,
    -- layer=1 filter=254 channel=13
    -9, -4, -15, -10, -12, -7, 0, -4, -5,
    -- layer=1 filter=254 channel=14
    -10, -2, -16, -5, -13, -10, 0, -11, -5,
    -- layer=1 filter=254 channel=15
    -8, 9, 0, -17, -10, -8, -7, -2, -1,
    -- layer=1 filter=254 channel=16
    6, -1, -4, -17, -13, -12, -2, -1, -1,
    -- layer=1 filter=254 channel=17
    -8, 3, -12, -6, -4, -4, -1, -5, -11,
    -- layer=1 filter=254 channel=18
    -5, -8, -3, -11, -8, -10, -4, 4, -12,
    -- layer=1 filter=254 channel=19
    -16, -4, -3, 0, 0, -12, 2, -6, -2,
    -- layer=1 filter=254 channel=20
    6, 5, 5, -1, 1, 1, -9, -10, -10,
    -- layer=1 filter=254 channel=21
    -8, -3, -5, -13, -17, -13, -12, -13, -11,
    -- layer=1 filter=254 channel=22
    -9, -1, 1, -6, -6, -10, -15, -7, 0,
    -- layer=1 filter=254 channel=23
    -13, 8, -5, -11, -1, -14, -8, 4, 0,
    -- layer=1 filter=254 channel=24
    -7, -14, 0, -8, -4, -15, -1, 0, -1,
    -- layer=1 filter=254 channel=25
    -16, -5, 2, -19, 0, 0, -15, -10, -14,
    -- layer=1 filter=254 channel=26
    7, -11, -13, 0, -12, -3, -2, -2, -14,
    -- layer=1 filter=254 channel=27
    -7, 6, -8, 0, -14, -5, 3, -4, -7,
    -- layer=1 filter=254 channel=28
    1, 3, -5, -11, -13, 5, -7, 3, -3,
    -- layer=1 filter=254 channel=29
    4, 5, 9, 0, 3, -3, 1, -6, -9,
    -- layer=1 filter=254 channel=30
    -13, 2, 0, 4, -6, -17, -9, 1, 2,
    -- layer=1 filter=254 channel=31
    -7, -11, 3, 0, -4, -17, -15, 3, -16,
    -- layer=1 filter=254 channel=32
    -8, 6, -3, -9, 4, 1, 0, -1, 4,
    -- layer=1 filter=254 channel=33
    -1, -8, -5, 0, -4, 2, -2, 3, 0,
    -- layer=1 filter=254 channel=34
    -7, 3, -11, 1, 5, 6, -3, 0, -6,
    -- layer=1 filter=254 channel=35
    -2, 3, -2, 5, -1, 3, -6, -7, 1,
    -- layer=1 filter=254 channel=36
    -5, -16, -17, 7, 2, 3, -11, -2, -5,
    -- layer=1 filter=254 channel=37
    -1, -2, 4, 1, -8, 1, -10, 0, -17,
    -- layer=1 filter=254 channel=38
    -13, -16, 2, -15, -5, -16, -4, -11, -11,
    -- layer=1 filter=254 channel=39
    1, -8, 5, 6, 1, 3, 3, -11, 0,
    -- layer=1 filter=254 channel=40
    2, -5, -8, -10, -7, -5, -8, -13, -15,
    -- layer=1 filter=254 channel=41
    -7, 0, -3, -2, -5, -8, -3, -2, -16,
    -- layer=1 filter=254 channel=42
    3, -6, -2, -4, -15, 0, 2, -1, -10,
    -- layer=1 filter=254 channel=43
    8, -10, 3, -14, 0, -6, -1, -8, -5,
    -- layer=1 filter=254 channel=44
    -6, -2, -9, 3, -2, 0, -1, -10, -3,
    -- layer=1 filter=254 channel=45
    6, -1, -7, -9, 1, -11, -4, -16, -10,
    -- layer=1 filter=254 channel=46
    -4, 0, 0, -6, -17, -12, -12, -15, -11,
    -- layer=1 filter=254 channel=47
    -16, 6, -11, 0, -1, 0, -6, -6, -6,
    -- layer=1 filter=254 channel=48
    -2, 1, 0, -2, -8, -3, -2, -11, -5,
    -- layer=1 filter=254 channel=49
    5, -9, 2, 4, -7, 0, 1, -11, -4,
    -- layer=1 filter=254 channel=50
    -9, -5, -3, -11, 5, 0, 0, -4, -6,
    -- layer=1 filter=254 channel=51
    -6, -2, -14, -2, -3, -15, -4, -11, -7,
    -- layer=1 filter=254 channel=52
    4, 8, -4, -9, -9, 7, 3, 5, -8,
    -- layer=1 filter=254 channel=53
    -6, -7, -1, 0, -5, -5, -3, -10, -8,
    -- layer=1 filter=254 channel=54
    0, 0, -2, -15, -12, -12, -6, -4, -14,
    -- layer=1 filter=254 channel=55
    -17, -15, -12, -5, -7, -15, 0, -1, -9,
    -- layer=1 filter=254 channel=56
    6, -6, 4, 6, -11, 4, -11, -10, 3,
    -- layer=1 filter=254 channel=57
    -15, -9, -7, -2, -2, -15, -14, -1, -13,
    -- layer=1 filter=254 channel=58
    -6, -14, -18, -7, -10, 2, 5, -9, -11,
    -- layer=1 filter=254 channel=59
    2, -12, 3, 6, -5, 7, -8, 1, 4,
    -- layer=1 filter=254 channel=60
    -1, 3, 7, -2, -7, -6, 0, -9, -5,
    -- layer=1 filter=254 channel=61
    -8, -5, 9, 4, 0, 5, 10, 8, -9,
    -- layer=1 filter=254 channel=62
    6, -4, 1, -11, 0, -3, -7, -9, -17,
    -- layer=1 filter=254 channel=63
    -5, -6, -10, 6, 6, -13, -11, -10, -1,
    -- layer=1 filter=254 channel=64
    -5, -3, 5, -11, -10, 3, 0, -9, 4,
    -- layer=1 filter=254 channel=65
    -14, 0, 0, 8, 1, -11, -9, 0, 6,
    -- layer=1 filter=254 channel=66
    0, -12, 3, -1, 0, -11, -7, 3, 6,
    -- layer=1 filter=254 channel=67
    0, -10, -10, -2, 9, 4, 7, 5, 0,
    -- layer=1 filter=254 channel=68
    5, -13, 3, 0, -6, -14, -13, -8, -5,
    -- layer=1 filter=254 channel=69
    4, -1, -10, -1, -14, -9, -13, -3, -8,
    -- layer=1 filter=254 channel=70
    -8, -2, 1, 6, -9, -5, -7, 2, -14,
    -- layer=1 filter=254 channel=71
    -6, -8, -12, -1, -7, -16, -13, -11, -10,
    -- layer=1 filter=254 channel=72
    -5, 8, -2, 9, 4, -10, 5, 0, -2,
    -- layer=1 filter=254 channel=73
    8, -10, -7, -7, 2, -11, -7, -7, -3,
    -- layer=1 filter=254 channel=74
    -1, -1, -15, 5, -3, 7, 0, -1, -10,
    -- layer=1 filter=254 channel=75
    2, 0, 0, -9, -9, -16, -8, -17, -2,
    -- layer=1 filter=254 channel=76
    -7, -4, -2, -10, -5, 2, -6, 5, 9,
    -- layer=1 filter=254 channel=77
    5, -7, 0, 0, 4, 7, 1, 1, 3,
    -- layer=1 filter=254 channel=78
    -4, -9, -7, -3, -3, 8, -8, -5, 0,
    -- layer=1 filter=254 channel=79
    -3, 5, 6, -4, 7, -14, -7, -9, 0,
    -- layer=1 filter=254 channel=80
    2, 8, 8, -7, -9, 4, 0, 3, 3,
    -- layer=1 filter=254 channel=81
    -2, -2, 3, -11, -5, -10, -2, -14, -14,
    -- layer=1 filter=254 channel=82
    -14, -6, -10, -7, -14, -1, -11, -2, -11,
    -- layer=1 filter=254 channel=83
    -5, 4, 8, -8, 3, -7, -7, 3, 0,
    -- layer=1 filter=254 channel=84
    0, -10, -9, -5, -4, -9, -5, -9, -8,
    -- layer=1 filter=254 channel=85
    -9, -11, 0, -11, 4, -8, 8, 5, -8,
    -- layer=1 filter=254 channel=86
    -6, -3, -6, 6, -8, 0, 1, -2, -8,
    -- layer=1 filter=254 channel=87
    -10, 1, -8, -9, -7, 0, -15, -3, -4,
    -- layer=1 filter=254 channel=88
    -8, 4, 10, -3, -14, -6, 3, -14, -8,
    -- layer=1 filter=254 channel=89
    2, -4, -9, 1, -13, -5, 2, -14, 0,
    -- layer=1 filter=254 channel=90
    -1, 1, -10, -4, -8, -4, -5, -10, -9,
    -- layer=1 filter=254 channel=91
    -5, 0, -3, -9, -4, -4, -5, -16, -2,
    -- layer=1 filter=254 channel=92
    1, -2, 0, -14, -14, 0, 1, -17, -6,
    -- layer=1 filter=254 channel=93
    1, 0, -9, -10, -8, -1, -18, -8, -10,
    -- layer=1 filter=254 channel=94
    2, 0, 0, 0, -4, -10, 5, -3, 5,
    -- layer=1 filter=254 channel=95
    -8, -11, -9, -8, -12, 0, -12, 2, 6,
    -- layer=1 filter=254 channel=96
    -1, 3, -9, -7, 6, 4, -7, -11, 0,
    -- layer=1 filter=254 channel=97
    -5, -15, -4, -10, 2, 0, -13, -4, 0,
    -- layer=1 filter=254 channel=98
    -3, -11, -1, -13, -4, -16, -4, -18, -9,
    -- layer=1 filter=254 channel=99
    -7, -12, -7, 4, -3, -9, -1, 9, -6,
    -- layer=1 filter=254 channel=100
    -13, -11, -15, 4, -7, -5, -3, 4, 1,
    -- layer=1 filter=254 channel=101
    -16, -17, -18, -10, -7, -11, -19, -4, -12,
    -- layer=1 filter=254 channel=102
    -10, -15, -9, -7, 0, -4, -2, 3, -11,
    -- layer=1 filter=254 channel=103
    -8, -9, -7, -5, -6, -3, 5, -5, -3,
    -- layer=1 filter=254 channel=104
    -2, 5, -10, 8, 7, -10, -1, 4, -5,
    -- layer=1 filter=254 channel=105
    -11, -4, -9, -3, 3, 0, -8, -7, 5,
    -- layer=1 filter=254 channel=106
    1, -13, -1, -11, 0, -15, -13, 1, -6,
    -- layer=1 filter=254 channel=107
    -1, 3, -5, -3, -3, -1, 6, -9, 0,
    -- layer=1 filter=254 channel=108
    11, -8, 0, -8, -12, -1, -10, -13, -3,
    -- layer=1 filter=254 channel=109
    2, 0, 2, 1, 0, 2, -10, -6, -2,
    -- layer=1 filter=254 channel=110
    -3, -7, -7, 0, 8, 4, -5, -10, 4,
    -- layer=1 filter=254 channel=111
    1, 0, -7, 4, 5, 0, -5, 0, 3,
    -- layer=1 filter=254 channel=112
    -11, -14, 0, -8, 0, -5, -11, 5, 4,
    -- layer=1 filter=254 channel=113
    -13, -2, -6, -14, 3, -12, -4, -4, -4,
    -- layer=1 filter=254 channel=114
    9, 0, -8, -4, -10, -3, -1, -10, 0,
    -- layer=1 filter=254 channel=115
    -13, -3, -11, -1, 3, -5, 2, -5, -13,
    -- layer=1 filter=254 channel=116
    -7, -9, -6, 2, 7, 0, 7, 5, -2,
    -- layer=1 filter=254 channel=117
    -11, 1, -16, 5, -9, 0, -8, -12, 1,
    -- layer=1 filter=254 channel=118
    2, 2, -14, 0, -10, -7, -12, -8, 1,
    -- layer=1 filter=254 channel=119
    0, -5, -12, 12, 3, 8, -7, -11, 8,
    -- layer=1 filter=254 channel=120
    -11, -3, -10, -18, -11, 1, -2, -7, -3,
    -- layer=1 filter=254 channel=121
    -2, -5, 2, -8, -7, -4, -13, -13, -7,
    -- layer=1 filter=254 channel=122
    -2, -9, 9, -7, -5, -6, 9, -1, 9,
    -- layer=1 filter=254 channel=123
    0, -13, -1, -16, -16, 0, -17, -8, -1,
    -- layer=1 filter=254 channel=124
    7, -4, -7, -8, 3, 0, 8, -2, -2,
    -- layer=1 filter=254 channel=125
    3, 0, -7, 10, 5, 9, -2, -10, -4,
    -- layer=1 filter=254 channel=126
    6, -3, -9, 4, -2, 8, 7, 2, 5,
    -- layer=1 filter=254 channel=127
    -5, -3, 2, -12, -5, -8, -11, -9, -12,
    -- layer=1 filter=255 channel=0
    3, -4, -10, -10, -11, -7, -7, -7, 3,
    -- layer=1 filter=255 channel=1
    2, 0, -11, 6, 3, -4, 8, 7, -9,
    -- layer=1 filter=255 channel=2
    9, -8, -7, -9, -3, 4, 9, -2, -8,
    -- layer=1 filter=255 channel=3
    7, 8, 10, 8, -2, -10, 0, -7, 10,
    -- layer=1 filter=255 channel=4
    -4, -9, -3, 0, -1, 2, -7, -4, 4,
    -- layer=1 filter=255 channel=5
    0, -3, 5, 0, -3, -4, 6, 2, 4,
    -- layer=1 filter=255 channel=6
    5, -9, -2, 9, 6, -10, 1, 6, -2,
    -- layer=1 filter=255 channel=7
    -8, -1, -10, -2, -5, -5, -6, 7, -10,
    -- layer=1 filter=255 channel=8
    0, 9, -1, 0, 7, 3, 7, -5, 10,
    -- layer=1 filter=255 channel=9
    7, -4, -5, 0, 4, -4, -1, 5, -7,
    -- layer=1 filter=255 channel=10
    6, -6, 7, -3, -2, -4, 6, -5, -6,
    -- layer=1 filter=255 channel=11
    0, 5, -2, -11, 6, 0, 6, -8, -1,
    -- layer=1 filter=255 channel=12
    8, -10, 0, 4, 0, -9, -10, 7, 0,
    -- layer=1 filter=255 channel=13
    -1, 6, 7, -4, 7, 7, -11, -4, -8,
    -- layer=1 filter=255 channel=14
    -8, 6, -9, 0, 6, 5, -6, 9, 6,
    -- layer=1 filter=255 channel=15
    -3, -4, -10, 0, -10, -10, -8, -3, 9,
    -- layer=1 filter=255 channel=16
    -7, 9, -12, -6, 0, 7, -4, -7, -9,
    -- layer=1 filter=255 channel=17
    7, -10, -10, -10, 0, 4, -11, 6, -5,
    -- layer=1 filter=255 channel=18
    5, 3, 7, -10, 3, 0, 2, -6, -9,
    -- layer=1 filter=255 channel=19
    6, 1, -10, -8, 3, -4, 7, -7, -8,
    -- layer=1 filter=255 channel=20
    -4, 1, 0, 1, -6, 5, 4, 0, -8,
    -- layer=1 filter=255 channel=21
    -9, 9, -7, -10, -1, 7, -9, -6, 6,
    -- layer=1 filter=255 channel=22
    2, -8, -8, -2, -7, -10, -8, -7, -5,
    -- layer=1 filter=255 channel=23
    9, 0, -6, -3, -3, -7, -7, 0, -8,
    -- layer=1 filter=255 channel=24
    2, -5, -8, -7, 5, -7, -8, 1, -4,
    -- layer=1 filter=255 channel=25
    -2, -3, 5, 3, 2, 4, 2, 7, 2,
    -- layer=1 filter=255 channel=26
    -3, -3, -6, -9, -10, -11, -6, 4, -9,
    -- layer=1 filter=255 channel=27
    0, 6, 4, 2, -8, 2, -5, 9, 1,
    -- layer=1 filter=255 channel=28
    2, -2, 0, -3, 1, -2, -6, 0, -6,
    -- layer=1 filter=255 channel=29
    -10, 9, 3, 6, -6, 7, -6, 3, -9,
    -- layer=1 filter=255 channel=30
    7, -1, 0, 5, 0, -1, 8, -5, 3,
    -- layer=1 filter=255 channel=31
    -9, -5, 3, -6, 0, -4, -8, 5, -1,
    -- layer=1 filter=255 channel=32
    -8, -2, -8, 0, 0, -5, -5, 0, -6,
    -- layer=1 filter=255 channel=33
    1, 2, 9, 9, 8, 5, 9, -4, -4,
    -- layer=1 filter=255 channel=34
    -1, -7, 2, 2, -4, 7, -4, 9, 7,
    -- layer=1 filter=255 channel=35
    -2, 2, -5, -6, -8, -4, 0, -7, 2,
    -- layer=1 filter=255 channel=36
    -5, -2, -10, 8, -6, 3, -6, 4, -6,
    -- layer=1 filter=255 channel=37
    -6, 3, 7, 6, 6, 3, 6, -5, -3,
    -- layer=1 filter=255 channel=38
    2, 7, -3, 5, 0, -9, 2, 7, 0,
    -- layer=1 filter=255 channel=39
    -5, 4, 0, -3, 3, 2, 8, 0, -5,
    -- layer=1 filter=255 channel=40
    -10, 5, 1, -6, 3, 4, 6, -6, 8,
    -- layer=1 filter=255 channel=41
    -8, 8, -10, -5, 9, 6, 1, -4, 7,
    -- layer=1 filter=255 channel=42
    0, -7, 3, 0, -5, -10, 3, -9, 7,
    -- layer=1 filter=255 channel=43
    -5, -10, 7, 9, 0, -1, -10, -2, -5,
    -- layer=1 filter=255 channel=44
    0, -2, -4, 8, -3, -6, 5, 6, 9,
    -- layer=1 filter=255 channel=45
    6, 4, 5, 0, -3, -11, -4, -4, 3,
    -- layer=1 filter=255 channel=46
    3, 5, 0, 4, 5, 4, 2, 5, -9,
    -- layer=1 filter=255 channel=47
    3, 8, 0, -2, 3, 2, -2, 0, -5,
    -- layer=1 filter=255 channel=48
    5, 0, -9, 0, -3, 2, -5, 1, -6,
    -- layer=1 filter=255 channel=49
    -10, 8, 3, -1, 6, 2, 3, -11, 1,
    -- layer=1 filter=255 channel=50
    -5, 8, 2, 4, 9, -4, 0, -6, 8,
    -- layer=1 filter=255 channel=51
    -4, 3, -3, 8, 5, -8, -10, -8, -8,
    -- layer=1 filter=255 channel=52
    9, 6, -5, 0, 4, 7, -6, -3, 8,
    -- layer=1 filter=255 channel=53
    -10, 0, 1, 10, -9, -4, 6, -7, 5,
    -- layer=1 filter=255 channel=54
    -7, -3, 0, 8, -4, -8, -6, -2, -10,
    -- layer=1 filter=255 channel=55
    -9, -8, 4, -7, -1, -5, -5, 4, -1,
    -- layer=1 filter=255 channel=56
    0, -7, -5, -1, 0, 2, 4, -3, 3,
    -- layer=1 filter=255 channel=57
    0, -9, 5, -2, -4, 3, 0, -3, -3,
    -- layer=1 filter=255 channel=58
    0, -1, 0, 0, 0, -2, -2, 1, -8,
    -- layer=1 filter=255 channel=59
    3, -3, -10, 3, 4, -7, 3, -3, -9,
    -- layer=1 filter=255 channel=60
    -6, 9, -7, -7, 9, 5, -8, 8, 7,
    -- layer=1 filter=255 channel=61
    -6, 8, -5, 4, 2, 1, -10, 6, -10,
    -- layer=1 filter=255 channel=62
    -4, 0, 6, 7, 2, 4, 5, 0, -9,
    -- layer=1 filter=255 channel=63
    8, -7, 8, 7, -7, -4, -10, 2, -10,
    -- layer=1 filter=255 channel=64
    -7, -5, -2, -9, 2, -3, -11, 3, -1,
    -- layer=1 filter=255 channel=65
    -7, -2, 4, -8, 3, -1, -9, 2, 4,
    -- layer=1 filter=255 channel=66
    5, -2, 6, -4, 0, -9, -5, 8, -11,
    -- layer=1 filter=255 channel=67
    5, -7, -8, 9, 2, 4, -4, 2, 9,
    -- layer=1 filter=255 channel=68
    -9, -3, -3, 1, 6, -1, 5, -7, 4,
    -- layer=1 filter=255 channel=69
    3, -9, -9, 4, -4, 0, -1, -7, -2,
    -- layer=1 filter=255 channel=70
    -5, 9, 3, -10, 5, 5, -10, -10, 5,
    -- layer=1 filter=255 channel=71
    2, -9, -5, -5, -5, 0, 2, 0, -7,
    -- layer=1 filter=255 channel=72
    6, 0, 8, -2, -3, 5, -6, 0, -10,
    -- layer=1 filter=255 channel=73
    5, 8, 0, -8, 8, -7, 2, 5, 1,
    -- layer=1 filter=255 channel=74
    -1, 2, 7, -3, -5, -3, -7, -5, 5,
    -- layer=1 filter=255 channel=75
    5, 3, 7, 3, -9, -3, -2, -2, -6,
    -- layer=1 filter=255 channel=76
    7, 2, -7, -9, -8, 8, 0, 9, -1,
    -- layer=1 filter=255 channel=77
    -11, 0, -10, 2, 9, 0, 6, -8, 0,
    -- layer=1 filter=255 channel=78
    -2, -9, -5, 6, -6, -9, -6, -4, -9,
    -- layer=1 filter=255 channel=79
    -7, 0, 0, -9, 10, 4, 0, 0, -5,
    -- layer=1 filter=255 channel=80
    -11, -6, -1, -4, 9, 9, 4, 8, -2,
    -- layer=1 filter=255 channel=81
    -7, -1, -6, 2, -4, 7, 6, -11, -5,
    -- layer=1 filter=255 channel=82
    3, 2, 8, -3, -6, 4, 0, 4, -8,
    -- layer=1 filter=255 channel=83
    8, -2, 2, -3, 7, -2, 1, -2, -7,
    -- layer=1 filter=255 channel=84
    -7, 8, 0, -7, 8, -3, 0, -4, 5,
    -- layer=1 filter=255 channel=85
    -3, 9, 9, 0, -3, 0, 2, 10, 6,
    -- layer=1 filter=255 channel=86
    -5, -1, 3, 0, 0, -8, -2, 5, 8,
    -- layer=1 filter=255 channel=87
    -6, -1, 0, 2, -8, 8, 4, -7, -8,
    -- layer=1 filter=255 channel=88
    3, -8, 9, -1, -5, 0, 4, 4, -2,
    -- layer=1 filter=255 channel=89
    1, -11, -10, -4, -5, 8, 0, -11, -3,
    -- layer=1 filter=255 channel=90
    -5, 3, 4, 8, -9, -2, 3, 8, -9,
    -- layer=1 filter=255 channel=91
    -5, -5, 5, -6, 4, -12, -5, 4, -3,
    -- layer=1 filter=255 channel=92
    7, -8, -1, 7, 0, 7, -9, -3, 8,
    -- layer=1 filter=255 channel=93
    -1, 2, -7, 7, -10, -6, -3, -1, -5,
    -- layer=1 filter=255 channel=94
    -5, 1, 2, -9, -2, -3, -8, 6, -1,
    -- layer=1 filter=255 channel=95
    3, -5, 0, 7, 0, 6, 0, -9, -6,
    -- layer=1 filter=255 channel=96
    1, 0, -8, -9, -7, 10, 8, -8, -6,
    -- layer=1 filter=255 channel=97
    -5, 3, -10, 4, -6, -4, -4, -5, -8,
    -- layer=1 filter=255 channel=98
    3, 7, -4, -8, 0, 4, -3, 4, -7,
    -- layer=1 filter=255 channel=99
    -8, -8, -1, -10, -2, -7, -7, 4, 8,
    -- layer=1 filter=255 channel=100
    -8, 2, -3, 3, -1, 0, -3, -8, 6,
    -- layer=1 filter=255 channel=101
    -10, -1, -7, 0, 3, 3, -2, 5, -7,
    -- layer=1 filter=255 channel=102
    3, 6, -10, 0, -3, -9, -10, -3, 10,
    -- layer=1 filter=255 channel=103
    2, -9, 0, -6, -10, -1, -6, -8, 1,
    -- layer=1 filter=255 channel=104
    3, -2, 4, 2, 0, -8, -8, 3, -6,
    -- layer=1 filter=255 channel=105
    -1, 6, 0, -7, -2, 3, -3, -6, -3,
    -- layer=1 filter=255 channel=106
    -10, -2, -10, 1, -5, -12, 0, 1, -10,
    -- layer=1 filter=255 channel=107
    1, 8, -3, 0, 8, -6, -7, 6, -5,
    -- layer=1 filter=255 channel=108
    4, -9, 5, 5, 1, -7, 2, -8, -1,
    -- layer=1 filter=255 channel=109
    0, 6, -5, 6, -4, -1, -6, -5, 9,
    -- layer=1 filter=255 channel=110
    7, -4, -6, 1, -10, -8, -8, -8, -6,
    -- layer=1 filter=255 channel=111
    -11, -4, 7, 2, 6, -6, 10, 0, -10,
    -- layer=1 filter=255 channel=112
    -10, 0, 3, -3, 4, 5, 3, 3, -1,
    -- layer=1 filter=255 channel=113
    0, 0, 0, 1, -2, 7, 2, 9, 5,
    -- layer=1 filter=255 channel=114
    6, -4, -7, 5, -6, 7, -6, -7, 4,
    -- layer=1 filter=255 channel=115
    -5, -10, -7, 6, -8, 8, -8, -7, 0,
    -- layer=1 filter=255 channel=116
    7, 0, 5, -3, -8, 8, 6, -4, -7,
    -- layer=1 filter=255 channel=117
    3, 6, -9, -9, 4, 4, 8, 8, 5,
    -- layer=1 filter=255 channel=118
    -3, 1, -10, -4, -7, 7, -7, 0, -1,
    -- layer=1 filter=255 channel=119
    -4, 1, -2, -9, -5, -3, -9, 6, 8,
    -- layer=1 filter=255 channel=120
    -8, 7, 6, -9, -9, 0, -6, -7, 6,
    -- layer=1 filter=255 channel=121
    -5, -10, 8, -7, -3, 7, -5, 8, 1,
    -- layer=1 filter=255 channel=122
    5, 0, -8, -4, -8, -4, 5, 8, -9,
    -- layer=1 filter=255 channel=123
    8, -10, 0, -4, 0, -11, -6, -1, -9,
    -- layer=1 filter=255 channel=124
    1, -6, -8, 9, -7, 0, -8, 4, 7,
    -- layer=1 filter=255 channel=125
    -3, 0, -9, -6, 5, -4, 5, 1, 3,
    -- layer=1 filter=255 channel=126
    4, 2, 2, -2, 1, -5, -2, 8, 0,
    -- layer=1 filter=255 channel=127
    8, 0, -2, -6, -8, -7, -7, -7, -3,

    others => 0);
end iwght_package;
