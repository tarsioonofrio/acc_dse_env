library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    588, 408, 450, 449, 458, 153, 35, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 114, 147, 83, 0, 0, 40, 222, 208, 308, 196, 123, 136, 113, 230, 129, 0, 14, 24, 0, 0, 85, 0, 53, 230, 0, 0, 202, 0, 0, 0, 234, 0, 0, 0, 0, 0, 59, 0, 0, 0, 156, 189, 471, 173, 52, 272, 234, 253, 0, 270, 242, 0, 210, 203, 360, 301, 0, 0, 184, 76, 141, 192, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 91, 0, 0, 0, 0, 0, 0, 0, 0, 297, 235, 231, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 110, 0, 0, 26, 0, 0, 0, 112, 152, 0, 0, 0, 14, 209, 259, 182, 7, 28, 0, 0, 0, 18, 0, 47, 0, 97, 215, 13, 0, 190, 239, 210, 332, 374, 0, 0, 0, 0, 0, 0, 0, 0, 0, 417, 62, 266, 82, 528, 429, 110, 287, 339, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 198, 0, 158, 0, 21, 138, 191, 119, 44, 0, 297, 142, 136, 253, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 351, 297, 308, 129, 416, 358, 0, 19, 0, 0, 87, 99, 110, 0, 0, 0, 0, 0, 310, 83, 80, 0, 0, 158, 0, 41, 132, 0, 91, 0, 0, 0, 0, 599, 811, 1065, 476, 417, 214, 60, 27, 0, 0, 0, 0, 47, 274, 173, 241, 191, 15, 167, 98, 174, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 100, 0, 0, 0, 0, 0, 0, 240, 360, 444, 0, 353, 264, 0, 0, 194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 90, 21, 299, 156, 0, 0, 0, 164, 0, 28, 168, 0, 49, 0, 103, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 97, 0, 243, 287, 310, 701, 71, 156, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 224, 140, 0, 0, 235, 0, 328, 56, 577, 463, 280, 249, 245, 0, 0, 0, 199, 35, 0, 0, 0, 0, 0, 0, 0, 153, 214, 85, 173, 106, 22, 0, 69, 0, 89, 82, 86, 562, 209, 68, 428, 338, 192, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 47, 0, 0, 0, 0, 58, 0, 0, 0, 0, 399, 49, 261, 73, 13, 0, 0, 0, 539, 632, 592, 290, 578, 329, 144, 100, 141, 28, 175, 58, 0, 0, 0, 53, 0, 0, 192, 0, 0, 0, 171, 40, 236, 0, 0, 0, 0, 0, 0, 0, 0, 70, 166, 0, 585, 486, 455, 407, 330, 364, 0, 0, 0, 0, 0, 0, 24, 0, 0, 295, 177, 80, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 113, 9, 40, 2, 0, 0, 0, 525, 303, 140, 361, 106, 0, 171, 0, 182, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 193, 0, 0, 146, 0, 0, 0, 398, 423, 487, 454, 237, 226, 195, 0, 0, 285, 179, 204, 474, 322, 225, 95, 173, 166, 0, 0, 0, 0, 0, 0, 0, 0, 0,
    others => 0);
end ifmap_package;
