library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    115, 174, 163, 174, 107, 112, 111, 82, 
    50, 151, 140, 169, 70, 65, 99, 165, 
    0, 0, 0, 32, 0, 0, 8, 109, 
    0, 0, 0, 0, 0, 0, 1, 104, 
    0, 0, 0, 0, 0, 0, 0, 53, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 2, 0, 9, 78, 
    0, 0, 0, 0, 6, 0, 67, 89, 
    0, 0, 0, 0, 0, 0, 57, 61, 
    0, 5, 0, 0, 25, 42, 50, 12, 
    0, 0, 0, 88, 50, 49, 0, 23, 
    0, 0, 17, 161, 63, 28, 2, 41, 
    0, 0, 57, 84, 0, 0, 0, 68, 
    
    -- channel=3
    467, 401, 345, 234, 182, 192, 154, 0, 
    812, 514, 370, 120, 131, 84, 0, 0, 
    849, 343, 191, 0, 41, 0, 0, 0, 
    921, 55, 23, 0, 0, 0, 0, 0, 
    928, 0, 0, 0, 0, 0, 0, 0, 
    1072, 0, 0, 0, 0, 0, 0, 0, 
    1094, 0, 0, 0, 0, 0, 0, 0, 
    866, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    301, 108, 124, 78, 24, 26, 21, 0, 
    316, 25, 45, 15, 0, 0, 0, 0, 
    265, 0, 0, 0, 0, 0, 9, 0, 
    192, 0, 48, 117, 20, 47, 99, 0, 
    166, 0, 31, 0, 40, 14, 97, 0, 
    134, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 23, 8, 0, 0, 0, 158, 
    
    -- channel=5
    0, 27, 35, 15, 3, 0, 37, 77, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 150, 74, 0, 0, 
    61, 277, 252, 205, 344, 151, 4, 0, 
    211, 333, 292, 127, 386, 145, 57, 0, 
    462, 418, 196, 0, 0, 0, 0, 0, 
    570, 866, 679, 490, 221, 390, 401, 262, 
    492, 690, 650, 784, 702, 959, 1204, 637, 
    443, 345, 274, 558, 829, 1184, 1304, 599, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 19, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 92, 0, 95, 79, 0, 0, 
    0, 0, 0, 4, 12, 0, 0, 0, 
    0, 0, 0, 76, 0, 0, 0, 1, 
    135, 278, 212, 48, 0, 0, 0, 0, 
    499, 612, 445, 329, 385, 463, 482, 262, 
    
    -- channel=8
    104, 211, 179, 145, 96, 91, 170, 125, 
    118, 349, 369, 309, 248, 208, 370, 336, 
    0, 67, 126, 92, 42, 85, 281, 269, 
    0, 0, 0, 38, 1, 101, 240, 206, 
    0, 0, 0, 0, 0, 0, 70, 106, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=9
    347, 509, 539, 518, 625, 541, 346, 109, 
    607, 770, 711, 616, 621, 352, 114, 20, 
    570, 559, 516, 414, 433, 156, 136, 89, 
    341, 224, 87, 0, 0, 0, 0, 33, 
    366, 564, 388, 149, 0, 191, 568, 341, 
    117, 343, 162, 70, 269, 675, 859, 332, 
    0, 0, 0, 0, 190, 406, 349, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    560, 554, 562, 457, 352, 344, 317, 0, 
    912, 761, 812, 628, 445, 394, 374, 0, 
    779, 568, 667, 558, 341, 239, 277, 0, 
    573, 250, 447, 448, 298, 206, 285, 0, 
    506, 139, 336, 234, 152, 85, 198, 0, 
    363, 0, 0, 0, 0, 0, 0, 0, 
    93, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    0, 225, 176, 347, 204, 259, 466, 396, 
    0, 203, 60, 321, 135, 199, 540, 363, 
    0, 251, 0, 247, 144, 217, 599, 441, 
    0, 287, 0, 89, 186, 214, 404, 451, 
    0, 121, 142, 191, 145, 20, 79, 481, 
    0, 0, 293, 319, 0, 0, 0, 600, 
    0, 0, 4, 134, 0, 0, 0, 738, 
    0, 0, 0, 0, 0, 0, 0, 292, 
    
    -- channel=12
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=13
    6, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 49, 37, 0, 0, 0, 0, 
    0, 0, 0, 90, 206, 27, 59, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 160, 118, 80, 0, 0, 0, 0, 
    209, 535, 564, 413, 85, 3, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    105, 167, 38, 13, 0, 0, 0, 0, 
    269, 465, 206, 359, 261, 361, 391, 164, 
    419, 804, 573, 742, 809, 979, 1147, 728, 
    486, 719, 609, 735, 848, 997, 1119, 672, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 32, 
    0, 0, 0, 0, 0, 0, 55, 122, 
    0, 0, 0, 0, 0, 10, 24, 133, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 0, 
    160, 196, 23, 7, 0, 0, 57, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 153, 101, 0, 0, 0, 0, 0, 
    0, 0, 102, 179, 128, 126, 91, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    107, 0, 0, 0, 0, 0, 0, 0, 
    208, 122, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 56, 59, 121, 121, 72, 6, 
    93, 126, 157, 95, 199, 150, 78, 0, 
    311, 356, 326, 252, 360, 268, 178, 14, 
    492, 529, 370, 214, 270, 155, 85, 39, 
    585, 854, 677, 449, 322, 268, 295, 211, 
    572, 953, 856, 726, 561, 683, 807, 500, 
    565, 828, 670, 719, 810, 1036, 1228, 721, 
    292, 317, 122, 251, 404, 508, 600, 293, 
    
    -- channel=19
    101, 0, 0, 0, 0, 0, 0, 0, 
    503, 92, 0, 0, 0, 0, 0, 0, 
    585, 54, 0, 0, 0, 0, 0, 0, 
    756, 0, 0, 0, 0, 0, 0, 0, 
    811, 0, 0, 0, 0, 0, 0, 0, 
    1078, 0, 0, 0, 0, 0, 0, 0, 
    1340, 193, 0, 0, 0, 0, 4, 0, 
    1137, 321, 0, 0, 0, 19, 0, 0, 
    
    -- channel=20
    346, 389, 293, 257, 154, 117, 244, 152, 
    437, 522, 381, 272, 224, 137, 279, 131, 
    244, 323, 195, 60, 68, 0, 93, 18, 
    69, 0, 99, 0, 1, 37, 40, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    147, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=21
    241, 107, 160, 27, 115, 98, 0, 0, 
    201, 0, 0, 0, 0, 0, 0, 0, 
    456, 0, 80, 0, 27, 0, 0, 0, 
    616, 0, 13, 0, 0, 0, 0, 0, 
    788, 103, 0, 0, 0, 0, 55, 0, 
    898, 437, 0, 0, 34, 157, 278, 0, 
    790, 436, 42, 99, 380, 535, 574, 0, 
    338, 136, 93, 302, 415, 496, 511, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    297, 0, 20, 0, 145, 16, 0, 0, 
    722, 153, 166, 39, 45, 0, 0, 0, 
    984, 432, 260, 170, 207, 143, 87, 0, 
    1188, 717, 474, 390, 484, 652, 713, 48, 
    1334, 933, 655, 623, 905, 1163, 1215, 157, 
    1045, 559, 349, 479, 697, 831, 868, 17, 
    
    -- channel=23
    0, 0, 0, 0, 0, 31, 0, 0, 
    267, 71, 130, 169, 29, 336, 166, 100, 
    469, 154, 152, 236, 35, 375, 155, 109, 
    628, 275, 130, 297, 63, 311, 130, 136, 
    618, 399, 266, 278, 261, 294, 268, 345, 
    545, 463, 463, 274, 413, 371, 508, 663, 
    541, 605, 654, 343, 424, 411, 579, 774, 
    372, 503, 467, 215, 258, 247, 389, 580, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 53, 
    0, 34, 107, 118, 62, 51, 86, 136, 
    0, 0, 0, 0, 0, 12, 40, 86, 
    0, 0, 20, 22, 6, 3, 0, 49, 
    0, 0, 45, 104, 180, 136, 81, 84, 
    0, 0, 0, 35, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 23, 0, 0, 0, 0, 0, 0, 
    
    -- channel=25
    53, 113, 151, 149, 109, 131, 128, 116, 
    19, 140, 126, 116, 71, 63, 59, 32, 
    0, 74, 37, 49, 80, 57, 0, 45, 
    0, 33, 62, 0, 29, 0, 0, 22, 
    0, 0, 111, 48, 7, 0, 0, 88, 
    0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=26
    145, 273, 296, 330, 267, 252, 238, 161, 
    13, 211, 181, 242, 120, 107, 33, 88, 
    0, 160, 111, 150, 88, 85, 18, 97, 
    0, 68, 68, 3, 0, 0, 0, 109, 
    0, 4, 159, 74, 0, 47, 24, 275, 
    0, 0, 0, 0, 0, 0, 0, 213, 
    0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    110, 124, 80, 44, 0, 1, 86, 126, 
    100, 350, 327, 277, 187, 175, 281, 343, 
    0, 31, 68, 22, 0, 59, 166, 269, 
    0, 0, 74, 19, 0, 61, 108, 200, 
    0, 0, 0, 0, 0, 0, 0, 155, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=28
    351, 276, 245, 166, 149, 131, 122, 53, 
    304, 235, 164, 137, 61, 75, 56, 54, 
    189, 20, 25, 59, 0, 8, 36, 56, 
    89, 0, 0, 10, 0, 0, 82, 67, 
    40, 0, 0, 0, 0, 0, 36, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    95, 4, 0, 0, 0, 0, 0, 0, 
    304, 173, 106, 0, 41, 0, 0, 0, 
    477, 161, 154, 0, 0, 0, 0, 0, 
    598, 103, 136, 0, 0, 0, 0, 0, 
    714, 82, 0, 53, 0, 0, 0, 0, 
    882, 172, 0, 0, 0, 42, 197, 0, 
    958, 303, 0, 0, 0, 129, 156, 0, 
    623, 44, 0, 0, 0, 0, 0, 0, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    125, 0, 0, 0, 0, 0, 0, 0, 
    340, 109, 0, 0, 0, 0, 0, 0, 
    581, 469, 289, 125, 102, 229, 334, 50, 
    829, 792, 548, 636, 854, 1137, 1327, 722, 
    771, 729, 502, 710, 972, 1194, 1274, 620, 
    
    -- channel=31
    25, 87, 41, 51, 62, 25, 71, 8, 
    0, 0, 0, 0, 21, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=32
    750, 901, 878, 739, 598, 563, 564, 254, 
    785, 904, 874, 706, 531, 461, 474, 242, 
    483, 467, 512, 467, 269, 236, 348, 195, 
    34, 0, 133, 195, 154, 139, 386, 194, 
    0, 0, 0, 0, 0, 0, 101, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=33
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 100, 89, 
    0, 0, 0, 0, 0, 0, 38, 0, 
    0, 0, 0, 16, 0, 0, 66, 0, 
    0, 0, 0, 22, 54, 149, 112, 0, 
    0, 0, 0, 21, 102, 39, 0, 0, 
    0, 5, 82, 12, 0, 0, 0, 0, 
    5, 315, 350, 101, 0, 0, 0, 36, 
    
    -- channel=34
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=35
    439, 534, 434, 371, 365, 233, 388, 179, 
    462, 607, 460, 324, 381, 203, 376, 168, 
    290, 430, 384, 161, 255, 103, 298, 88, 
    109, 107, 253, 137, 159, 191, 280, 57, 
    35, 0, 0, 92, 0, 58, 102, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=36
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 41, 0, 0, 0, 
    109, 239, 81, 0, 74, 0, 0, 0, 
    278, 425, 279, 218, 159, 192, 132, 0, 
    473, 611, 460, 530, 493, 618, 573, 185, 
    646, 750, 672, 845, 878, 1018, 1057, 524, 
    542, 569, 580, 638, 659, 784, 822, 386, 
    
    -- channel=38
    17, 19, 0, 0, 26, 0, 0, 0, 
    113, 166, 92, 59, 124, 0, 11, 0, 
    33, 107, 45, 0, 84, 0, 0, 0, 
    15, 139, 85, 9, 35, 0, 1, 0, 
    27, 62, 50, 48, 89, 122, 139, 0, 
    129, 0, 0, 28, 116, 137, 66, 0, 
    203, 73, 0, 106, 55, 71, 0, 0, 
    67, 32, 0, 27, 0, 0, 0, 0, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 26, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    6, 0, 0, 0, 0, 0, 0, 0, 
    208, 294, 292, 167, 0, 0, 0, 0, 
    789, 1257, 1314, 1116, 968, 1106, 1189, 855, 
    
    -- channel=40
    0, 0, 0, 0, 0, 0, 0, 0, 
    107, 0, 0, 0, 10, 105, 0, 0, 
    444, 0, 29, 36, 72, 150, 0, 0, 
    934, 195, 211, 185, 71, 34, 0, 0, 
    1083, 543, 429, 370, 403, 439, 403, 65, 
    1217, 740, 559, 511, 791, 870, 904, 322, 
    1403, 1000, 903, 875, 1058, 1146, 1220, 455, 
    934, 721, 697, 587, 584, 622, 685, 256, 
    
    -- channel=41
    261, 277, 270, 230, 267, 235, 203, 0, 
    455, 628, 538, 435, 378, 263, 199, 0, 
    394, 430, 343, 229, 198, 92, 132, 0, 
    209, 174, 84, 0, 0, 0, 0, 0, 
    127, 275, 198, 174, 0, 113, 315, 102, 
    0, 0, 0, 0, 6, 230, 395, 93, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    0, 0, 0, 92, 0, 63, 372, 434, 
    0, 0, 0, 287, 0, 296, 781, 729, 
    0, 0, 0, 316, 0, 479, 999, 869, 
    0, 312, 0, 339, 153, 615, 740, 910, 
    0, 228, 218, 432, 334, 319, 227, 1179, 
    0, 0, 723, 704, 241, 0, 0, 1632, 
    0, 0, 941, 694, 0, 0, 0, 2184, 
    0, 83, 641, 335, 0, 0, 0, 1635, 
    
    -- channel=43
    154, 396, 458, 382, 257, 245, 316, 125, 
    83, 525, 597, 532, 393, 290, 461, 207, 
    0, 294, 402, 417, 297, 127, 405, 178, 
    0, 78, 394, 351, 411, 186, 429, 145, 
    0, 0, 253, 263, 244, 45, 124, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=44
    75, 20, 6, 9, 0, 14, 12, 0, 
    144, 0, 0, 0, 0, 0, 54, 0, 
    90, 0, 0, 16, 0, 33, 92, 0, 
    80, 44, 0, 47, 0, 59, 78, 0, 
    44, 84, 4, 0, 0, 0, 0, 0, 
    0, 0, 62, 0, 0, 0, 0, 37, 
    0, 0, 59, 0, 0, 0, 0, 194, 
    0, 98, 47, 0, 0, 0, 22, 340, 
    
    -- channel=45
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    202, 534, 350, 464, 196, 94, 98, 0, 
    777, 1473, 1368, 1297, 1166, 1304, 1434, 1007, 
    
    -- channel=46
    43, 0, 0, 0, 0, 0, 0, 0, 
    33, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 80, 80, 9, 32, 0, 0, 0, 
    0, 118, 129, 65, 134, 67, 63, 0, 
    37, 72, 0, 0, 0, 0, 0, 0, 
    21, 141, 102, 245, 66, 77, 0, 0, 
    26, 232, 150, 204, 86, 98, 66, 54, 
    
    -- channel=47
    0, 0, 0, 0, 0, 0, 0, 0, 
    38, 0, 0, 0, 0, 0, 0, 0, 
    169, 0, 0, 0, 0, 0, 0, 0, 
    346, 0, 0, 0, 0, 0, 0, 0, 
    536, 0, 0, 0, 0, 0, 0, 0, 
    788, 0, 0, 0, 0, 0, 0, 0, 
    920, 74, 0, 0, 0, 0, 0, 0, 
    994, 361, 0, 0, 114, 204, 226, 0, 
    
    -- channel=48
    546, 734, 722, 607, 500, 450, 551, 276, 
    593, 761, 726, 579, 452, 352, 488, 220, 
    274, 387, 449, 338, 235, 154, 326, 149, 
    0, 0, 185, 165, 151, 133, 254, 122, 
    0, 0, 0, 12, 0, 0, 61, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=49
    39, 76, 34, 0, 0, 0, 0, 0, 
    188, 278, 280, 264, 137, 164, 143, 113, 
    0, 0, 40, 24, 0, 0, 52, 66, 
    0, 0, 0, 0, 0, 0, 35, 0, 
    0, 0, 0, 0, 0, 0, 16, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=50
    62, 187, 196, 266, 277, 301, 280, 105, 
    251, 570, 470, 455, 403, 325, 229, 62, 
    274, 614, 412, 324, 365, 179, 82, 78, 
    125, 315, 81, 0, 0, 0, 0, 0, 
    29, 374, 482, 228, 0, 0, 0, 329, 
    0, 36, 274, 262, 52, 349, 657, 687, 
    0, 0, 0, 0, 0, 242, 350, 241, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=51
    0, 0, 0, 0, 0, 0, 0, 0, 
    133, 272, 172, 191, 230, 66, 0, 0, 
    129, 228, 97, 96, 176, 24, 77, 0, 
    187, 421, 236, 143, 61, 0, 0, 0, 
    229, 660, 563, 450, 409, 377, 599, 292, 
    214, 579, 475, 446, 584, 760, 807, 384, 
    183, 389, 338, 591, 663, 785, 713, 428, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=52
    42, 38, 54, 30, 0, 0, 0, 203, 
    74, 27, 119, 57, 0, 51, 97, 353, 
    0, 0, 62, 0, 0, 0, 0, 196, 
    0, 0, 0, 0, 0, 64, 0, 172, 
    0, 0, 0, 0, 0, 0, 0, 27, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=53
    55, 9, 0, 0, 36, 0, 0, 0, 
    93, 0, 0, 0, 0, 0, 0, 0, 
    61, 0, 0, 0, 0, 0, 0, 0, 
    93, 0, 0, 0, 0, 0, 0, 0, 
    143, 0, 0, 0, 0, 0, 52, 0, 
    118, 0, 0, 0, 0, 4, 19, 0, 
    0, 0, 0, 11, 8, 16, 25, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=55
    570, 634, 625, 473, 418, 331, 347, 198, 
    706, 696, 688, 455, 356, 272, 349, 213, 
    424, 290, 425, 287, 136, 60, 232, 128, 
    41, 0, 50, 131, 46, 57, 306, 99, 
    0, 0, 0, 0, 0, 0, 75, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=56
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 50, 116, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 342, 248, 202, 0, 0, 0, 0, 
    743, 1452, 1332, 1219, 997, 1077, 1205, 1029, 
    
    -- channel=57
    5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=58
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 0, 141, 111, 78, 
    134, 80, 40, 100, 24, 182, 131, 84, 
    160, 96, 86, 131, 136, 189, 108, 84, 
    149, 34, 3, 49, 40, 0, 0, 51, 
    174, 157, 201, 92, 53, 33, 112, 221, 
    279, 340, 226, 106, 134, 136, 233, 350, 
    513, 514, 416, 390, 401, 427, 517, 373, 
    
    -- channel=59
    0, 0, 0, 8, 0, 3, 174, 286, 
    0, 0, 0, 161, 0, 120, 394, 438, 
    0, 14, 0, 111, 0, 243, 497, 481, 
    0, 205, 45, 205, 122, 309, 352, 481, 
    0, 110, 221, 381, 251, 278, 164, 687, 
    0, 0, 345, 409, 123, 0, 0, 829, 
    0, 0, 506, 355, 0, 0, 0, 1064, 
    0, 52, 323, 74, 0, 0, 0, 717, 
    
    -- channel=60
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    130, 0, 0, 0, 0, 0, 0, 0, 
    291, 0, 0, 0, 0, 0, 0, 0, 
    453, 239, 0, 40, 40, 126, 167, 0, 
    548, 566, 397, 446, 558, 713, 883, 634, 
    539, 741, 589, 615, 781, 941, 1077, 861, 
    
    -- channel=61
    324, 185, 165, 4, 132, 16, 27, 0, 
    444, 344, 222, 0, 316, 0, 0, 0, 
    474, 313, 216, 0, 326, 0, 0, 0, 
    439, 93, 267, 0, 212, 0, 0, 0, 
    471, 0, 70, 0, 7, 0, 114, 0, 
    632, 119, 0, 0, 0, 96, 217, 0, 
    660, 201, 0, 0, 13, 179, 125, 0, 
    331, 30, 0, 45, 92, 149, 35, 0, 
    
    -- channel=62
    281, 331, 141, 33, 276, 0, 26, 0, 
    256, 418, 98, 0, 273, 0, 0, 0, 
    141, 374, 165, 0, 316, 0, 0, 0, 
    93, 226, 133, 0, 99, 0, 113, 0, 
    257, 310, 0, 0, 0, 119, 239, 0, 
    458, 252, 0, 0, 28, 272, 192, 0, 
    285, 26, 0, 189, 199, 348, 129, 0, 
    0, 0, 0, 83, 51, 116, 0, 0, 
    
    -- channel=63
    0, 0, 0, 0, 0, 18, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 
    80, 0, 0, 0, 0, 0, 0, 0, 
    95, 0, 0, 0, 0, 0, 0, 88, 
    99, 0, 0, 0, 0, 61, 97, 178, 
    84, 0, 0, 0, 50, 119, 102, 105, 
    0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end ifmap_package;
