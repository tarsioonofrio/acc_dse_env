library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 8, 11, 8, 7, 6, 3, 9, 0, 0, 0, 0, 8, 5, 
    10, 14, 12, 9, 11, 60, 33, 0, 0, 0, 26, 6, 0, 0, 6, 
    0, 0, 6, 6, 7, 0, 0, 0, 5, 18, 21, 9, 15, 0, 0, 
    37, 31, 10, 8, 14, 0, 48, 25, 3, 0, 0, 0, 0, 0, 0, 
    37, 79, 26, 19, 118, 100, 16, 12, 0, 0, 37, 37, 11, 16, 0, 
    6, 0, 19, 0, 0, 0, 30, 29, 29, 40, 14, 0, 0, 10, 32, 
    27, 0, 0, 4, 0, 22, 0, 17, 10, 11, 0, 12, 0, 14, 28, 
    35, 7, 39, 19, 20, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    26, 7, 21, 0, 40, 0, 0, 17, 2, 0, 0, 0, 0, 0, 33, 
    0, 1, 10, 1, 17, 5, 0, 61, 31, 0, 0, 0, 16, 29, 2, 
    0, 8, 0, 59, 130, 125, 37, 0, 0, 0, 24, 48, 13, 0, 0, 
    0, 0, 17, 66, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 2, 0, 0, 0, 0, 0, 1, 5, 16, 0, 0, 15, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 16, 3, 0, 31, 35, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 5, 0, 0, 10, 6, 0, 0, 0, 0, 11, 11, 0, 0, 0, 
    34, 7, 0, 0, 0, 0, 3, 0, 1, 0, 15, 0, 0, 0, 0, 
    29, 7, 0, 0, 0, 0, 28, 6, 2, 0, 9, 1, 0, 0, 0, 
    33, 20, 29, 0, 0, 6, 0, 0, 0, 0, 0, 14, 0, 0, 0, 
    27, 25, 26, 0, 12, 0, 0, 0, 2, 7, 13, 0, 0, 0, 0, 
    8, 13, 27, 0, 3, 3, 20, 41, 41, 0, 6, 15, 24, 8, 9, 
    66, 39, 25, 0, 71, 75, 50, 49, 57, 50, 56, 60, 64, 65, 69, 
    82, 57, 26, 22, 86, 56, 58, 54, 56, 58, 64, 65, 74, 78, 71, 
    92, 68, 54, 61, 64, 57, 56, 55, 60, 64, 76, 82, 79, 79, 100, 
    89, 80, 66, 58, 62, 66, 72, 62, 56, 59, 71, 70, 60, 81, 89, 
    
    -- channel=2
    82, 81, 83, 77, 78, 79, 87, 89, 78, 71, 69, 76, 71, 67, 62, 
    79, 85, 90, 80, 87, 50, 55, 72, 69, 38, 0, 14, 54, 74, 63, 
    51, 114, 87, 82, 92, 99, 28, 27, 25, 44, 0, 0, 0, 53, 71, 
    0, 75, 74, 89, 53, 64, 2, 0, 2, 86, 0, 21, 0, 0, 98, 
    0, 26, 41, 120, 0, 23, 0, 0, 0, 87, 0, 0, 1, 0, 58, 
    0, 16, 27, 84, 94, 45, 0, 0, 0, 124, 0, 0, 21, 0, 0, 
    0, 0, 57, 21, 98, 56, 9, 0, 0, 113, 0, 0, 9, 8, 0, 
    0, 0, 2, 10, 78, 78, 0, 23, 0, 90, 0, 0, 27, 27, 25, 
    0, 3, 0, 30, 15, 59, 1, 0, 33, 23, 38, 0, 36, 39, 60, 
    0, 7, 0, 45, 0, 35, 44, 0, 8, 29, 0, 6, 38, 73, 61, 
    43, 9, 0, 84, 0, 0, 44, 1, 0, 0, 0, 0, 0, 8, 0, 
    45, 33, 0, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 37, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 94, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    19, 21, 29, 27, 26, 20, 28, 28, 21, 6, 4, 11, 24, 21, 17, 
    28, 27, 28, 27, 29, 60, 24, 13, 0, 0, 6, 0, 0, 7, 21, 
    0, 18, 27, 27, 21, 0, 0, 0, 0, 11, 0, 10, 1, 0, 19, 
    0, 21, 21, 26, 17, 16, 12, 3, 1, 0, 12, 0, 0, 0, 0, 
    22, 31, 32, 28, 82, 57, 0, 0, 0, 7, 0, 4, 0, 5, 0, 
    0, 3, 37, 0, 0, 0, 25, 0, 0, 17, 6, 0, 0, 4, 11, 
    1, 0, 0, 15, 0, 20, 0, 27, 0, 3, 0, 0, 0, 0, 4, 
    6, 4, 6, 20, 4, 0, 11, 0, 0, 0, 0, 0, 0, 0, 15, 
    7, 0, 0, 5, 4, 0, 0, 0, 6, 0, 0, 0, 0, 6, 25, 
    0, 0, 0, 0, 0, 14, 17, 18, 0, 0, 0, 0, 10, 32, 17, 
    0, 0, 0, 18, 100, 20, 23, 0, 10, 2, 0, 7, 0, 0, 0, 
    0, 0, 17, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    90, 93, 99, 96, 95, 93, 102, 105, 96, 69, 57, 68, 81, 85, 81, 
    98, 105, 102, 98, 99, 116, 89, 79, 52, 50, 37, 34, 42, 64, 78, 
    44, 68, 101, 103, 103, 62, 55, 33, 32, 43, 16, 17, 15, 25, 70, 
    16, 67, 94, 101, 85, 71, 52, 20, 16, 26, 30, 22, 13, 9, 52, 
    15, 53, 78, 86, 81, 69, 38, 26, 7, 54, 44, 25, 23, 11, 25, 
    5, 33, 78, 86, 43, 52, 58, 30, 15, 67, 25, 10, 16, 12, 21, 
    20, 23, 54, 75, 49, 75, 28, 40, 7, 53, 20, 20, 23, 28, 22, 
    33, 26, 26, 59, 52, 36, 7, 19, 20, 53, 31, 14, 16, 21, 47, 
    26, 25, 10, 38, 50, 25, 36, 34, 29, 54, 21, 0, 19, 50, 80, 
    31, 26, 6, 39, 7, 25, 47, 43, 20, 6, 0, 1, 28, 77, 74, 
    32, 34, 7, 66, 52, 18, 13, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 4, 18, 70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 30, 23, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=5
    0, 0, 0, 2, 6, 0, 2, 3, 4, 0, 0, 0, 0, 8, 9, 
    2, 0, 0, 4, 0, 0, 38, 2, 5, 0, 21, 20, 0, 0, 5, 
    11, 0, 0, 3, 0, 0, 36, 12, 0, 0, 18, 14, 42, 0, 0, 
    83, 0, 7, 0, 22, 0, 12, 27, 12, 0, 50, 1, 26, 25, 0, 
    71, 0, 53, 0, 0, 46, 48, 45, 22, 0, 13, 60, 0, 37, 0, 
    66, 0, 63, 26, 0, 4, 42, 34, 65, 0, 66, 58, 0, 22, 33, 
    67, 31, 0, 44, 0, 0, 0, 48, 49, 0, 67, 46, 2, 0, 30, 
    56, 21, 51, 26, 0, 0, 80, 2, 22, 0, 33, 48, 0, 0, 16, 
    52, 0, 111, 0, 48, 0, 14, 11, 0, 52, 0, 48, 0, 0, 0, 
    0, 0, 93, 0, 25, 24, 0, 18, 35, 0, 42, 0, 0, 0, 10, 
    0, 1, 84, 0, 112, 38, 0, 0, 53, 48, 0, 0, 0, 0, 11, 
    0, 0, 17, 0, 88, 38, 0, 0, 1, 0, 0, 0, 0, 0, 4, 
    28, 0, 0, 9, 93, 1, 4, 2, 2, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 39, 22, 0, 18, 1, 0, 0, 0, 0, 5, 0, 14, 
    38, 0, 4, 0, 11, 0, 0, 0, 0, 5, 14, 0, 0, 24, 46, 
    
    -- channel=6
    56, 66, 58, 60, 57, 63, 58, 56, 58, 64, 63, 59, 56, 47, 44, 
    53, 57, 59, 62, 61, 106, 58, 68, 68, 69, 67, 47, 47, 52, 48, 
    72, 65, 57, 59, 58, 113, 85, 46, 36, 98, 106, 88, 65, 30, 58, 
    66, 36, 55, 63, 73, 67, 92, 64, 68, 95, 119, 80, 72, 31, 43, 
    122, 111, 66, 77, 163, 108, 124, 79, 65, 64, 116, 75, 69, 49, 13, 
    128, 170, 80, 75, 197, 149, 158, 89, 65, 100, 153, 91, 76, 70, 32, 
    121, 179, 78, 67, 110, 142, 190, 125, 91, 136, 145, 80, 67, 81, 63, 
    151, 180, 73, 79, 75, 184, 163, 125, 87, 121, 146, 84, 75, 88, 63, 
    191, 194, 116, 131, 78, 113, 98, 97, 81, 85, 98, 78, 49, 65, 59, 
    208, 192, 150, 126, 110, 69, 104, 142, 75, 107, 81, 34, 51, 71, 73, 
    200, 181, 151, 159, 200, 105, 164, 199, 128, 67, 47, 65, 87, 107, 99, 
    160, 201, 160, 232, 251, 142, 116, 112, 103, 94, 101, 107, 115, 118, 117, 
    116, 135, 168, 259, 156, 105, 101, 96, 94, 96, 107, 115, 127, 130, 134, 
    126, 108, 139, 253, 120, 108, 104, 95, 102, 109, 118, 127, 122, 130, 150, 
    128, 118, 113, 134, 94, 102, 115, 108, 111, 118, 111, 107, 130, 155, 115, 
    
    -- channel=7
    62, 71, 67, 69, 69, 63, 69, 78, 73, 56, 48, 48, 56, 60, 65, 
    66, 71, 67, 73, 64, 70, 60, 63, 58, 24, 14, 11, 17, 37, 57, 
    55, 41, 70, 77, 68, 59, 71, 28, 1, 0, 7, 9, 17, 0, 41, 
    48, 0, 56, 68, 72, 36, 29, 10, 8, 0, 47, 9, 28, 8, 0, 
    29, 0, 56, 6, 34, 12, 40, 30, 19, 0, 14, 26, 7, 20, 0, 
    2, 0, 63, 65, 16, 30, 58, 23, 38, 0, 38, 37, 0, 13, 4, 
    0, 28, 23, 94, 3, 10, 26, 36, 34, 0, 42, 21, 0, 0, 10, 
    5, 24, 0, 44, 0, 0, 56, 22, 32, 0, 45, 28, 0, 5, 37, 
    18, 0, 32, 0, 22, 15, 28, 21, 0, 43, 1, 45, 1, 16, 35, 
    26, 0, 49, 0, 1, 5, 0, 22, 0, 22, 41, 0, 0, 18, 52, 
    0, 0, 46, 0, 47, 0, 0, 8, 18, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 53, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 19, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    0, 0, 3, 6, 7, 3, 1, 2, 7, 0, 0, 0, 0, 8, 12, 
    6, 9, 5, 6, 4, 44, 16, 0, 0, 4, 35, 18, 0, 0, 10, 
    0, 0, 4, 5, 4, 0, 0, 0, 9, 23, 23, 17, 37, 0, 0, 
    62, 21, 6, 4, 15, 1, 44, 23, 19, 0, 16, 2, 10, 16, 0, 
    39, 55, 11, 0, 69, 44, 19, 20, 14, 0, 33, 36, 26, 38, 0, 
    0, 0, 0, 0, 0, 0, 36, 33, 57, 1, 6, 0, 8, 26, 37, 
    0, 32, 0, 23, 0, 0, 4, 16, 34, 4, 4, 23, 17, 22, 28, 
    0, 27, 11, 27, 15, 0, 0, 0, 4, 2, 0, 17, 1, 0, 0, 
    4, 0, 14, 0, 13, 0, 0, 33, 1, 31, 0, 0, 0, 6, 20, 
    0, 0, 28, 15, 5, 0, 0, 65, 11, 0, 0, 5, 21, 21, 5, 
    0, 0, 20, 8, 96, 66, 3, 0, 0, 29, 37, 46, 27, 0, 0, 
    0, 0, 6, 27, 0, 0, 0, 0, 0, 12, 16, 17, 22, 23, 20, 
    29, 0, 0, 10, 0, 17, 20, 18, 23, 26, 29, 31, 18, 10, 28, 
    22, 18, 0, 0, 2, 19, 30, 22, 17, 21, 19, 8, 16, 23, 3, 
    28, 20, 10, 0, 9, 0, 0, 12, 30, 36, 30, 19, 36, 51, 31, 
    
    -- channel=9
    74, 72, 73, 75, 74, 66, 75, 81, 76, 64, 57, 60, 63, 65, 71, 
    73, 71, 72, 75, 74, 63, 59, 61, 54, 44, 25, 30, 44, 60, 69, 
    56, 72, 77, 78, 78, 70, 59, 46, 32, 24, 20, 26, 21, 35, 61, 
    31, 35, 71, 74, 65, 58, 34, 24, 27, 20, 35, 24, 35, 25, 44, 
    17, 8, 59, 49, 24, 7, 26, 29, 30, 21, 23, 21, 29, 27, 24, 
    7, 20, 58, 50, 38, 24, 32, 27, 30, 9, 24, 33, 26, 27, 19, 
    6, 13, 47, 75, 31, 28, 24, 31, 28, 10, 27, 26, 24, 24, 26, 
    1, 20, 6, 54, 26, 15, 39, 33, 40, 30, 33, 30, 21, 29, 52, 
    5, 6, 13, 21, 31, 31, 36, 31, 25, 39, 34, 44, 32, 44, 52, 
    27, 10, 21, 5, 14, 24, 27, 20, 12, 39, 38, 24, 16, 43, 59, 
    18, 11, 24, 5, 2, 0, 0, 15, 13, 21, 8, 0, 0, 11, 17, 
    0, 13, 11, 0, 12, 21, 6, 7, 3, 1, 0, 0, 0, 0, 0, 
    0, 0, 8, 12, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 39, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 16, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=10
    29, 42, 38, 40, 34, 40, 38, 39, 32, 16, 6, 15, 29, 25, 21, 
    37, 45, 41, 40, 44, 115, 23, 19, 0, 25, 25, 0, 0, 13, 24, 
    0, 15, 37, 41, 36, 47, 10, 0, 0, 75, 57, 49, 14, 0, 34, 
    15, 35, 33, 42, 31, 34, 65, 16, 22, 50, 62, 20, 16, 0, 15, 
    71, 111, 28, 56, 166, 77, 65, 27, 5, 44, 83, 26, 35, 14, 0, 
    29, 120, 41, 1, 115, 69, 119, 51, 26, 106, 68, 15, 33, 28, 4, 
    45, 105, 18, 30, 71, 107, 117, 71, 39, 114, 63, 25, 23, 51, 29, 
    71, 130, 12, 46, 47, 132, 55, 42, 39, 92, 75, 22, 30, 38, 40, 
    107, 123, 25, 91, 16, 26, 43, 52, 52, 24, 29, 0, 2, 52, 46, 
    131, 121, 74, 88, 42, 1, 67, 121, 13, 21, 0, 0, 37, 60, 31, 
    139, 109, 68, 168, 181, 71, 93, 89, 36, 0, 6, 27, 15, 2, 0, 
    39, 107, 106, 202, 73, 0, 8, 4, 12, 12, 25, 29, 45, 47, 41, 
    30, 29, 104, 147, 8, 36, 29, 27, 27, 32, 44, 50, 47, 44, 73, 
    39, 28, 36, 114, 31, 41, 38, 27, 32, 39, 36, 39, 38, 58, 33, 
    42, 43, 22, 29, 5, 17, 29, 39, 52, 59, 38, 40, 89, 84, 32, 
    
    -- channel=11
    0, 2, 0, 0, 0, 0, 0, 0, 0, 9, 23, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 45, 0, 0, 0, 11, 4, 0, 
    44, 30, 0, 0, 0, 65, 26, 12, 0, 0, 0, 0, 0, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 6, 17, 14, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 6, 
    3, 0, 0, 44, 73, 11, 0, 0, 0, 0, 14, 18, 0, 0, 0, 
    0, 20, 6, 9, 23, 0, 15, 0, 0, 0, 10, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 61, 41, 10, 4, 15, 6, 0, 21, 0, 
    0, 0, 1, 0, 0, 54, 1, 0, 0, 8, 34, 62, 24, 0, 0, 
    15, 0, 0, 0, 0, 4, 0, 0, 0, 53, 57, 3, 0, 0, 0, 
    0, 0, 16, 0, 0, 0, 0, 47, 18, 0, 0, 0, 0, 0, 2, 
    63, 23, 0, 0, 113, 76, 46, 39, 14, 4, 0, 2, 0, 0, 0, 
    0, 45, 0, 45, 73, 0, 1, 0, 0, 0, 0, 0, 4, 5, 0, 
    2, 0, 26, 101, 16, 0, 0, 0, 0, 0, 7, 16, 4, 0, 59, 
    6, 0, 12, 57, 27, 26, 28, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=12
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 7, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 19, 32, 24, 22, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 11, 20, 15, 14, 15, 19, 19, 0, 
    32, 28, 0, 0, 0, 0, 15, 16, 25, 6, 18, 16, 19, 21, 1, 
    39, 40, 0, 0, 22, 1, 16, 14, 26, 13, 23, 19, 21, 21, 20, 
    34, 52, 0, 0, 0, 0, 22, 12, 26, 26, 28, 25, 24, 24, 19, 
    37, 45, 19, 0, 0, 19, 23, 21, 15, 8, 19, 26, 24, 19, 0, 
    49, 56, 41, 24, 0, 13, 11, 18, 15, 0, 14, 15, 17, 0, 0, 
    37, 49, 48, 43, 35, 5, 8, 30, 27, 4, 18, 23, 23, 0, 0, 
    52, 40, 48, 36, 46, 46, 47, 51, 46, 35, 54, 62, 70, 61, 54, 
    106, 64, 42, 41, 69, 79, 86, 86, 90, 88, 98, 102, 108, 108, 107, 
    125, 97, 46, 60, 72, 94, 96, 93, 93, 99, 108, 112, 113, 111, 119, 
    130, 117, 86, 81, 79, 97, 98, 97, 97, 105, 114, 120, 119, 127, 133, 
    126, 123, 111, 99, 92, 99, 98, 95, 97, 106, 112, 109, 111, 131, 126, 
    
    -- channel=13
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 19, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 36, 34, 27, 15, 0, 0, 
    12, 23, 0, 0, 0, 0, 23, 24, 19, 15, 14, 7, 5, 3, 0, 
    35, 56, 0, 0, 56, 54, 19, 20, 8, 23, 33, 23, 24, 17, 0, 
    38, 32, 0, 0, 0, 0, 26, 24, 24, 60, 27, 4, 18, 23, 23, 
    48, 30, 0, 0, 0, 33, 18, 26, 14, 50, 14, 23, 23, 30, 24, 
    53, 41, 30, 0, 13, 36, 11, 0, 3, 30, 10, 13, 19, 14, 0, 
    55, 50, 37, 17, 28, 0, 0, 26, 20, 2, 0, 0, 3, 0, 0, 
    36, 49, 31, 44, 20, 22, 26, 49, 37, 0, 0, 1, 18, 2, 0, 
    38, 46, 23, 92, 91, 82, 62, 23, 20, 26, 48, 65, 57, 27, 20, 
    41, 34, 43, 88, 10, 2, 25, 26, 38, 54, 63, 67, 76, 78, 76, 
    87, 47, 50, 51, 12, 64, 62, 61, 64, 73, 81, 90, 78, 75, 99, 
    85, 74, 61, 12, 48, 71, 70, 65, 66, 76, 79, 73, 76, 103, 70, 
    88, 80, 64, 24, 51, 55, 54, 64, 78, 85, 79, 78, 105, 110, 74, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 0, 0, 24, 22, 10, 0, 0, 15, 0, 10, 0, 0, 
    58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 34, 4, 14, 0, 0, 
    22, 0, 0, 0, 0, 0, 44, 19, 21, 0, 2, 17, 0, 0, 0, 
    32, 8, 0, 13, 22, 0, 39, 6, 38, 0, 58, 35, 0, 0, 0, 
    0, 77, 0, 21, 0, 0, 47, 17, 41, 0, 58, 20, 0, 0, 0, 
    14, 43, 0, 2, 0, 0, 82, 25, 15, 0, 34, 37, 0, 0, 0, 
    46, 25, 62, 0, 6, 12, 14, 15, 0, 33, 16, 46, 0, 0, 0, 
    40, 22, 79, 0, 30, 0, 0, 21, 8, 15, 40, 0, 0, 0, 0, 
    4, 22, 87, 0, 27, 0, 0, 54, 42, 16, 0, 0, 0, 16, 30, 
    24, 7, 0, 0, 183, 84, 50, 45, 27, 13, 9, 14, 12, 13, 21, 
    30, 7, 0, 114, 117, 10, 16, 10, 9, 2, 1, 5, 20, 16, 0, 
    36, 12, 0, 154, 31, 5, 16, 11, 5, 9, 23, 27, 23, 4, 71, 
    45, 17, 20, 62, 31, 13, 14, 4, 0, 11, 26, 3, 0, 46, 44, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 26, 27, 12, 0, 0, 
    12, 0, 0, 0, 0, 0, 7, 16, 14, 0, 21, 3, 13, 0, 0, 
    55, 23, 0, 0, 38, 33, 22, 19, 5, 12, 26, 20, 14, 15, 0, 
    49, 29, 0, 0, 0, 19, 34, 20, 18, 18, 30, 18, 10, 21, 17, 
    60, 31, 0, 0, 0, 20, 20, 29, 20, 17, 32, 22, 15, 22, 13, 
    61, 52, 21, 0, 0, 13, 25, 7, 10, 0, 27, 16, 12, 5, 0, 
    68, 55, 45, 19, 5, 0, 7, 15, 12, 0, 0, 0, 0, 0, 0, 
    48, 51, 51, 38, 22, 11, 25, 41, 15, 0, 4, 6, 7, 0, 0, 
    38, 45, 45, 55, 101, 58, 45, 40, 41, 31, 39, 55, 46, 25, 24, 
    36, 49, 56, 52, 43, 45, 41, 43, 55, 59, 66, 71, 81, 80, 81, 
    89, 39, 54, 41, 59, 70, 68, 66, 67, 73, 83, 86, 81, 85, 99, 
    96, 79, 39, 47, 64, 72, 76, 67, 72, 78, 83, 80, 88, 97, 80, 
    97, 89, 72, 40, 57, 58, 63, 71, 79, 86, 82, 83, 100, 107, 93, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 18, 22, 0, 0, 0, 0, 0, 
    0, 72, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 12, 0, 65, 13, 0, 0, 0, 0, 95, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 122, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 31, 0, 0, 0, 27, 0, 0, 0, 14, 0, 
    0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 5, 0, 0, 0, 0, 28, 0, 0, 0, 0, 14, 0, 
    0, 0, 0, 20, 0, 0, 42, 0, 0, 0, 0, 0, 31, 0, 0, 
    0, 0, 0, 129, 3, 0, 0, 0, 0, 0, 35, 39, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 62, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 0, 0, 
    
    -- channel=17
    1, 0, 0, 0, 5, 3, 0, 3, 11, 10, 8, 4, 3, 2, 5, 
    5, 3, 0, 0, 0, 0, 18, 9, 23, 30, 31, 36, 29, 6, 1, 
    5, 1, 6, 3, 8, 18, 31, 55, 21, 4, 0, 0, 8, 13, 0, 
    25, 14, 9, 10, 19, 34, 8, 0, 0, 0, 0, 5, 7, 0, 0, 
    6, 0, 5, 9, 0, 6, 7, 1, 2, 18, 14, 5, 0, 0, 16, 
    21, 0, 0, 39, 0, 2, 0, 7, 6, 0, 0, 8, 0, 0, 2, 
    16, 6, 10, 9, 5, 7, 0, 5, 0, 0, 15, 15, 18, 4, 0, 
    15, 1, 22, 24, 9, 0, 0, 2, 0, 0, 3, 19, 0, 0, 0, 
    9, 5, 18, 0, 25, 31, 25, 15, 0, 68, 5, 1, 5, 0, 0, 
    0, 0, 0, 33, 0, 1, 18, 3, 8, 0, 1, 11, 0, 0, 15, 
    12, 14, 20, 0, 0, 0, 0, 0, 0, 40, 27, 5, 17, 48, 58, 
    7, 0, 0, 0, 37, 46, 53, 48, 17, 13, 3, 11, 7, 7, 7, 
    7, 10, 4, 10, 27, 2, 1, 6, 8, 5, 6, 1, 0, 4, 2, 
    1, 9, 2, 0, 4, 5, 10, 4, 0, 0, 8, 1, 12, 0, 0, 
    0, 0, 23, 26, 18, 1, 0, 0, 0, 7, 5, 4, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    17, 14, 0, 11, 41, 21, 0, 0, 0, 7, 10, 0, 0, 0, 0, 
    15, 1, 0, 0, 6, 9, 9, 0, 0, 18, 0, 0, 0, 0, 0, 
    21, 0, 0, 0, 0, 26, 20, 0, 0, 21, 0, 0, 0, 0, 0, 
    25, 22, 0, 0, 0, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 32, 0, 3, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 
    17, 26, 0, 30, 0, 0, 11, 10, 0, 0, 0, 0, 0, 0, 0, 
    22, 25, 4, 51, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 32, 46, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 42, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    11, 7, 9, 10, 10, 6, 12, 11, 7, 7, 6, 6, 7, 7, 7, 
    13, 8, 8, 11, 10, 11, 7, 4, 3, 1, 5, 2, 2, 11, 10, 
    1, 16, 13, 10, 12, 0, 2, 0, 0, 4, 0, 0, 6, 7, 13, 
    0, 17, 18, 9, 4, 2, 4, 0, 7, 4, 2, 0, 0, 5, 12, 
    0, 18, 14, 0, 6, 0, 0, 0, 1, 3, 0, 0, 1, 4, 1, 
    0, 11, 13, 0, 0, 0, 2, 0, 3, 7, 0, 0, 1, 1, 2, 
    0, 12, 12, 4, 0, 2, 3, 3, 0, 10, 0, 0, 2, 5, 6, 
    0, 0, 2, 13, 5, 4, 0, 1, 2, 5, 4, 0, 0, 6, 6, 
    0, 0, 0, 10, 4, 0, 0, 2, 7, 8, 0, 0, 0, 10, 13, 
    0, 0, 2, 3, 0, 0, 0, 8, 0, 0, 1, 0, 11, 17, 10, 
    11, 0, 0, 0, 14, 2, 6, 0, 0, 0, 0, 5, 2, 11, 10, 
    5, 6, 3, 14, 0, 0, 0, 0, 0, 2, 6, 3, 3, 5, 3, 
    11, 4, 3, 8, 0, 1, 1, 2, 3, 4, 4, 4, 5, 2, 4, 
    6, 7, 0, 8, 2, 1, 3, 1, 1, 1, 3, 4, 5, 3, 10, 
    5, 3, 9, 0, 5, 3, 4, 4, 3, 3, 3, 3, 6, 5, 7, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 2, 0, 0, 1, 4, 
    0, 0, 0, 0, 0, 0, 32, 6, 17, 0, 18, 17, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 43, 19, 0, 0, 32, 15, 54, 0, 0, 
    123, 0, 0, 0, 18, 0, 17, 30, 12, 0, 60, 11, 40, 38, 0, 
    98, 0, 45, 0, 0, 11, 62, 52, 35, 0, 18, 74, 1, 53, 0, 
    71, 0, 58, 0, 0, 2, 54, 46, 85, 0, 78, 77, 0, 28, 31, 
    59, 54, 5, 58, 0, 0, 25, 42, 89, 0, 91, 57, 0, 0, 38, 
    46, 39, 41, 34, 0, 0, 92, 13, 44, 0, 47, 68, 0, 0, 8, 
    54, 0, 120, 0, 27, 0, 27, 17, 0, 32, 0, 70, 0, 0, 0, 
    1, 0, 130, 0, 70, 0, 0, 32, 27, 15, 65, 6, 0, 0, 11, 
    0, 0, 117, 0, 114, 52, 0, 25, 89, 45, 1, 0, 0, 0, 19, 
    0, 0, 30, 0, 156, 71, 2, 6, 25, 6, 4, 0, 0, 4, 18, 
    38, 0, 0, 32, 144, 9, 18, 10, 12, 3, 0, 0, 10, 2, 0, 
    45, 7, 0, 101, 42, 0, 27, 14, 1, 1, 6, 6, 15, 0, 41, 
    56, 7, 2, 14, 26, 0, 0, 7, 0, 7, 29, 0, 0, 39, 79, 
    
    -- channel=21
    3, 0, 6, 0, 0, 5, 0, 0, 0, 0, 0, 6, 2, 0, 0, 
    3, 3, 9, 0, 12, 14, 0, 0, 0, 19, 0, 0, 9, 11, 0, 
    0, 28, 4, 0, 10, 0, 0, 0, 23, 59, 0, 0, 0, 21, 12, 
    0, 85, 0, 11, 0, 27, 0, 0, 0, 83, 0, 0, 0, 0, 59, 
    0, 40, 0, 95, 0, 19, 0, 0, 0, 115, 0, 0, 0, 0, 42, 
    0, 1, 0, 35, 44, 1, 0, 0, 0, 198, 0, 0, 13, 0, 0, 
    0, 0, 0, 0, 66, 67, 0, 0, 0, 148, 0, 0, 10, 21, 0, 
    0, 0, 0, 0, 70, 75, 0, 0, 0, 89, 0, 0, 29, 2, 0, 
    0, 2, 0, 25, 7, 3, 0, 0, 31, 0, 14, 0, 22, 15, 17, 
    0, 5, 0, 66, 0, 25, 46, 0, 3, 0, 0, 0, 42, 39, 0, 
    51, 5, 0, 172, 0, 0, 71, 0, 0, 0, 15, 34, 32, 17, 0, 
    61, 32, 0, 118, 0, 0, 0, 0, 0, 6, 7, 10, 8, 8, 0, 
    0, 67, 102, 0, 0, 0, 0, 0, 0, 10, 14, 15, 3, 9, 18, 
    0, 8, 152, 0, 0, 10, 0, 1, 10, 10, 7, 2, 0, 37, 0, 
    0, 4, 18, 0, 0, 17, 4, 0, 17, 3, 0, 9, 52, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=23
    50, 57, 55, 57, 57, 51, 59, 65, 64, 55, 50, 48, 53, 54, 56, 
    59, 60, 55, 61, 53, 51, 63, 61, 58, 25, 24, 19, 19, 42, 53, 
    50, 42, 58, 63, 53, 22, 63, 26, 11, 0, 5, 15, 29, 7, 40, 
    55, 0, 56, 58, 64, 32, 29, 18, 13, 0, 41, 8, 28, 22, 5, 
    50, 0, 64, 14, 42, 13, 31, 28, 17, 0, 15, 35, 9, 35, 0, 
    5, 0, 70, 21, 0, 22, 47, 27, 39, 0, 30, 40, 0, 21, 22, 
    9, 17, 40, 81, 0, 0, 22, 35, 42, 0, 42, 24, 0, 0, 19, 
    8, 22, 15, 57, 0, 0, 36, 12, 32, 0, 34, 24, 0, 0, 33, 
    11, 0, 34, 7, 16, 0, 24, 14, 0, 25, 0, 39, 0, 11, 31, 
    3, 0, 52, 0, 22, 5, 0, 24, 0, 26, 44, 14, 0, 26, 59, 
    0, 0, 41, 0, 68, 4, 0, 13, 44, 25, 0, 0, 0, 0, 0, 
    0, 0, 15, 0, 32, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 5, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 5, 9, 0, 
    0, 47, 0, 0, 0, 45, 0, 0, 0, 14, 0, 0, 0, 19, 3, 
    0, 5, 0, 0, 0, 0, 0, 0, 0, 84, 0, 6, 0, 0, 51, 
    0, 0, 0, 48, 0, 0, 0, 0, 0, 58, 0, 0, 0, 0, 18, 
    0, 21, 0, 0, 115, 34, 0, 0, 0, 94, 0, 0, 14, 0, 0, 
    0, 0, 21, 0, 61, 17, 11, 0, 0, 92, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 31, 81, 0, 28, 0, 66, 0, 0, 24, 14, 0, 
    0, 22, 0, 25, 0, 59, 0, 0, 19, 0, 42, 0, 19, 5, 0, 
    21, 29, 0, 33, 0, 8, 22, 0, 0, 41, 0, 0, 9, 4, 0, 
    63, 18, 0, 79, 0, 0, 49, 46, 0, 0, 0, 0, 6, 24, 2, 
    135, 81, 0, 64, 4, 33, 42, 41, 16, 14, 16, 18, 11, 17, 11, 
    0, 110, 97, 16, 0, 7, 7, 9, 7, 8, 10, 9, 23, 31, 11, 
    5, 16, 160, 9, 2, 15, 0, 7, 18, 16, 20, 35, 17, 27, 37, 
    0, 19, 25, 58, 15, 44, 45, 16, 8, 0, 1, 19, 22, 0, 0, 
    
    -- channel=25
    15, 12, 21, 17, 19, 19, 13, 17, 21, 5, 0, 11, 19, 12, 15, 
    24, 19, 20, 12, 29, 48, 0, 2, 0, 46, 21, 10, 14, 22, 15, 
    0, 28, 20, 18, 19, 0, 0, 16, 38, 48, 0, 11, 0, 12, 24, 
    0, 75, 10, 29, 6, 57, 8, 0, 3, 29, 0, 0, 0, 0, 41, 
    0, 18, 0, 92, 23, 6, 0, 0, 0, 98, 8, 0, 15, 0, 15, 
    0, 0, 0, 0, 6, 2, 0, 0, 0, 120, 0, 0, 12, 5, 15, 
    14, 0, 6, 0, 19, 57, 0, 0, 0, 66, 0, 0, 20, 31, 0, 
    3, 0, 4, 5, 39, 0, 0, 0, 0, 28, 0, 0, 21, 0, 13, 
    0, 0, 0, 27, 4, 0, 3, 4, 41, 0, 0, 0, 18, 32, 17, 
    0, 0, 0, 48, 0, 14, 64, 0, 0, 0, 0, 17, 30, 23, 5, 
    27, 0, 0, 126, 0, 0, 0, 0, 0, 5, 39, 35, 14, 15, 10, 
    0, 14, 0, 32, 0, 0, 0, 0, 0, 7, 4, 5, 11, 1, 0, 
    0, 0, 82, 0, 0, 5, 0, 1, 5, 11, 16, 11, 0, 0, 27, 
    0, 0, 34, 0, 0, 9, 0, 0, 5, 5, 0, 0, 0, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 11, 10, 0, 12, 47, 0, 0, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 14, 10, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 29, 0, 0, 53, 20, 0, 0, 0, 8, 12, 0, 0, 0, 0, 
    0, 33, 0, 0, 25, 0, 45, 0, 0, 38, 2, 0, 0, 0, 0, 
    0, 26, 0, 0, 2, 61, 22, 10, 0, 25, 0, 0, 0, 1, 0, 
    19, 41, 0, 9, 0, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 39, 0, 19, 1, 0, 0, 5, 0, 1, 0, 0, 0, 0, 0, 
    41, 30, 2, 22, 0, 0, 46, 54, 4, 0, 0, 0, 0, 0, 0, 
    61, 47, 24, 73, 61, 0, 2, 0, 0, 0, 0, 0, 0, 3, 0, 
    0, 39, 25, 67, 0, 0, 0, 0, 0, 0, 0, 0, 12, 10, 1, 
    0, 1, 50, 51, 0, 0, 0, 0, 0, 0, 3, 9, 0, 0, 32, 
    3, 4, 3, 22, 0, 0, 7, 0, 0, 0, 0, 0, 4, 16, 0, 
    
    -- channel=28
    2, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 4, 9, 0, 
    0, 40, 0, 0, 0, 50, 0, 0, 0, 0, 0, 0, 0, 14, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 0, 5, 0, 0, 37, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 11, 
    0, 0, 0, 16, 102, 13, 0, 0, 0, 29, 0, 0, 1, 0, 0, 
    0, 0, 12, 0, 42, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 40, 0, 20, 0, 43, 0, 0, 9, 15, 1, 
    0, 0, 0, 0, 0, 46, 0, 0, 0, 0, 46, 8, 25, 10, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 38, 0, 0, 0, 0, 0, 
    14, 0, 0, 1, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 
    75, 26, 0, 0, 0, 20, 21, 20, 0, 0, 0, 0, 0, 0, 0, 
    0, 60, 18, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 83, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 35, 0, 16, 13, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 0, 0, 2, 0, 0, 
    8, 0, 0, 0, 0, 20, 23, 19, 0, 0, 9, 1, 8, 0, 0, 
    19, 0, 0, 0, 0, 0, 0, 3, 2, 0, 16, 18, 26, 15, 0, 
    7, 0, 0, 0, 0, 0, 18, 17, 22, 0, 0, 12, 0, 11, 0, 
    16, 0, 1, 20, 31, 23, 7, 9, 16, 0, 12, 30, 2, 6, 0, 
    6, 11, 5, 24, 0, 0, 9, 1, 27, 0, 27, 15, 1, 0, 3, 
    1, 9, 0, 0, 0, 0, 26, 24, 22, 0, 21, 28, 4, 9, 11, 
    2, 0, 22, 0, 0, 34, 25, 4, 0, 6, 31, 45, 15, 0, 0, 
    9, 0, 30, 0, 20, 0, 0, 0, 0, 28, 34, 20, 0, 0, 0, 
    0, 0, 34, 0, 0, 0, 0, 17, 16, 4, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 67, 60, 35, 35, 21, 5, 1, 3, 1, 2, 7, 
    0, 2, 0, 6, 67, 7, 11, 9, 8, 1, 0, 0, 1, 3, 0, 
    10, 0, 0, 48, 18, 0, 5, 9, 7, 3, 4, 11, 9, 0, 21, 
    12, 8, 6, 38, 17, 15, 14, 5, 0, 0, 9, 4, 0, 0, 19, 
    
    -- channel=30
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 0, 0, 0, 
    0, 29, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 49, 0, 1, 49, 22, 0, 0, 0, 32, 18, 0, 0, 0, 0, 
    0, 26, 0, 0, 0, 0, 21, 0, 0, 84, 0, 0, 0, 0, 0, 
    10, 0, 0, 0, 0, 46, 0, 0, 0, 58, 0, 0, 0, 9, 0, 
    21, 24, 0, 0, 0, 14, 0, 0, 0, 34, 0, 0, 0, 0, 0, 
    27, 31, 0, 12, 0, 0, 0, 2, 4, 0, 0, 0, 0, 4, 0, 
    24, 33, 0, 42, 0, 0, 23, 28, 0, 0, 0, 0, 0, 0, 0, 
    33, 25, 0, 131, 75, 27, 10, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 10, 12, 102, 0, 0, 0, 0, 0, 0, 0, 4, 18, 22, 11, 
    10, 0, 53, 10, 0, 8, 0, 2, 4, 13, 23, 29, 8, 5, 48, 
    9, 10, 17, 0, 0, 15, 12, 4, 4, 14, 11, 5, 10, 43, 0, 
    9, 19, 4, 0, 0, 0, 0, 5, 23, 33, 11, 21, 67, 42, 0, 
    
    -- channel=31
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 1, 7, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 3, 7, 3, 0, 6, 1, 6, 0, 
    6, 10, 0, 0, 0, 0, 2, 4, 11, 0, 0, 5, 1, 5, 0, 
    21, 20, 0, 0, 5, 0, 0, 0, 9, 0, 16, 1, 4, 3, 0, 
    6, 39, 0, 0, 0, 0, 20, 0, 12, 7, 9, 6, 0, 3, 6, 
    16, 17, 0, 0, 0, 28, 13, 6, 0, 0, 2, 6, 7, 11, 0, 
    26, 30, 27, 3, 0, 0, 0, 4, 0, 0, 13, 1, 0, 0, 0, 
    18, 26, 29, 4, 29, 0, 0, 13, 15, 10, 5, 2, 3, 0, 0, 
    29, 20, 24, 3, 20, 36, 49, 45, 35, 6, 24, 38, 44, 31, 30, 
    81, 36, 17, 27, 68, 44, 47, 47, 56, 58, 67, 67, 71, 73, 74, 
    90, 70, 9, 61, 39, 61, 65, 60, 61, 66, 70, 77, 83, 77, 75, 
    92, 79, 65, 67, 53, 61, 63, 65, 66, 72, 80, 86, 78, 91, 109, 
    92, 85, 77, 59, 63, 70, 72, 63, 64, 67, 78, 69, 68, 96, 87, 
    
    
    others => 0);
end gold_package;
