library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package iwght_package is
  type mem is array(0 to 4000000) of integer;

  constant input_wght : mem := (
    -- bias
    1667, -2120, 7432, 241, -3858, -5338, -7391, -9255, -5555, -10569, 8651, -10870, -4125, 4217, -4600, -428, 1219, -1023, -2754, -941, 89, -575, -4742, -4741, -3326, -2324, 10239, 3129, -4241, -1941, -8043, -2158, -1838, -5539, -3575, -4860, 2573, 1278, -3056, -1078, -586, -6735, -3412, 8011, -4375, -1911, 4223, -1340, -9774, -1503, -5391, 10268, -2565, 19, -19, 1739, -7715, 5495, -166, -5499, 17173, -8026, 3916, -6577,

    -- weights
    -- filter=0 channel=0
    -8, -14, 3, 3, -3, -4, -7, -5, -8,
    -- filter=0 channel=1
    3, 11, 0, 6, -15, -16, -8, 10, 7,
    -- filter=0 channel=2
    -2, 1, 4, 9, -13, 1, 9, 9, 10,
    -- filter=0 channel=3
    -13, 4, -8, 4, 14, -9, 3, -11, 13,
    -- filter=0 channel=4
    10, 9, 2, -5, 12, 12, -8, 6, 0,
    -- filter=0 channel=5
    -6, 3, -7, -10, 5, 12, 5, 10, -14,
    -- filter=0 channel=6
    8, -8, 13, -3, -11, 1, -11, -1, -14,
    -- filter=0 channel=7
    18, 1, -22, 13, 3, -14, 9, 3, -7,
    -- filter=0 channel=8
    6, 5, 1, -3, 16, -9, -8, 0, -10,
    -- filter=0 channel=9
    -9, 11, -11, -13, 2, 13, -7, -6, 0,
    -- filter=0 channel=10
    -3, -10, -2, -2, -12, -4, -2, 4, 15,
    -- filter=0 channel=11
    -10, 7, -2, -5, -1, 4, -14, 0, -7,
    -- filter=0 channel=12
    15, 9, -20, 0, -4, -14, 6, -14, -7,
    -- filter=0 channel=13
    -8, 5, -10, 16, -9, -12, -2, -4, -14,
    -- filter=0 channel=14
    5, -3, -4, -14, -6, -13, 6, 4, 13,
    -- filter=0 channel=15
    9, 13, 8, 12, 6, 0, 14, -6, -14,
    -- filter=0 channel=16
    -3, 3, -1, -8, 13, 9, -10, 0, -15,
    -- filter=0 channel=17
    24, 16, -9, 19, 1, -4, 21, -7, -9,
    -- filter=0 channel=18
    -1, -5, -10, -9, -7, -8, -6, 2, 11,
    -- filter=0 channel=19
    -1, -5, -5, -7, 14, 7, -3, 3, 5,
    -- filter=0 channel=20
    -9, -16, -10, -6, -7, -11, -6, 7, -20,
    -- filter=0 channel=21
    5, 12, -2, 3, -12, -8, 20, -5, 1,
    -- filter=0 channel=22
    -6, -3, 12, 1, 5, 7, -9, 7, 12,
    -- filter=0 channel=23
    2, 10, -9, 8, -11, 16, 11, -6, -1,
    -- filter=0 channel=24
    -4, 2, 10, -7, -13, -15, -7, 10, -6,
    -- filter=0 channel=25
    -11, -4, 6, 0, 2, -4, -8, -5, 6,
    -- filter=0 channel=26
    16, 11, 0, 12, 0, -2, 8, -2, 12,
    -- filter=0 channel=27
    -7, 12, -6, -7, 13, -1, -1, 14, 4,
    -- filter=0 channel=28
    7, -2, 0, -6, -11, 7, 5, 1, -2,
    -- filter=0 channel=29
    4, 16, 18, 15, 0, 16, -4, 2, 6,
    -- filter=0 channel=30
    -6, -5, -13, -6, -7, -12, 6, -6, -2,
    -- filter=0 channel=31
    7, -9, -15, 12, 4, -11, -5, -15, 6,
    -- filter=1 channel=0
    7, 15, 11, 12, 3, 1, -10, 0, 0,
    -- filter=1 channel=1
    9, -13, 1, -3, -9, -3, 2, 8, 0,
    -- filter=1 channel=2
    5, 11, 5, -2, 1, 11, 8, 3, 0,
    -- filter=1 channel=3
    3, -1, -5, 6, -12, -7, -13, -7, -4,
    -- filter=1 channel=4
    1, -14, 7, 0, -17, -5, 9, -9, 0,
    -- filter=1 channel=5
    -11, -14, -7, -2, 11, -4, -14, 5, -13,
    -- filter=1 channel=6
    3, 12, 0, -7, 13, -11, 3, 6, 12,
    -- filter=1 channel=7
    1, -11, 17, 8, -4, 14, 9, 9, 3,
    -- filter=1 channel=8
    -14, 12, -9, -15, 8, 9, -10, 10, 5,
    -- filter=1 channel=9
    5, -10, 12, -9, -5, 15, 3, 9, 7,
    -- filter=1 channel=10
    7, -1, 13, 9, 3, 8, -9, -2, -10,
    -- filter=1 channel=11
    -12, 7, -7, 10, 5, 8, 0, 0, 11,
    -- filter=1 channel=12
    17, 16, -2, -11, 2, 10, -13, 10, 10,
    -- filter=1 channel=13
    5, 0, 14, 5, -12, -4, 13, 4, 0,
    -- filter=1 channel=14
    -7, -6, -7, -7, 9, 10, -13, -15, 8,
    -- filter=1 channel=15
    -8, 4, -7, 8, 2, -7, -1, 0, -8,
    -- filter=1 channel=16
    9, -3, 0, -9, -5, -10, -8, 11, 13,
    -- filter=1 channel=17
    1, -6, 8, 3, 6, 13, 2, -15, -13,
    -- filter=1 channel=18
    -16, -14, -5, 4, -9, -7, -2, -14, 6,
    -- filter=1 channel=19
    -6, 8, 3, 14, -5, 12, -1, 8, -4,
    -- filter=1 channel=20
    -2, -10, -7, 8, -2, 3, 7, 3, -3,
    -- filter=1 channel=21
    11, -3, 5, -12, -6, 8, 3, -13, -6,
    -- filter=1 channel=22
    4, 9, 16, 6, 6, 10, 0, 5, 22,
    -- filter=1 channel=23
    -15, -9, 5, 5, -13, 11, 6, 9, 10,
    -- filter=1 channel=24
    -9, 6, -9, -14, 0, -4, -6, -2, 15,
    -- filter=1 channel=25
    -15, -21, 1, -14, 7, 7, -2, -9, -9,
    -- filter=1 channel=26
    9, -6, -6, -2, -6, 0, -11, -9, -15,
    -- filter=1 channel=27
    13, 8, -1, 1, -11, 9, 12, 1, 4,
    -- filter=1 channel=28
    5, 7, 16, 5, -3, -10, -6, -1, 14,
    -- filter=1 channel=29
    0, -1, 9, 2, -14, -1, -3, 3, 14,
    -- filter=1 channel=30
    2, -12, -9, 14, 5, 12, -2, 4, 7,
    -- filter=1 channel=31
    4, 11, -12, 15, 10, 5, -6, -8, -14,
    -- filter=2 channel=0
    8, 6, 13, 5, -10, -11, 13, 4, -10,
    -- filter=2 channel=1
    -17, -15, 0, 0, -4, 5, -17, 10, 11,
    -- filter=2 channel=2
    7, 1, 10, 0, -9, 0, -7, 8, 7,
    -- filter=2 channel=3
    0, -13, 9, 7, -1, 6, 11, -2, -14,
    -- filter=2 channel=4
    2, -8, 3, -6, 0, 9, -3, 4, 14,
    -- filter=2 channel=5
    -8, 11, 9, -15, -10, 10, -16, 6, -8,
    -- filter=2 channel=6
    -4, -11, 1, 0, -13, 4, -14, 1, -8,
    -- filter=2 channel=7
    11, -1, 12, 10, 16, 13, 8, 16, 12,
    -- filter=2 channel=8
    -6, 10, 10, -4, -13, 9, -1, -9, -12,
    -- filter=2 channel=9
    -11, 7, -13, -12, -13, 0, -2, -3, -3,
    -- filter=2 channel=10
    -6, -1, 2, -9, -1, -8, -3, 7, -4,
    -- filter=2 channel=11
    6, 11, -8, 17, 2, -9, 14, 7, -15,
    -- filter=2 channel=12
    7, -12, 14, 3, 3, 5, 0, 2, -5,
    -- filter=2 channel=13
    4, 0, -15, -20, -6, -11, 0, -13, 0,
    -- filter=2 channel=14
    -8, 6, 15, -5, 5, 14, 7, -3, 12,
    -- filter=2 channel=15
    5, -5, 0, -10, -15, 8, -13, 3, 5,
    -- filter=2 channel=16
    -4, 3, -11, -5, -4, -2, -10, -6, -15,
    -- filter=2 channel=17
    -7, -16, -3, -20, -19, -13, 5, 10, -1,
    -- filter=2 channel=18
    3, -2, -6, -5, 4, 0, -16, 0, 2,
    -- filter=2 channel=19
    12, 0, -12, -4, 14, 12, -2, 10, 14,
    -- filter=2 channel=20
    -3, 14, 6, -15, -1, 10, -9, -7, 16,
    -- filter=2 channel=21
    -17, -15, -5, -3, 2, 4, 4, 7, -8,
    -- filter=2 channel=22
    4, -1, 16, 0, -12, 8, 8, 1, -9,
    -- filter=2 channel=23
    2, 3, -12, 10, 0, 3, -9, 8, 7,
    -- filter=2 channel=24
    4, -11, 3, -9, 0, -9, 5, 0, 2,
    -- filter=2 channel=25
    -18, 7, 6, 2, 11, 10, -8, 15, 22,
    -- filter=2 channel=26
    4, -21, -16, -18, -1, -19, 1, -16, -15,
    -- filter=2 channel=27
    -3, 14, 0, -11, -7, -5, -12, -5, 4,
    -- filter=2 channel=28
    -5, -11, 12, -1, -3, -5, -7, -3, 4,
    -- filter=2 channel=29
    16, -5, 5, 5, -1, 1, 10, -10, -7,
    -- filter=2 channel=30
    -5, -12, -1, 8, -13, -5, 4, -1, 14,
    -- filter=2 channel=31
    -14, -7, 5, -6, -16, -11, -17, -4, -10,
    -- filter=3 channel=0
    4, 15, 8, 10, 9, -13, 9, -5, 12,
    -- filter=3 channel=1
    -8, 11, 9, 7, 2, 3, 0, -6, 2,
    -- filter=3 channel=2
    6, -8, -13, 6, 14, -6, -11, 5, -9,
    -- filter=3 channel=3
    -5, -2, 0, 12, 10, 1, -9, 8, 0,
    -- filter=3 channel=4
    3, 10, -5, -6, 3, -15, -11, -15, -7,
    -- filter=3 channel=5
    -9, -8, 11, 8, -15, 5, 14, -11, 4,
    -- filter=3 channel=6
    -2, 2, 11, -4, -11, 12, -10, 5, 0,
    -- filter=3 channel=7
    -14, -3, -7, -10, 1, -10, 16, -6, 17,
    -- filter=3 channel=8
    0, -5, 6, 7, -5, -2, 6, -3, 4,
    -- filter=3 channel=9
    8, -6, 8, -5, -1, 6, 4, -13, 10,
    -- filter=3 channel=10
    6, 12, 14, -5, -7, -9, -2, 9, -13,
    -- filter=3 channel=11
    1, 12, -8, 0, 9, 7, -8, -14, -7,
    -- filter=3 channel=12
    2, -11, -9, -4, 7, 4, 10, 4, -4,
    -- filter=3 channel=13
    -18, -20, 0, -14, -4, 3, 8, 11, 15,
    -- filter=3 channel=14
    0, -10, -2, -8, -1, -12, 12, 4, -4,
    -- filter=3 channel=15
    4, -9, 4, -9, -6, -4, 12, -9, -2,
    -- filter=3 channel=16
    0, -12, 16, -8, -6, 2, 14, 15, 6,
    -- filter=3 channel=17
    -12, -14, -12, -17, -5, 9, 12, 4, 20,
    -- filter=3 channel=18
    14, 10, 6, 13, 0, -15, -16, -16, 0,
    -- filter=3 channel=19
    -4, -13, -13, 13, 10, -11, 12, 0, 13,
    -- filter=3 channel=20
    -16, -17, -18, -12, 9, 0, 2, 3, 17,
    -- filter=3 channel=21
    6, 2, 10, -4, -5, -7, 11, 16, -3,
    -- filter=3 channel=22
    12, -3, 13, 7, 6, -11, -6, 0, -2,
    -- filter=3 channel=23
    -7, 1, 12, -12, 3, -15, -12, 10, 8,
    -- filter=3 channel=24
    9, -3, 8, 0, -4, 9, -14, 14, -8,
    -- filter=3 channel=25
    1, 6, 2, 10, 4, 0, 8, -1, 10,
    -- filter=3 channel=26
    2, -6, 13, 5, 6, -6, 0, 16, 3,
    -- filter=3 channel=27
    -7, -7, -1, -14, -5, -14, -5, 2, 14,
    -- filter=3 channel=28
    -4, -4, 13, -10, 13, -8, 1, -9, 17,
    -- filter=3 channel=29
    -8, 3, -1, -1, -5, 1, -6, 3, -12,
    -- filter=3 channel=30
    -1, 1, -7, -1, 8, 14, -12, -1, 4,
    -- filter=3 channel=31
    -5, -16, 11, 3, 3, 12, -8, 14, -11,
    -- filter=4 channel=0
    -12, -4, 0, -10, -4, 6, 18, -5, -4,
    -- filter=4 channel=1
    7, 14, 12, -5, 9, 6, 4, 9, -7,
    -- filter=4 channel=2
    7, -14, 9, -8, -6, -11, -10, -5, -6,
    -- filter=4 channel=3
    7, -3, -5, -12, 12, 4, -8, -3, -9,
    -- filter=4 channel=4
    -1, 14, -6, 8, -11, -9, -6, 3, 2,
    -- filter=4 channel=5
    -3, -8, 13, -9, 0, -9, 1, -14, -12,
    -- filter=4 channel=6
    -12, 3, -2, 6, -7, -7, 8, -2, -4,
    -- filter=4 channel=7
    8, 11, 0, -8, 1, 1, -6, 10, -2,
    -- filter=4 channel=8
    5, -6, -8, 5, -7, 5, 9, -1, 0,
    -- filter=4 channel=9
    10, 11, 17, 6, 17, 12, 17, 17, -10,
    -- filter=4 channel=10
    9, 5, 6, 0, 9, 9, 12, 9, -8,
    -- filter=4 channel=11
    0, 7, -9, -7, 3, 1, -9, -4, -4,
    -- filter=4 channel=12
    -5, 17, 14, -2, 3, -5, 8, 0, 15,
    -- filter=4 channel=13
    0, 4, 9, 0, -14, 1, -6, -6, 1,
    -- filter=4 channel=14
    11, 4, -3, 10, -14, 11, -2, -3, -7,
    -- filter=4 channel=15
    -13, 13, -5, -15, 11, 6, -10, -7, -8,
    -- filter=4 channel=16
    -5, 11, 0, 2, -14, -11, 7, 14, -15,
    -- filter=4 channel=17
    14, 15, 0, -9, 10, 0, -18, 0, -3,
    -- filter=4 channel=18
    -12, 7, -9, -7, 0, -10, 0, -10, 8,
    -- filter=4 channel=19
    -4, 11, -6, 2, 2, 12, 10, 3, -11,
    -- filter=4 channel=20
    16, 13, 1, -3, 11, 0, -15, -10, -12,
    -- filter=4 channel=21
    -3, 7, 5, 8, -10, -13, -20, -1, -18,
    -- filter=4 channel=22
    19, 17, 23, 20, 18, 20, 22, 27, 26,
    -- filter=4 channel=23
    6, -3, 6, 14, 1, -1, 16, 15, 4,
    -- filter=4 channel=24
    -9, -4, -7, 12, -11, -14, 13, -13, 11,
    -- filter=4 channel=25
    4, -4, -5, -15, 0, -13, -5, 8, 0,
    -- filter=4 channel=26
    0, 9, -5, 10, 0, -2, 6, -13, -15,
    -- filter=4 channel=27
    5, 2, -5, -8, -4, -5, -4, -8, -4,
    -- filter=4 channel=28
    -4, -3, -11, 6, -7, 5, -11, -7, -4,
    -- filter=4 channel=29
    2, -9, 7, 12, 13, 8, 1, 9, 10,
    -- filter=4 channel=30
    2, 9, 3, 12, -7, -12, -1, -10, -4,
    -- filter=4 channel=31
    3, -6, 13, 12, 6, 3, -17, -8, -16,
    -- filter=5 channel=0
    8, -12, 0, 3, -12, -14, 10, -13, -14,
    -- filter=5 channel=1
    6, -13, 6, -2, 0, 8, -5, -1, -14,
    -- filter=5 channel=2
    5, -7, -8, 6, -3, 13, -5, -9, 9,
    -- filter=5 channel=3
    -10, -1, -1, -11, 5, 3, 6, -8, 5,
    -- filter=5 channel=4
    17, 21, 2, -1, 6, 8, 13, 11, 20,
    -- filter=5 channel=5
    -12, 14, -12, 8, -14, 8, -14, -4, -3,
    -- filter=5 channel=6
    -6, 12, -4, 11, -7, -11, -4, -11, 6,
    -- filter=5 channel=7
    10, -3, 1, 2, -13, -20, -8, 4, -21,
    -- filter=5 channel=8
    0, -7, -7, 9, 9, -14, 3, 4, 11,
    -- filter=5 channel=9
    7, 8, 11, 13, -11, -15, 7, 11, 12,
    -- filter=5 channel=10
    -1, -3, -9, -4, -12, 9, 3, 10, 15,
    -- filter=5 channel=11
    -6, -17, -17, -8, -8, -18, 7, -16, 10,
    -- filter=5 channel=12
    -11, -12, 6, -7, -12, -18, -3, 5, -5,
    -- filter=5 channel=13
    13, 0, 7, 0, -2, -10, -13, 2, -13,
    -- filter=5 channel=14
    3, -2, 8, 1, -5, 1, 2, -1, 10,
    -- filter=5 channel=15
    -12, -8, -1, 2, -7, 14, -11, 4, 7,
    -- filter=5 channel=16
    13, 12, -7, 11, 7, -2, 4, 14, -2,
    -- filter=5 channel=17
    -14, -13, -1, -2, 4, 4, -19, -10, 7,
    -- filter=5 channel=18
    12, 8, 15, 20, 10, 7, 11, 18, 20,
    -- filter=5 channel=19
    0, 1, -9, -1, -9, -11, -10, -4, -4,
    -- filter=5 channel=20
    -13, -13, -4, 0, 11, 11, 8, 0, -14,
    -- filter=5 channel=21
    -12, 0, 5, -5, 6, -17, 10, -9, 0,
    -- filter=5 channel=22
    -10, -1, -16, -15, -12, -6, -9, 3, 0,
    -- filter=5 channel=23
    -6, 0, -1, 12, -11, -4, 14, 7, -1,
    -- filter=5 channel=24
    0, 7, 0, -2, 2, 8, 10, 15, -1,
    -- filter=5 channel=25
    18, -5, 15, 18, -3, 12, 9, 3, 10,
    -- filter=5 channel=26
    7, -3, -15, -2, 3, 8, -15, 11, 2,
    -- filter=5 channel=27
    13, 0, -7, 3, -9, -3, -11, 13, 7,
    -- filter=5 channel=28
    5, -8, 12, 2, -7, -10, -14, 10, 3,
    -- filter=5 channel=29
    -10, -1, -7, -5, -8, -2, -7, -15, 0,
    -- filter=5 channel=30
    4, -12, -2, 5, -2, -7, -2, 6, -10,
    -- filter=5 channel=31
    -1, 0, -14, -6, -11, -9, -7, 9, -15,
    -- filter=6 channel=0
    -19, -16, 1, -3, 2, -15, 8, -4, -19,
    -- filter=6 channel=1
    14, 2, 18, 0, 5, 16, -9, -3, -11,
    -- filter=6 channel=2
    -10, -7, 3, -14, 12, -8, -10, -3, -6,
    -- filter=6 channel=3
    -14, 0, 13, 3, -3, -1, -4, -7, -3,
    -- filter=6 channel=4
    0, 1, 20, 8, 0, 17, -17, 4, 1,
    -- filter=6 channel=5
    -9, -15, -10, -13, -16, 11, -8, 3, 1,
    -- filter=6 channel=6
    -6, -3, -2, 11, -2, 8, -5, 10, -5,
    -- filter=6 channel=7
    7, 18, -2, 5, 19, -2, -9, 5, 4,
    -- filter=6 channel=8
    -13, -1, -1, -8, 1, 9, 1, -16, -1,
    -- filter=6 channel=9
    13, 4, -12, -6, 7, -5, 5, -12, -10,
    -- filter=6 channel=10
    -20, -2, -8, 5, 7, -14, 5, -6, -15,
    -- filter=6 channel=11
    -7, -14, 4, -1, -10, -5, 13, 4, 5,
    -- filter=6 channel=12
    0, -11, -11, 12, 6, 11, 1, -6, 8,
    -- filter=6 channel=13
    -23, -2, -23, -4, -15, 5, -7, -13, -8,
    -- filter=6 channel=14
    10, -13, -5, 4, 1, 2, 5, 4, -3,
    -- filter=6 channel=15
    -14, 8, -6, -17, -1, 2, -14, -19, -10,
    -- filter=6 channel=16
    12, -2, -1, 4, 8, 11, 0, 3, 12,
    -- filter=6 channel=17
    3, 6, -1, -12, -12, 14, -18, -13, -7,
    -- filter=6 channel=18
    8, 1, 6, 5, 3, 2, 10, 9, 0,
    -- filter=6 channel=19
    -8, -8, -14, -4, -12, 9, -9, 4, -3,
    -- filter=6 channel=20
    13, 17, 16, 7, 12, 20, -8, 8, 18,
    -- filter=6 channel=21
    -10, 6, 15, -22, 0, -10, -13, -25, -18,
    -- filter=6 channel=22
    -11, -2, -6, -19, 5, 0, -3, -3, -1,
    -- filter=6 channel=23
    -13, -11, 6, 5, 6, -4, 4, -11, -11,
    -- filter=6 channel=24
    -8, 16, 9, 8, -11, 14, -7, 2, 1,
    -- filter=6 channel=25
    7, 11, 17, -20, -10, 2, -9, -9, -10,
    -- filter=6 channel=26
    -12, -16, -21, -5, -15, 0, 0, -11, -8,
    -- filter=6 channel=27
    0, -13, -13, 3, 12, -9, 12, 10, -7,
    -- filter=6 channel=28
    2, 11, 10, -6, -4, 8, -9, 14, 6,
    -- filter=6 channel=29
    -3, 7, 9, -5, -12, -11, -9, -8, -5,
    -- filter=6 channel=30
    12, 1, -14, 7, 8, -4, -9, -13, 10,
    -- filter=6 channel=31
    -11, -6, 4, 6, -9, 1, 2, -1, 2,
    -- filter=7 channel=0
    -8, 2, -13, -7, -12, -5, 0, 12, 5,
    -- filter=7 channel=1
    6, 6, -7, -10, 1, -3, 3, 6, -1,
    -- filter=7 channel=2
    -11, 11, -12, 10, 11, -8, 10, 0, 14,
    -- filter=7 channel=3
    14, 5, 1, -13, 7, -9, 2, 8, 4,
    -- filter=7 channel=4
    -10, 0, -8, -17, -1, 11, -19, -14, -13,
    -- filter=7 channel=5
    10, 16, 13, 7, -5, -4, -1, -9, -9,
    -- filter=7 channel=6
    2, 13, 2, 7, 7, 0, 12, -12, -9,
    -- filter=7 channel=7
    18, 6, 3, 8, 0, 11, 13, -11, -3,
    -- filter=7 channel=8
    8, 4, -15, 3, 0, -1, 15, 10, 0,
    -- filter=7 channel=9
    6, 12, 6, -10, 5, -1, 7, -10, 13,
    -- filter=7 channel=10
    5, 8, 12, -10, 11, -13, -14, -14, 0,
    -- filter=7 channel=11
    -20, -16, -5, -17, -7, 1, -9, 4, 0,
    -- filter=7 channel=12
    10, 0, -16, 6, 0, -13, -3, -3, -7,
    -- filter=7 channel=13
    13, 5, 9, 20, 18, -13, 14, 15, -10,
    -- filter=7 channel=14
    -8, -12, -2, -7, -13, -9, -3, -17, 10,
    -- filter=7 channel=15
    -5, 0, -11, -4, 10, 8, -10, -12, -15,
    -- filter=7 channel=16
    7, 1, 1, 4, 5, 4, -13, -14, 8,
    -- filter=7 channel=17
    9, 16, 5, 8, 17, 9, -10, 9, 3,
    -- filter=7 channel=18
    0, -3, 10, 1, 1, -5, 4, 12, -13,
    -- filter=7 channel=19
    -5, 8, 8, 0, 4, 10, 4, -8, 10,
    -- filter=7 channel=20
    0, 13, -3, -2, -4, 1, 5, 11, 3,
    -- filter=7 channel=21
    15, 12, 0, -4, -5, 10, -9, -9, 0,
    -- filter=7 channel=22
    -1, -4, 9, 16, 3, -4, 0, 2, 2,
    -- filter=7 channel=23
    0, -17, -4, -4, 1, 3, -6, -11, 0,
    -- filter=7 channel=24
    8, -17, -7, -16, -8, -8, 0, 6, -8,
    -- filter=7 channel=25
    -6, -5, 6, -15, -15, -16, -10, -13, -16,
    -- filter=7 channel=26
    16, -9, -13, 10, -4, -12, 16, -8, -8,
    -- filter=7 channel=27
    12, 7, -8, 12, -9, 1, 11, 14, 13,
    -- filter=7 channel=28
    -6, 2, 4, 5, -4, 6, -14, -13, 4,
    -- filter=7 channel=29
    -16, -6, -19, -14, 9, -14, -13, 8, -16,
    -- filter=7 channel=30
    6, -10, 3, -12, 7, -12, 3, -14, 7,
    -- filter=7 channel=31
    14, 17, -11, 13, 12, 12, 0, 7, -2,
    -- filter=8 channel=0
    1, -6, -13, -9, 4, 9, -4, 9, -4,
    -- filter=8 channel=1
    8, -1, 0, 7, 13, -4, -7, -4, -7,
    -- filter=8 channel=2
    6, 2, -8, -10, 0, 5, 0, -10, -6,
    -- filter=8 channel=3
    3, 4, -5, 1, -1, 14, 12, 5, -8,
    -- filter=8 channel=4
    15, 10, -7, 14, -12, -14, 0, 8, 0,
    -- filter=8 channel=5
    -3, 7, 12, 3, -9, -13, -12, 3, 2,
    -- filter=8 channel=6
    0, -8, 7, -12, 7, -6, 1, 13, 9,
    -- filter=8 channel=7
    -1, -11, -14, 10, 10, 9, -10, 10, 13,
    -- filter=8 channel=8
    3, 3, -1, 0, -1, -14, -14, -12, -7,
    -- filter=8 channel=9
    -7, 13, 12, 8, -13, 2, 1, 2, 13,
    -- filter=8 channel=10
    11, 8, -10, 8, 7, -2, 6, 0, -7,
    -- filter=8 channel=11
    -7, -2, 5, -9, 11, -1, -12, 4, -2,
    -- filter=8 channel=12
    -6, -6, 3, 0, 13, 12, -10, 9, -11,
    -- filter=8 channel=13
    -10, -9, -7, -6, 7, 3, -4, -7, 13,
    -- filter=8 channel=14
    12, 11, 8, 12, -13, 3, -10, -6, -4,
    -- filter=8 channel=15
    1, 3, 5, 8, 0, 13, 8, 12, 8,
    -- filter=8 channel=16
    0, -5, 8, -12, 10, 14, 12, -11, 14,
    -- filter=8 channel=17
    -11, 12, 2, -1, 9, 8, 1, -1, 1,
    -- filter=8 channel=18
    5, 4, 1, 3, -13, 13, -3, 5, 14,
    -- filter=8 channel=19
    -13, -13, 2, -1, -5, -6, -2, 11, 4,
    -- filter=8 channel=20
    -15, 9, -4, -13, -11, 7, -4, -9, 14,
    -- filter=8 channel=21
    7, 4, 1, 5, -10, -10, 12, -7, 1,
    -- filter=8 channel=22
    -15, 10, 0, 0, 4, 3, 17, 0, 11,
    -- filter=8 channel=23
    10, -13, 8, -8, 9, -8, 5, 13, 7,
    -- filter=8 channel=24
    1, 11, 5, 7, -6, -9, 14, 3, -2,
    -- filter=8 channel=25
    -10, -7, -5, -12, 6, -7, 5, -11, 12,
    -- filter=8 channel=26
    3, -15, 13, -9, 2, -1, -4, 6, 13,
    -- filter=8 channel=27
    -2, -14, -2, 11, -5, -10, 1, 4, -2,
    -- filter=8 channel=28
    8, 0, 10, 14, -12, 6, -9, 0, 6,
    -- filter=8 channel=29
    6, -6, -4, -7, -15, 11, 13, 10, 5,
    -- filter=8 channel=30
    3, 9, 14, -2, -5, 7, -6, -10, -2,
    -- filter=8 channel=31
    -15, -6, 8, 7, -7, -6, 4, -2, 4,
    -- filter=9 channel=0
    9, 0, -3, 6, 1, -11, -9, -6, 3,
    -- filter=9 channel=1
    -2, 11, 19, -14, -10, 9, -12, -15, 0,
    -- filter=9 channel=2
    11, 14, -9, 5, 8, 13, 6, 4, -14,
    -- filter=9 channel=3
    -8, 0, 11, 5, 9, 12, 7, 5, 0,
    -- filter=9 channel=4
    4, -1, 11, -2, -8, 7, 3, -9, 2,
    -- filter=9 channel=5
    3, -7, -5, 9, -4, 0, -3, 10, -5,
    -- filter=9 channel=6
    9, 2, -3, 7, -10, -5, -4, -11, 2,
    -- filter=9 channel=7
    0, 17, 2, 13, 12, -4, 3, -8, 11,
    -- filter=9 channel=8
    -3, -15, -5, 12, 5, 10, -8, 1, -4,
    -- filter=9 channel=9
    -5, 0, 4, 16, 5, 16, 4, -4, 0,
    -- filter=9 channel=10
    4, 8, -13, 1, -14, -8, 5, -6, -2,
    -- filter=9 channel=11
    -9, -14, -2, 10, -4, -10, 4, 5, -6,
    -- filter=9 channel=12
    12, 10, 4, 7, -4, 2, -11, 0, 9,
    -- filter=9 channel=13
    10, 0, 13, 15, 3, -8, -1, -18, 5,
    -- filter=9 channel=14
    -17, -20, -3, 3, -20, 5, -7, -11, 10,
    -- filter=9 channel=15
    14, 13, 5, 6, 2, 5, 5, 11, 3,
    -- filter=9 channel=16
    -12, -7, -11, 7, -5, 7, -13, 9, -8,
    -- filter=9 channel=17
    22, 17, 5, 12, -11, 6, 2, -2, -11,
    -- filter=9 channel=18
    -4, -5, -3, 5, -4, 7, -12, -2, 7,
    -- filter=9 channel=19
    2, 10, -12, 10, 13, -11, 10, -10, 11,
    -- filter=9 channel=20
    3, 0, 14, -14, 3, 17, -14, 6, 7,
    -- filter=9 channel=21
    1, -9, 17, 5, -2, 1, -12, -15, -11,
    -- filter=9 channel=22
    18, 1, 9, 20, 10, 3, 24, 10, 3,
    -- filter=9 channel=23
    -9, -17, 1, -8, 6, -12, 0, 5, 17,
    -- filter=9 channel=24
    -15, -7, -9, -13, 0, 9, 0, -1, -6,
    -- filter=9 channel=25
    -25, -10, -9, -19, -16, 12, -18, 9, 0,
    -- filter=9 channel=26
    -8, 13, 3, -4, -13, -16, 2, -8, -24,
    -- filter=9 channel=27
    -6, -7, 15, 4, 1, -8, 5, -6, -5,
    -- filter=9 channel=28
    1, 2, -4, 9, 12, 16, 0, -7, 2,
    -- filter=9 channel=29
    2, -5, 4, -13, -18, -4, -16, -12, -13,
    -- filter=9 channel=30
    -10, 4, -6, 14, -5, 5, 3, -10, 12,
    -- filter=9 channel=31
    23, 19, 13, 2, 9, -13, -9, -5, 10,
    -- filter=10 channel=0
    4, 17, 0, 16, 4, 2, -1, 19, 16,
    -- filter=10 channel=1
    -6, -4, -7, -14, -19, -14, -18, -18, -16,
    -- filter=10 channel=2
    -1, -5, 1, 5, -6, 5, 0, 10, 8,
    -- filter=10 channel=3
    8, -4, -1, -2, -9, 0, 14, -7, 14,
    -- filter=10 channel=4
    -14, -17, -18, 13, -11, 10, 6, 13, -11,
    -- filter=10 channel=5
    2, -8, -13, -14, 6, -13, 4, 5, -6,
    -- filter=10 channel=6
    14, 2, -1, -13, -14, -4, -2, -14, -10,
    -- filter=10 channel=7
    -4, -24, -16, -23, -2, -1, -2, 1, -11,
    -- filter=10 channel=8
    3, -8, 16, 14, -3, 19, 6, 2, 8,
    -- filter=10 channel=9
    -5, -9, -4, 3, 0, -13, -10, -7, -7,
    -- filter=10 channel=10
    7, 11, 6, 2, -7, 9, -6, 0, 11,
    -- filter=10 channel=11
    20, 21, 2, 0, 10, 4, -9, -7, 17,
    -- filter=10 channel=12
    -5, 11, -5, 2, -5, -12, 12, -14, -9,
    -- filter=10 channel=13
    -7, 11, -4, -5, 4, -2, 15, -12, 2,
    -- filter=10 channel=14
    -13, 5, -3, -5, -4, 11, -15, 6, 3,
    -- filter=10 channel=15
    15, -12, 9, -12, 4, -2, -13, 5, -14,
    -- filter=10 channel=16
    -16, 6, -6, -3, -7, -14, -13, -10, -6,
    -- filter=10 channel=17
    4, 3, -21, 0, -2, -15, -4, 6, -1,
    -- filter=10 channel=18
    -5, -11, 11, 2, 5, -2, 2, -3, 9,
    -- filter=10 channel=19
    7, -9, -9, -13, -9, 9, 6, -11, -7,
    -- filter=10 channel=20
    -12, -27, -16, -3, -23, -20, -23, -9, -26,
    -- filter=10 channel=21
    -16, -11, -4, -4, -3, -15, 0, 2, -17,
    -- filter=10 channel=22
    -2, 24, 1, 8, 0, 14, 4, 17, 2,
    -- filter=10 channel=23
    17, 8, 16, 12, 2, -10, 5, 0, 13,
    -- filter=10 channel=24
    9, 2, 8, 10, 0, -5, -12, -11, 10,
    -- filter=10 channel=25
    13, 3, 5, 21, 18, 16, 8, 12, 2,
    -- filter=10 channel=26
    9, -11, -13, 12, -7, 14, 8, 2, -5,
    -- filter=10 channel=27
    0, 12, 12, 5, 3, -1, 7, -10, 1,
    -- filter=10 channel=28
    4, -13, -9, -3, -14, 11, -9, 2, 7,
    -- filter=10 channel=29
    8, 14, 14, -2, 0, -6, 16, -8, -3,
    -- filter=10 channel=30
    -6, -14, -3, -4, -6, 11, 13, -14, -13,
    -- filter=10 channel=31
    -9, 11, -11, -10, -4, -15, 11, -6, 5,
    -- filter=11 channel=0
    -8, 11, 7, -11, -14, 4, -13, 5, 0,
    -- filter=11 channel=1
    -8, 12, 10, -5, 8, -10, -7, 0, 4,
    -- filter=11 channel=2
    -12, 6, 10, -7, 14, 7, -4, 9, 4,
    -- filter=11 channel=3
    -1, 4, 12, -13, -8, 0, 0, -13, 3,
    -- filter=11 channel=4
    -12, -10, -9, -3, -16, 12, 8, 12, 7,
    -- filter=11 channel=5
    15, 9, -15, 0, 11, -3, 4, -5, -14,
    -- filter=11 channel=6
    -10, -10, 11, 4, 13, 0, 9, 9, -10,
    -- filter=11 channel=7
    14, 2, 0, 16, 2, -8, 12, -2, 8,
    -- filter=11 channel=8
    12, -9, -14, 8, -5, -2, 3, 6, -7,
    -- filter=11 channel=9
    -10, -4, -6, -7, -8, -4, 9, 5, -8,
    -- filter=11 channel=10
    -14, -9, -4, -15, 9, 9, -8, -12, -2,
    -- filter=11 channel=11
    1, 3, -1, 10, -2, 12, 3, 13, -3,
    -- filter=11 channel=12
    -5, -19, 0, 5, -18, 9, 14, -2, 5,
    -- filter=11 channel=13
    16, -4, -9, 10, -6, 13, 7, 5, -10,
    -- filter=11 channel=14
    5, 1, 11, -1, 3, 0, -14, 12, -9,
    -- filter=11 channel=15
    5, -16, -7, 15, 5, -8, -6, 1, 1,
    -- filter=11 channel=16
    7, -7, 11, -2, 8, 0, 3, -6, 1,
    -- filter=11 channel=17
    -2, -15, -3, 14, -1, 8, 15, 7, 9,
    -- filter=11 channel=18
    1, 9, 0, 8, 0, 10, 4, -11, 3,
    -- filter=11 channel=19
    0, -1, 0, -1, -11, -8, -9, 2, 4,
    -- filter=11 channel=20
    6, -14, -16, 17, 2, -6, 22, 16, -3,
    -- filter=11 channel=21
    5, 9, -15, -7, -14, 2, -2, -2, -2,
    -- filter=11 channel=22
    -14, -5, -2, -12, -18, 0, 8, 10, -13,
    -- filter=11 channel=23
    4, -2, -13, 6, 5, -7, 0, -5, 10,
    -- filter=11 channel=24
    -12, 0, 6, -11, -2, 13, 12, 14, 11,
    -- filter=11 channel=25
    -3, -9, -20, -1, -12, -7, 1, -17, -15,
    -- filter=11 channel=26
    0, 10, -14, 8, 0, -12, -2, -16, 4,
    -- filter=11 channel=27
    -8, 8, 12, -9, 3, 3, 0, -7, 3,
    -- filter=11 channel=28
    6, 10, 6, 3, 4, 9, -1, 10, -5,
    -- filter=11 channel=29
    -1, 12, 6, -11, 13, 15, 12, 0, -2,
    -- filter=11 channel=30
    3, 3, -14, -3, 8, 4, -7, 11, 9,
    -- filter=11 channel=31
    -7, -2, 2, -11, 0, -7, 8, 10, 10,
    -- filter=12 channel=0
    -5, -9, 12, 0, 10, 6, -12, -6, -10,
    -- filter=12 channel=1
    0, 8, 7, -4, -9, 8, 0, -7, -1,
    -- filter=12 channel=2
    -4, 3, 4, -13, -14, 1, 8, -9, 7,
    -- filter=12 channel=3
    -6, 10, 10, 6, 13, 5, 11, 8, -4,
    -- filter=12 channel=4
    -4, -8, 15, -5, 12, 6, 3, -6, 11,
    -- filter=12 channel=5
    3, 0, 6, 8, -7, -9, -4, -8, -6,
    -- filter=12 channel=6
    -4, 0, 0, 3, -5, -7, 10, 6, -13,
    -- filter=12 channel=7
    17, 16, -12, 0, 4, -17, -5, -8, -5,
    -- filter=12 channel=8
    -1, 5, 4, 1, -6, 0, 10, -7, -13,
    -- filter=12 channel=9
    -14, 7, 7, 8, -13, 4, 7, -8, 7,
    -- filter=12 channel=10
    -3, -7, 0, 9, -2, -12, 2, 0, 4,
    -- filter=12 channel=11
    13, 13, -16, 5, 0, -14, -2, -4, 13,
    -- filter=12 channel=12
    -4, 4, 8, -10, 2, -11, 2, 8, -2,
    -- filter=12 channel=13
    13, -10, -3, 14, 8, -13, 12, -2, -12,
    -- filter=12 channel=14
    -3, 6, 9, -5, 4, 17, -13, 14, 6,
    -- filter=12 channel=15
    0, 0, -11, 7, -4, 6, 16, 9, -1,
    -- filter=12 channel=16
    11, 0, 8, 12, 12, -13, 12, 9, 5,
    -- filter=12 channel=17
    24, 11, -12, 0, -10, 2, 12, -9, -24,
    -- filter=12 channel=18
    1, 10, -2, -5, 4, 1, -8, 2, -6,
    -- filter=12 channel=19
    -7, 7, 6, -2, 13, -10, -9, 3, 7,
    -- filter=12 channel=20
    9, 3, 18, 18, -6, 12, 3, 14, -11,
    -- filter=12 channel=21
    14, 5, -8, 7, 0, -8, 2, -13, -2,
    -- filter=12 channel=22
    -3, -8, -3, -14, -1, -18, -16, 1, -10,
    -- filter=12 channel=23
    -15, -11, 2, -1, -1, 1, -13, -10, -3,
    -- filter=12 channel=24
    8, -3, 10, 13, 12, 19, -12, 0, -3,
    -- filter=12 channel=25
    -11, 2, 12, -2, -3, -2, -18, -8, -13,
    -- filter=12 channel=26
    2, -14, -15, 18, 8, 7, 21, -13, -7,
    -- filter=12 channel=27
    -6, -15, -7, -9, -2, -1, -13, -10, 0,
    -- filter=12 channel=28
    -6, 14, 1, 3, 11, -6, -7, -7, 0,
    -- filter=12 channel=29
    8, -10, 9, -9, 5, 6, 6, -9, 5,
    -- filter=12 channel=30
    -4, -10, 7, 6, 1, -9, 0, -11, -7,
    -- filter=12 channel=31
    16, 11, -2, 14, 1, -2, -6, 9, -11,
    -- filter=13 channel=0
    6, -3, -9, -1, -13, 1, -7, 2, 14,
    -- filter=13 channel=1
    6, 3, 12, 4, -13, 13, -5, 6, -6,
    -- filter=13 channel=2
    7, 14, 5, -4, -3, -8, -12, -7, -3,
    -- filter=13 channel=3
    14, -5, 11, -2, 11, 12, -3, -9, 13,
    -- filter=13 channel=4
    -9, -13, 5, 6, -2, 9, -5, -6, -8,
    -- filter=13 channel=5
    0, -5, 10, 9, -4, 10, -5, 10, 10,
    -- filter=13 channel=6
    -12, -4, 8, 6, 8, 10, -10, -10, 9,
    -- filter=13 channel=7
    -16, 8, 10, 11, 13, 8, 8, 0, 6,
    -- filter=13 channel=8
    -8, 9, 0, 12, 0, -9, 13, -6, -4,
    -- filter=13 channel=9
    -7, -9, -3, 0, -7, -16, -1, -5, -15,
    -- filter=13 channel=10
    11, 11, 8, 9, 9, -7, 9, 2, 14,
    -- filter=13 channel=11
    5, -9, 5, -5, -7, -7, 9, -10, 18,
    -- filter=13 channel=12
    5, 10, 5, -5, -2, -10, -3, -13, 11,
    -- filter=13 channel=13
    -6, 9, -2, 6, 9, 2, 0, 10, 19,
    -- filter=13 channel=14
    -14, -11, 4, -14, -10, 1, -16, -11, 5,
    -- filter=13 channel=15
    3, 13, -5, -2, 5, 11, 15, 7, -11,
    -- filter=13 channel=16
    13, 1, 0, -10, -9, 5, -14, -3, 15,
    -- filter=13 channel=17
    -7, -3, 8, 15, 11, -11, -7, 16, 2,
    -- filter=13 channel=18
    -1, -12, -12, -15, -5, -4, 0, -14, -16,
    -- filter=13 channel=19
    12, 2, -3, 0, -9, -12, 8, -9, 6,
    -- filter=13 channel=20
    -9, -2, 7, 1, 1, 12, -5, 5, -9,
    -- filter=13 channel=21
    -12, -10, 4, -12, 8, -5, 10, 3, -10,
    -- filter=13 channel=22
    -11, -20, -8, -7, -5, -1, -9, 5, 2,
    -- filter=13 channel=23
    -17, -14, -7, 2, -17, -9, 11, -6, -9,
    -- filter=13 channel=24
    1, -11, -9, -2, 1, 10, -2, -7, 0,
    -- filter=13 channel=25
    -15, -8, -6, -8, -21, -16, 0, -18, -20,
    -- filter=13 channel=26
    8, 0, 0, 20, 8, 5, 20, 12, 12,
    -- filter=13 channel=27
    1, 7, -3, -12, 9, 3, 4, -3, -5,
    -- filter=13 channel=28
    -5, 5, -10, 8, 1, -10, 11, -7, -7,
    -- filter=13 channel=29
    -11, 11, -4, 15, 7, -4, 13, 9, -5,
    -- filter=13 channel=30
    0, -14, -7, 10, -13, -12, 0, -8, -5,
    -- filter=13 channel=31
    16, -1, 12, -4, -4, 0, 13, 5, -14,
    -- filter=14 channel=0
    -8, 10, -15, 3, 11, -10, 13, -12, -3,
    -- filter=14 channel=1
    11, 2, 19, 9, 5, 11, -13, 14, -5,
    -- filter=14 channel=2
    1, 9, -12, -5, -12, 4, -5, 7, 14,
    -- filter=14 channel=3
    7, 0, 0, 4, -14, 6, 2, -8, -6,
    -- filter=14 channel=4
    8, 7, 17, -1, 11, 18, -1, 7, 8,
    -- filter=14 channel=5
    -4, -1, -15, -11, 6, -12, -7, -8, -15,
    -- filter=14 channel=6
    -7, 10, 1, 4, 11, -13, 11, -12, -12,
    -- filter=14 channel=7
    -12, -10, 14, 6, -2, -5, -13, 0, 10,
    -- filter=14 channel=8
    11, 12, 6, -10, 9, -9, -2, -9, -13,
    -- filter=14 channel=9
    14, -6, 0, -1, -1, 11, 13, 6, -5,
    -- filter=14 channel=10
    12, -2, 1, 2, 0, -9, -9, 12, -11,
    -- filter=14 channel=11
    -16, -4, -4, -14, -2, -15, 10, -16, -17,
    -- filter=14 channel=12
    -12, 3, -13, -9, -14, 6, 4, 10, -1,
    -- filter=14 channel=13
    4, 13, 10, 15, 14, 5, 15, -3, 1,
    -- filter=14 channel=14
    -16, -14, -13, 0, 12, -4, -5, 11, 10,
    -- filter=14 channel=15
    11, -14, -11, 8, -14, 7, 1, -9, -6,
    -- filter=14 channel=16
    -10, -7, 15, -9, -1, -2, -7, 0, -4,
    -- filter=14 channel=17
    3, -12, 12, 3, 10, 12, 13, -9, 6,
    -- filter=14 channel=18
    -2, 10, -6, 1, -1, 0, -7, -11, 14,
    -- filter=14 channel=19
    -1, 6, -14, 0, 5, 14, 9, -4, -1,
    -- filter=14 channel=20
    8, -5, 1, -1, -5, 17, -2, -19, -7,
    -- filter=14 channel=21
    9, 11, 3, 12, -1, 13, -1, -5, -9,
    -- filter=14 channel=22
    -2, -20, -2, 0, -7, -9, -8, -7, -17,
    -- filter=14 channel=23
    -13, 7, -14, 2, 10, 5, -3, -6, 4,
    -- filter=14 channel=24
    4, -16, 7, -6, -5, 15, 7, 7, -13,
    -- filter=14 channel=25
    -15, 8, 13, -12, 8, 4, -1, 1, -5,
    -- filter=14 channel=26
    15, -3, -15, 3, 3, -4, 17, 10, 0,
    -- filter=14 channel=27
    0, -6, -5, 14, -12, -1, 1, 7, -7,
    -- filter=14 channel=28
    9, 13, 7, 12, -6, -8, -7, -15, 5,
    -- filter=14 channel=29
    -13, -5, 4, -10, -7, 5, -2, -13, -14,
    -- filter=14 channel=30
    6, 2, 8, 0, 3, -1, -10, -7, -11,
    -- filter=14 channel=31
    -3, 1, -11, 4, -5, 4, -2, -8, 9,
    -- filter=15 channel=0
    17, 14, -9, 13, -3, 0, 8, -1, 5,
    -- filter=15 channel=1
    -5, 4, -8, -12, -6, -4, 1, -5, 9,
    -- filter=15 channel=2
    8, -6, -10, 7, -6, 11, -14, -8, -3,
    -- filter=15 channel=3
    4, 5, -3, 10, 12, 5, -13, 6, -13,
    -- filter=15 channel=4
    -8, -18, 12, 1, -11, 10, -20, -10, 0,
    -- filter=15 channel=5
    -16, -6, -9, 7, 4, -15, 3, 5, -10,
    -- filter=15 channel=6
    10, 0, -9, -4, 4, 1, -7, -1, 5,
    -- filter=15 channel=7
    -6, 0, 7, -16, 0, 0, 4, -3, 6,
    -- filter=15 channel=8
    7, 0, -11, -10, -1, -12, -8, -8, 2,
    -- filter=15 channel=9
    -10, 12, 9, 6, 7, -7, -6, 11, 9,
    -- filter=15 channel=10
    -9, 6, 0, 11, -5, 3, 4, -8, 12,
    -- filter=15 channel=11
    -6, 18, 13, 11, -5, 13, 19, 0, 3,
    -- filter=15 channel=12
    -13, -12, 4, 9, -3, 17, -3, -7, -8,
    -- filter=15 channel=13
    23, 16, 25, 23, 25, 27, 18, 2, 10,
    -- filter=15 channel=14
    12, 4, 1, -12, 6, 1, 0, -14, -9,
    -- filter=15 channel=15
    10, -3, 2, -11, 1, 6, 5, -11, 11,
    -- filter=15 channel=16
    7, -3, 10, -12, -8, -12, 5, -9, 2,
    -- filter=15 channel=17
    4, 0, -1, -14, 4, 16, -4, -6, 5,
    -- filter=15 channel=18
    -12, -2, 8, -3, -6, 10, -9, 3, -13,
    -- filter=15 channel=19
    -14, 14, -12, -9, -12, 8, -1, -6, 5,
    -- filter=15 channel=20
    -24, 7, 12, -21, -12, 11, 0, 1, 4,
    -- filter=15 channel=21
    -20, -16, 9, -13, -12, -7, 2, -21, -3,
    -- filter=15 channel=22
    0, -15, -14, -14, -3, -7, -8, 8, 3,
    -- filter=15 channel=23
    -17, -3, -13, 7, -7, -1, 0, -3, 0,
    -- filter=15 channel=24
    -7, -10, -3, 7, 2, -2, -17, -4, -10,
    -- filter=15 channel=25
    -16, 4, -5, 3, 1, -11, -15, -18, -19,
    -- filter=15 channel=26
    12, 2, 12, 8, -1, -1, -2, 7, 1,
    -- filter=15 channel=27
    -12, -10, -13, 0, 10, 13, -6, -1, 0,
    -- filter=15 channel=28
    9, -4, -3, 8, -17, -11, -6, -11, 7,
    -- filter=15 channel=29
    6, -12, -6, -8, -3, -11, 16, 15, -11,
    -- filter=15 channel=30
    -1, -8, 12, 1, 11, 14, 3, -8, 6,
    -- filter=15 channel=31
    -8, -8, 3, -5, -2, 7, 3, -15, -4,
    -- filter=16 channel=0
    -16, 0, -1, -14, -6, 13, -15, -14, 2,
    -- filter=16 channel=1
    -8, -5, -4, 12, -13, 7, 8, 2, 11,
    -- filter=16 channel=2
    14, -8, 12, 12, -1, 2, 2, 13, -5,
    -- filter=16 channel=3
    10, -8, -9, -7, 8, 1, 13, 11, -7,
    -- filter=16 channel=4
    -5, -12, 1, 1, -8, 3, 7, -9, 4,
    -- filter=16 channel=5
    -7, -3, -10, -1, -9, -1, 2, 7, -1,
    -- filter=16 channel=6
    11, 1, 0, -9, 0, -3, 0, -9, 5,
    -- filter=16 channel=7
    7, -16, -3, 1, 12, -14, -13, -16, 6,
    -- filter=16 channel=8
    -9, -2, -5, 7, 1, -4, 10, 6, -7,
    -- filter=16 channel=9
    0, 2, -13, -3, -5, 1, 0, -5, -12,
    -- filter=16 channel=10
    1, 9, -12, 0, 9, -9, 13, 3, 8,
    -- filter=16 channel=11
    2, 5, 12, -15, 10, -4, 12, -10, -9,
    -- filter=16 channel=12
    12, -2, 12, 1, -12, 1, -11, 4, 7,
    -- filter=16 channel=13
    0, -13, -7, 3, -12, 4, 11, 11, 3,
    -- filter=16 channel=14
    -8, 0, -9, -14, -10, 8, 1, 10, 12,
    -- filter=16 channel=15
    -7, 3, -4, -3, 4, 0, 7, -8, 2,
    -- filter=16 channel=16
    -6, -2, -5, -9, 3, 1, -13, 0, -3,
    -- filter=16 channel=17
    11, 5, 6, 9, 12, -11, 15, 1, 1,
    -- filter=16 channel=18
    11, -8, 11, -1, -10, -11, -1, 0, -3,
    -- filter=16 channel=19
    -5, -12, -6, 10, 1, -12, 9, -3, -12,
    -- filter=16 channel=20
    5, 0, 5, 0, -4, 9, 5, -2, -5,
    -- filter=16 channel=21
    9, 11, 11, 2, 8, 10, 5, 4, 7,
    -- filter=16 channel=22
    -4, -16, -21, 6, -11, -13, -13, -10, -6,
    -- filter=16 channel=23
    5, 1, 3, 11, 13, 2, -11, 6, -1,
    -- filter=16 channel=24
    4, 10, 7, 7, -11, 10, -11, -8, -5,
    -- filter=16 channel=25
    -13, 0, -11, -1, 0, 9, -15, 0, -13,
    -- filter=16 channel=26
    16, 6, -12, 16, -1, -3, 10, 12, -5,
    -- filter=16 channel=27
    -11, -3, -2, 11, 0, 4, -10, 1, -5,
    -- filter=16 channel=28
    2, -8, -8, -2, 5, -3, 1, -5, -15,
    -- filter=16 channel=29
    8, -5, 12, -7, -4, 0, -1, 13, 7,
    -- filter=16 channel=30
    13, 6, -1, -6, 1, -6, 9, -13, 12,
    -- filter=16 channel=31
    -2, -7, -16, 10, -14, -18, 1, 9, 1,
    -- filter=17 channel=0
    -14, -4, -11, 14, 2, 12, -2, -13, 5,
    -- filter=17 channel=1
    -8, 9, -5, 2, -4, 5, 1, 8, 4,
    -- filter=17 channel=2
    7, -13, 0, -11, -11, -8, -8, 13, 10,
    -- filter=17 channel=3
    0, 12, 10, 0, 13, -10, -12, 14, -11,
    -- filter=17 channel=4
    8, -7, 11, -3, -14, -12, -10, -6, 0,
    -- filter=17 channel=5
    -10, -8, 2, 5, 14, 14, 13, -7, 13,
    -- filter=17 channel=6
    -2, 12, 13, -10, 1, 3, -14, -10, -5,
    -- filter=17 channel=7
    -12, -4, 10, 12, 12, -11, 12, -1, 1,
    -- filter=17 channel=8
    10, -1, 1, -1, 8, -4, 2, 0, 0,
    -- filter=17 channel=9
    13, 3, 7, -7, -1, 8, -7, 4, -13,
    -- filter=17 channel=10
    0, 9, -12, -8, 9, -9, -12, -9, 1,
    -- filter=17 channel=11
    14, -5, 3, -2, 9, 1, 10, -8, -8,
    -- filter=17 channel=12
    4, 0, -10, -10, 7, -4, -3, 0, 9,
    -- filter=17 channel=13
    7, 14, -7, -12, 12, -8, 1, -14, 2,
    -- filter=17 channel=14
    -11, 8, 7, -6, 10, -1, 2, 0, -11,
    -- filter=17 channel=15
    -3, 12, -7, 6, -12, 5, -10, -9, -6,
    -- filter=17 channel=16
    -7, -10, -8, -10, -6, 3, 2, -11, -9,
    -- filter=17 channel=17
    8, 5, -14, 6, -11, -1, -13, -1, 1,
    -- filter=17 channel=18
    5, -7, -13, 12, 8, 0, -1, 14, -10,
    -- filter=17 channel=19
    -14, 2, 10, -14, -10, -6, -13, -2, -13,
    -- filter=17 channel=20
    2, -11, 7, 8, -8, -1, -8, -3, 8,
    -- filter=17 channel=21
    -8, -6, -13, 14, 13, 9, -5, 0, -5,
    -- filter=17 channel=22
    5, 8, 11, 0, -3, 9, 9, 8, -13,
    -- filter=17 channel=23
    14, -13, -13, 11, -5, 8, 0, -5, 11,
    -- filter=17 channel=24
    -3, -9, 9, 12, -1, -2, 7, 1, -14,
    -- filter=17 channel=25
    11, 1, -3, 5, -4, -11, 0, -10, 1,
    -- filter=17 channel=26
    10, 0, 1, 9, -14, 9, -6, -10, -9,
    -- filter=17 channel=27
    5, -1, 6, -9, -2, 0, 7, -1, -11,
    -- filter=17 channel=28
    14, 8, -1, -8, -1, -9, 11, -7, 0,
    -- filter=17 channel=29
    0, -9, -6, -11, -8, 0, 0, 5, -1,
    -- filter=17 channel=30
    2, 4, 1, 0, -6, 0, -14, 1, -15,
    -- filter=17 channel=31
    -12, 0, -5, 6, -11, -10, -10, -13, -14,
    -- filter=18 channel=0
    -11, 2, -8, 3, 10, -4, 0, 8, 15,
    -- filter=18 channel=1
    1, -3, -6, -12, -3, 3, 4, -16, -12,
    -- filter=18 channel=2
    9, -14, 14, -11, 6, 0, 14, 5, -14,
    -- filter=18 channel=3
    5, 2, -2, 6, -6, 14, -11, -6, -2,
    -- filter=18 channel=4
    3, -14, -2, -3, -8, 13, 9, 3, 10,
    -- filter=18 channel=5
    -8, -14, -8, 8, -5, 14, -1, 13, -12,
    -- filter=18 channel=6
    -8, -7, -8, 11, 10, 12, -4, 14, -13,
    -- filter=18 channel=7
    3, -2, -14, -18, 5, 0, -11, 3, 7,
    -- filter=18 channel=8
    1, -1, 2, -10, 2, -8, -4, -1, 4,
    -- filter=18 channel=9
    -12, -7, 0, 12, -6, -3, -1, -6, 12,
    -- filter=18 channel=10
    1, -2, 9, -4, 8, 0, -6, 6, 7,
    -- filter=18 channel=11
    -6, 10, 4, 0, -6, -3, 5, 3, 1,
    -- filter=18 channel=12
    -11, -3, 7, 13, -5, 9, -8, 1, 5,
    -- filter=18 channel=13
    14, 12, -3, -9, 8, 17, 13, 0, 9,
    -- filter=18 channel=14
    12, -5, 10, 12, -5, 4, -13, -14, -8,
    -- filter=18 channel=15
    2, -1, 0, -1, -6, 8, 2, -6, 1,
    -- filter=18 channel=16
    12, -9, 8, -9, -5, -2, 4, 7, -10,
    -- filter=18 channel=17
    -1, -16, 7, -1, -10, 5, 9, 0, 13,
    -- filter=18 channel=18
    -2, -2, -1, 11, 3, 8, 9, -13, 10,
    -- filter=18 channel=19
    -9, -13, 9, -1, 14, 13, -1, 5, 10,
    -- filter=18 channel=20
    -15, -14, 0, -12, -4, -5, 4, -16, -17,
    -- filter=18 channel=21
    -15, -12, -11, 2, 8, -15, 9, 3, 8,
    -- filter=18 channel=22
    6, 10, -3, -3, 5, -4, 6, 12, -14,
    -- filter=18 channel=23
    5, -9, 2, 2, 4, 11, 10, 10, -12,
    -- filter=18 channel=24
    -10, -7, -1, -11, -13, 0, -11, -11, -5,
    -- filter=18 channel=25
    -5, -5, -6, 2, -14, -10, -4, -4, 10,
    -- filter=18 channel=26
    -3, 2, -7, 13, -3, 8, 7, 13, -4,
    -- filter=18 channel=27
    11, -2, 4, 7, 4, 1, 2, 9, -1,
    -- filter=18 channel=28
    -5, 4, -10, 13, -4, 4, -3, 7, -9,
    -- filter=18 channel=29
    -11, -6, -15, -7, 1, -16, 14, -6, -11,
    -- filter=18 channel=30
    4, 6, 12, 9, -10, -10, -7, -6, 5,
    -- filter=18 channel=31
    9, 7, -6, 9, 9, 9, -8, 5, 12,
    -- filter=19 channel=0
    -8, -2, 6, 14, -10, 17, 0, 5, -6,
    -- filter=19 channel=1
    -6, 6, 10, 9, -9, 6, 4, -2, 14,
    -- filter=19 channel=2
    1, 8, 1, 10, 5, 7, 10, -10, 9,
    -- filter=19 channel=3
    -13, -13, 7, -14, 7, 15, -12, 4, 1,
    -- filter=19 channel=4
    2, 6, 15, 5, -7, 5, -2, 3, 12,
    -- filter=19 channel=5
    -13, -13, 8, -1, 14, -2, -11, 0, 11,
    -- filter=19 channel=6
    -11, -12, 5, -11, -11, -7, 3, -1, 14,
    -- filter=19 channel=7
    -14, -2, -6, 3, 15, -6, -1, -11, 2,
    -- filter=19 channel=8
    7, -2, 11, 7, 2, -6, -7, 0, 2,
    -- filter=19 channel=9
    6, 5, 14, 13, -8, -4, -4, 0, -4,
    -- filter=19 channel=10
    13, 2, 3, 10, 0, -7, -12, 1, 0,
    -- filter=19 channel=11
    -15, -16, 1, -15, -17, 4, -11, 4, -12,
    -- filter=19 channel=12
    16, -5, 8, -7, 3, 14, 0, -2, 0,
    -- filter=19 channel=13
    8, 3, -3, -5, -12, -6, 7, -8, 8,
    -- filter=19 channel=14
    14, 11, 8, 5, 5, 1, -6, 5, 1,
    -- filter=19 channel=15
    11, 8, -3, 13, 8, -10, 9, -9, 1,
    -- filter=19 channel=16
    -18, -9, 1, 0, 12, -7, -17, -17, 7,
    -- filter=19 channel=17
    13, -7, 11, 11, 0, 5, -17, -18, 1,
    -- filter=19 channel=18
    11, 1, 6, 0, 5, 11, 10, 10, -5,
    -- filter=19 channel=19
    3, -1, 10, -10, 4, 12, 2, 0, -13,
    -- filter=19 channel=20
    10, -16, 0, -19, -17, 14, -22, -7, 4,
    -- filter=19 channel=21
    -3, 10, 17, 1, 2, 17, -8, 0, -11,
    -- filter=19 channel=22
    -6, 12, 14, -1, 3, 0, 11, 11, 16,
    -- filter=19 channel=23
    9, 10, -7, -11, 1, -2, -2, 0, -7,
    -- filter=19 channel=24
    -12, 11, 0, 5, -12, 10, -16, -9, 0,
    -- filter=19 channel=25
    11, 20, 21, -6, -4, 13, 5, 3, 0,
    -- filter=19 channel=26
    -10, 9, 1, -11, 5, 10, -14, 14, -4,
    -- filter=19 channel=27
    10, 11, -9, 8, 6, 2, 0, -9, 13,
    -- filter=19 channel=28
    -5, 14, 9, 9, 7, 8, -8, -1, -13,
    -- filter=19 channel=29
    3, -13, -18, 11, -12, -18, -4, -15, -10,
    -- filter=19 channel=30
    -2, -6, 11, 4, 15, -9, -15, 0, -8,
    -- filter=19 channel=31
    -2, 8, 10, 0, 1, 16, 10, 7, -13,
    -- filter=20 channel=0
    -4, -7, 9, 10, 17, 0, 3, 0, 3,
    -- filter=20 channel=1
    -2, -6, -24, 7, -20, -7, -3, -6, -13,
    -- filter=20 channel=2
    -11, 7, 11, -5, -11, 0, 3, 0, 14,
    -- filter=20 channel=3
    0, 8, 6, -6, -13, 8, -4, 6, -10,
    -- filter=20 channel=4
    12, 0, 8, 6, -7, 0, 10, 14, -11,
    -- filter=20 channel=5
    6, -2, 12, 5, 6, -10, -7, 11, -3,
    -- filter=20 channel=6
    -10, -11, 7, 1, 4, 11, 6, -8, -9,
    -- filter=20 channel=7
    8, -7, -6, 10, -4, -3, 6, -16, -34,
    -- filter=20 channel=8
    -10, 11, -13, 2, -10, -9, -1, 7, -1,
    -- filter=20 channel=9
    0, 12, 16, 10, 2, 19, 0, 13, 16,
    -- filter=20 channel=10
    -6, 8, 10, 0, 20, 10, 4, -1, 16,
    -- filter=20 channel=11
    6, -13, 3, -15, 6, 6, 0, 9, 4,
    -- filter=20 channel=12
    18, 19, 19, 13, 1, -8, 13, 8, -1,
    -- filter=20 channel=13
    7, -2, -14, 14, -6, -8, 5, -19, 2,
    -- filter=20 channel=14
    -10, -8, 0, -19, -14, 4, -12, 4, -17,
    -- filter=20 channel=15
    19, -2, -1, 13, -7, 7, 8, 2, -8,
    -- filter=20 channel=16
    -16, -4, 0, -4, 7, -17, -10, -13, -4,
    -- filter=20 channel=17
    25, -11, -13, -2, -9, -27, -6, -20, -11,
    -- filter=20 channel=18
    -5, 3, 4, 13, 12, -5, -3, 4, 1,
    -- filter=20 channel=19
    -7, -7, -10, -4, 0, -6, 3, -12, -10,
    -- filter=20 channel=20
    25, 6, -3, 10, -23, -12, 0, -30, -34,
    -- filter=20 channel=21
    23, 19, 7, 21, -13, -27, 0, -20, -6,
    -- filter=20 channel=22
    27, 45, 30, 37, 42, 30, 14, 16, 31,
    -- filter=20 channel=23
    15, -1, 9, 4, 8, 16, 17, 6, 18,
    -- filter=20 channel=24
    2, -14, 1, -8, -19, -25, -9, -24, -16,
    -- filter=20 channel=25
    29, 23, -1, 28, -1, 3, 24, 15, 0,
    -- filter=20 channel=26
    4, 14, 5, 15, 17, -11, 24, 4, -10,
    -- filter=20 channel=27
    -12, 11, -4, -12, 8, -14, -13, 6, 7,
    -- filter=20 channel=28
    10, -10, 2, 3, -10, 0, 17, -11, -8,
    -- filter=20 channel=29
    -3, -15, 3, -17, -17, -3, -20, 6, -3,
    -- filter=20 channel=30
    10, -9, 2, 4, -4, 0, 8, 4, -11,
    -- filter=20 channel=31
    20, -2, -7, 5, -5, -18, 15, -12, 1,
    -- filter=21 channel=0
    1, -10, 11, 11, -13, 6, -6, 12, 9,
    -- filter=21 channel=1
    -13, -5, -2, 0, 7, 6, -14, -4, -12,
    -- filter=21 channel=2
    3, -9, 14, 1, 5, 6, -7, -14, -10,
    -- filter=21 channel=3
    3, -6, 3, 0, 3, -1, 7, 13, 11,
    -- filter=21 channel=4
    -3, 5, -2, -4, 1, 10, -2, -9, -2,
    -- filter=21 channel=5
    0, 8, 12, -12, 0, -14, 6, 0, -4,
    -- filter=21 channel=6
    4, -5, 0, 2, 1, 4, -3, 13, -2,
    -- filter=21 channel=7
    6, 11, -3, -9, -3, -5, 9, -10, -11,
    -- filter=21 channel=8
    4, 14, -2, -14, -6, 11, 10, -11, -5,
    -- filter=21 channel=9
    10, -8, 15, 14, 12, 4, -1, 7, -7,
    -- filter=21 channel=10
    0, 13, 0, -9, 0, 4, -10, -2, 4,
    -- filter=21 channel=11
    -13, -13, 4, 0, 10, 13, -9, 6, 14,
    -- filter=21 channel=12
    -12, -1, -13, 15, 10, 11, -9, 6, 15,
    -- filter=21 channel=13
    3, 2, 7, 2, 5, -10, -3, 9, 11,
    -- filter=21 channel=14
    15, -5, -9, 13, -1, 0, -9, 12, 6,
    -- filter=21 channel=15
    -3, -8, 8, 12, -9, 5, -14, -2, 8,
    -- filter=21 channel=16
    3, 0, 2, 11, 5, -11, 11, -10, -9,
    -- filter=21 channel=17
    -12, -5, -5, -3, 5, 11, -6, -13, 8,
    -- filter=21 channel=18
    4, 8, 7, -7, -10, 0, 11, 6, 4,
    -- filter=21 channel=19
    11, -12, -7, -14, -14, 13, -14, -13, 12,
    -- filter=21 channel=20
    -6, -1, 13, -11, -1, 10, -11, 8, 8,
    -- filter=21 channel=21
    8, -6, 13, 0, -2, -10, -8, -11, 11,
    -- filter=21 channel=22
    -2, 2, 6, 14, 2, 5, 3, -7, 5,
    -- filter=21 channel=23
    10, 5, 4, 0, 11, -9, -9, 13, 10,
    -- filter=21 channel=24
    -12, -9, -3, -11, -4, -4, 11, 6, 3,
    -- filter=21 channel=25
    2, 3, 3, 8, 2, 4, -9, -3, -10,
    -- filter=21 channel=26
    -11, 0, -6, 4, -1, -13, -2, -2, -11,
    -- filter=21 channel=27
    8, -3, 8, 11, -2, -11, -13, 12, -1,
    -- filter=21 channel=28
    8, 9, 13, -5, -9, -4, 9, 4, -8,
    -- filter=21 channel=29
    -11, -7, 12, -5, 0, -1, -8, -11, 10,
    -- filter=21 channel=30
    -2, -14, 0, -4, -13, -7, 1, -14, -1,
    -- filter=21 channel=31
    9, -9, -12, -11, -5, -3, -10, -12, 9,
    -- filter=22 channel=0
    -19, -18, 5, -20, 0, -6, -13, -16, -14,
    -- filter=22 channel=1
    -1, 17, 9, 12, 7, 3, 8, 3, -15,
    -- filter=22 channel=2
    7, 8, 14, 3, -1, -5, 4, -5, 0,
    -- filter=22 channel=3
    11, -4, -3, -3, 8, -13, -13, 13, -7,
    -- filter=22 channel=4
    1, -11, 15, 2, -9, 4, 1, 8, -14,
    -- filter=22 channel=5
    -7, 11, -9, 0, 0, 12, -6, 0, 11,
    -- filter=22 channel=6
    3, -14, -4, 15, 4, 9, -5, -1, 14,
    -- filter=22 channel=7
    13, 17, -5, -3, -5, -8, -10, 4, -13,
    -- filter=22 channel=8
    9, 0, 8, -2, 11, -5, 7, 9, 7,
    -- filter=22 channel=9
    -8, -11, -1, -13, -17, -2, 2, -2, -14,
    -- filter=22 channel=10
    -3, 9, -11, -1, -5, 11, 7, -15, 7,
    -- filter=22 channel=11
    -1, -8, 6, 8, 11, 1, 0, 4, -5,
    -- filter=22 channel=12
    -6, -3, -6, 4, 1, -6, 4, -9, -19,
    -- filter=22 channel=13
    18, 11, 17, -6, 2, 2, 19, 0, 14,
    -- filter=22 channel=14
    8, 8, 3, -13, 6, 13, -15, 7, 6,
    -- filter=22 channel=15
    -11, -1, 7, 0, 7, -3, 6, 3, -4,
    -- filter=22 channel=16
    -2, 2, 17, 3, 10, 3, 9, 2, -7,
    -- filter=22 channel=17
    10, 13, 2, 17, 10, 6, -6, 1, -11,
    -- filter=22 channel=18
    14, 0, 17, -6, -9, 4, -6, 13, 7,
    -- filter=22 channel=19
    13, 11, 5, 14, 12, 4, -8, 7, -9,
    -- filter=22 channel=20
    19, -2, 5, 8, 19, 8, 13, -4, 4,
    -- filter=22 channel=21
    0, 9, -17, 2, -22, -12, -22, -28, -11,
    -- filter=22 channel=22
    -13, -11, 0, -21, -13, -6, 0, -8, -16,
    -- filter=22 channel=23
    -4, 3, -11, 8, -12, -13, -6, 2, -4,
    -- filter=22 channel=24
    0, 4, 10, 1, 9, 15, 11, 2, 11,
    -- filter=22 channel=25
    -18, -2, -11, -3, -19, -13, -16, 1, 0,
    -- filter=22 channel=26
    9, 6, 3, 15, -8, -13, -10, -6, -16,
    -- filter=22 channel=27
    9, 9, 6, 0, 11, -1, -2, 10, 0,
    -- filter=22 channel=28
    -2, 12, 4, -7, 8, -7, 0, 13, -14,
    -- filter=22 channel=29
    -1, 8, 0, 3, 0, 16, 10, 11, 11,
    -- filter=22 channel=30
    -9, -10, 12, -6, 12, 12, 6, 8, -8,
    -- filter=22 channel=31
    -2, -14, 0, 8, -10, 1, 9, -12, 2,
    -- filter=23 channel=0
    3, 9, 12, 9, 0, -7, -13, 7, 9,
    -- filter=23 channel=1
    -16, 0, -10, 11, 0, 8, 8, -13, 10,
    -- filter=23 channel=2
    -5, -11, -10, 0, -11, 1, 2, 8, -7,
    -- filter=23 channel=3
    0, 2, 6, 3, -5, 7, 6, -7, -5,
    -- filter=23 channel=4
    12, 5, 6, -1, 4, 8, 10, 21, 1,
    -- filter=23 channel=5
    15, 3, -1, 6, 12, 12, 6, 3, -13,
    -- filter=23 channel=6
    14, -7, -8, 7, 6, -7, -7, 6, -8,
    -- filter=23 channel=7
    -21, -5, -19, 3, -1, -23, -16, 4, -15,
    -- filter=23 channel=8
    -2, -1, -4, -6, 0, -12, 8, -3, -13,
    -- filter=23 channel=9
    -10, -3, -5, 10, 13, 7, -3, 14, 9,
    -- filter=23 channel=10
    -4, -10, 5, 11, -8, -8, -9, -2, 10,
    -- filter=23 channel=11
    -17, -8, -16, -23, -7, 2, 2, -6, 3,
    -- filter=23 channel=12
    -9, 9, -9, -3, -3, -12, 3, -2, -5,
    -- filter=23 channel=13
    -13, -2, 8, 14, -6, -7, -1, -7, -8,
    -- filter=23 channel=14
    -10, -4, -4, -7, -12, -12, 9, 4, 11,
    -- filter=23 channel=15
    12, 13, 4, -9, 8, 0, 7, -6, 4,
    -- filter=23 channel=16
    -8, -7, 1, 1, 10, -8, -13, 6, -3,
    -- filter=23 channel=17
    -8, -16, 5, -7, -20, 3, 2, -4, -15,
    -- filter=23 channel=18
    10, 8, 13, 14, 13, 11, -5, 15, 10,
    -- filter=23 channel=19
    12, 2, 0, 6, -8, 12, -12, -13, 9,
    -- filter=23 channel=20
    -12, -13, -19, -9, -23, -11, -14, 6, -5,
    -- filter=23 channel=21
    12, 1, -13, -3, -7, -6, 8, -13, 9,
    -- filter=23 channel=22
    -7, 12, -4, -3, 4, -1, 9, 14, -9,
    -- filter=23 channel=23
    -8, 11, 8, 6, 1, 5, 7, -2, -6,
    -- filter=23 channel=24
    -8, -10, -5, 2, -1, -1, -15, 8, -5,
    -- filter=23 channel=25
    23, 13, -7, 24, 16, -2, 25, 21, 17,
    -- filter=23 channel=26
    -9, 9, 5, -7, 1, -8, 6, -10, -4,
    -- filter=23 channel=27
    1, 11, 9, 6, 0, 4, 10, 0, 8,
    -- filter=23 channel=28
    -10, -2, 2, -3, 12, 12, 12, 12, -16,
    -- filter=23 channel=29
    -4, 9, 6, -14, -15, -4, -1, -11, -11,
    -- filter=23 channel=30
    -11, 6, 13, 4, 11, 8, 5, -6, 3,
    -- filter=23 channel=31
    -13, 15, -2, 0, -10, -13, -9, -6, 0,
    -- filter=24 channel=0
    -5, 2, -14, -22, -8, -1, -24, -13, -13,
    -- filter=24 channel=1
    9, 11, 16, 9, 5, 15, 14, -11, 10,
    -- filter=24 channel=2
    -6, -4, 7, -9, 11, -10, -8, -3, -5,
    -- filter=24 channel=3
    8, -6, -1, -3, 0, -9, -7, 4, -1,
    -- filter=24 channel=4
    -3, -8, 4, 6, -9, 7, -6, 3, -9,
    -- filter=24 channel=5
    13, -3, -6, 13, 3, -7, 4, -6, -16,
    -- filter=24 channel=6
    8, 0, -5, 9, 10, 9, 11, 5, 14,
    -- filter=24 channel=7
    -5, 1, -11, 14, 13, 1, 2, -1, -5,
    -- filter=24 channel=8
    9, 6, -13, -5, 10, 6, 5, 4, 8,
    -- filter=24 channel=9
    -8, -5, -15, 2, -11, 5, -15, 5, -1,
    -- filter=24 channel=10
    6, 0, 0, -1, 7, -13, -2, -18, 9,
    -- filter=24 channel=11
    -10, -5, 8, -17, -15, -5, 9, -13, 11,
    -- filter=24 channel=12
    -12, -16, -13, -16, 0, 6, -7, 4, 4,
    -- filter=24 channel=13
    7, -21, -2, 4, -13, -25, -15, -11, -6,
    -- filter=24 channel=14
    -7, 9, 2, -9, -11, 9, 5, -19, -4,
    -- filter=24 channel=15
    0, -2, -3, -3, -12, -16, -11, -15, -25,
    -- filter=24 channel=16
    -2, 9, 9, 7, 10, -12, -4, -15, 5,
    -- filter=24 channel=17
    25, 7, -10, 8, 13, 2, 12, 11, -5,
    -- filter=24 channel=18
    2, -4, -12, -17, -9, 10, -5, -13, 10,
    -- filter=24 channel=19
    7, 14, 0, 7, 11, 0, 0, 4, 8,
    -- filter=24 channel=20
    17, 0, 14, 23, 21, -1, 18, 11, 16,
    -- filter=24 channel=21
    10, -12, 8, 2, -8, 3, 19, 4, 5,
    -- filter=24 channel=22
    -21, -24, -18, -5, -11, -8, 6, -22, -8,
    -- filter=24 channel=23
    9, -2, -16, 9, -11, 0, 11, -7, 11,
    -- filter=24 channel=24
    -13, 13, 8, 4, -6, 14, 10, 3, 8,
    -- filter=24 channel=25
    -4, -2, 10, 5, 3, -4, -6, -15, 12,
    -- filter=24 channel=26
    8, -11, -15, 9, -17, -25, -13, 5, -9,
    -- filter=24 channel=27
    -6, -8, -14, 10, 0, 0, 10, 6, -11,
    -- filter=24 channel=28
    -9, 13, 5, -5, 11, -6, 11, -6, -11,
    -- filter=24 channel=29
    3, 6, 10, -9, -2, -4, -5, -10, -15,
    -- filter=24 channel=30
    0, -15, 10, 5, 9, 0, 10, 13, 4,
    -- filter=24 channel=31
    3, 1, 0, 3, -21, 0, -9, -14, 0,
    -- filter=25 channel=0
    -1, 5, 8, -8, 6, 6, -7, 12, -14,
    -- filter=25 channel=1
    6, -5, 4, 7, 8, 14, -1, 12, -13,
    -- filter=25 channel=2
    -10, 1, 7, -10, -9, 4, 0, -12, 12,
    -- filter=25 channel=3
    -3, 7, -6, -4, 10, -11, 10, -14, 8,
    -- filter=25 channel=4
    -10, -11, -4, -6, 14, 12, 0, 4, -4,
    -- filter=25 channel=5
    7, 5, -1, -1, -3, 2, 9, -6, 2,
    -- filter=25 channel=6
    1, -12, 14, 11, -3, 8, 12, 11, -7,
    -- filter=25 channel=7
    -9, -13, -14, 1, 4, 12, 0, -7, -10,
    -- filter=25 channel=8
    3, 1, -8, 2, -5, -6, 6, 1, 10,
    -- filter=25 channel=9
    5, -10, -13, -13, -1, 7, 1, -6, 0,
    -- filter=25 channel=10
    -13, 5, -12, -11, -10, 4, 8, 8, 8,
    -- filter=25 channel=11
    2, -1, -6, -10, 9, -6, 4, -4, 8,
    -- filter=25 channel=12
    13, -2, -10, -9, 13, 0, 6, -14, -6,
    -- filter=25 channel=13
    0, -4, 2, 11, -13, 0, -7, 12, 5,
    -- filter=25 channel=14
    -9, -6, -7, 7, -7, 8, -6, 12, 1,
    -- filter=25 channel=15
    -13, 0, 12, 7, -12, 11, 13, 13, -8,
    -- filter=25 channel=16
    -14, -2, 1, -4, 3, -5, -10, 0, 2,
    -- filter=25 channel=17
    2, 11, 0, -13, 7, -1, 6, 9, -2,
    -- filter=25 channel=18
    -12, -8, -8, 0, 6, -2, 12, 0, -2,
    -- filter=25 channel=19
    8, 8, -7, -8, 8, 13, -3, -1, -2,
    -- filter=25 channel=20
    -3, 4, 14, -14, -2, -3, -8, -14, -5,
    -- filter=25 channel=21
    9, -3, 0, 9, -12, -7, -5, -13, 4,
    -- filter=25 channel=22
    -3, 13, -1, 4, -9, -14, 10, 13, -10,
    -- filter=25 channel=23
    14, 6, 3, 0, -7, -11, 7, 2, 12,
    -- filter=25 channel=24
    0, 0, -2, -5, -1, 7, -10, -9, 2,
    -- filter=25 channel=25
    4, 3, -8, 4, -13, -4, -12, 6, 11,
    -- filter=25 channel=26
    -6, 2, 3, -13, 11, 10, 13, -13, -2,
    -- filter=25 channel=27
    13, -7, 13, 8, 9, -7, -11, 7, 4,
    -- filter=25 channel=28
    14, -10, 4, -9, -14, -12, 0, 12, 2,
    -- filter=25 channel=29
    0, 0, -12, -6, 7, -8, 12, 0, 10,
    -- filter=25 channel=30
    -13, -14, -4, -6, -13, 5, -5, -13, -2,
    -- filter=25 channel=31
    5, -10, 3, -3, 11, -2, -6, -12, 7,
    -- filter=26 channel=0
    11, -2, -11, 8, 0, -4, 7, 1, 1,
    -- filter=26 channel=1
    -2, -3, 16, 0, 0, 7, -15, 19, 22,
    -- filter=26 channel=2
    0, -5, 6, 12, 1, 1, 2, -10, 14,
    -- filter=26 channel=3
    -9, 14, 14, 11, 14, -10, 4, -10, 6,
    -- filter=26 channel=4
    -19, 8, 0, -10, -3, 2, -15, -2, 4,
    -- filter=26 channel=5
    1, -7, -16, -9, -13, -4, -12, -1, 4,
    -- filter=26 channel=6
    3, 2, -2, -9, -6, 5, 13, 13, -9,
    -- filter=26 channel=7
    -13, -9, 18, -12, -12, 23, -4, 8, 23,
    -- filter=26 channel=8
    13, 1, 7, 0, -11, -7, 5, -9, -14,
    -- filter=26 channel=9
    -17, -2, -17, -3, 1, -15, -8, 3, -11,
    -- filter=26 channel=10
    7, 2, -8, 6, -3, 1, 0, 9, -10,
    -- filter=26 channel=11
    16, 6, -8, 25, 24, 13, 23, 19, 14,
    -- filter=26 channel=12
    -17, 4, 5, -10, 9, -3, -13, -15, -4,
    -- filter=26 channel=13
    -1, -4, 4, -11, -12, 0, -23, 5, 13,
    -- filter=26 channel=14
    0, 17, 14, -4, 23, 6, 20, 15, 3,
    -- filter=26 channel=15
    -10, 0, -12, -13, -18, -7, -8, -14, 10,
    -- filter=26 channel=16
    7, 16, 17, -10, 13, 7, -9, 9, -7,
    -- filter=26 channel=17
    -20, -5, -11, -26, -20, 0, -3, -9, -5,
    -- filter=26 channel=18
    13, -8, -6, 2, -12, 9, -2, -2, -8,
    -- filter=26 channel=19
    -13, -3, 4, 2, 12, 13, -8, 10, 4,
    -- filter=26 channel=20
    11, -3, 9, -11, 17, 31, -6, 7, 29,
    -- filter=26 channel=21
    -6, -6, -3, -21, -21, 5, -10, -15, -7,
    -- filter=26 channel=22
    -16, -3, -19, 3, -17, -7, -20, -16, -20,
    -- filter=26 channel=23
    1, -17, -11, -9, 10, -8, -7, 5, -16,
    -- filter=26 channel=24
    0, 3, 25, 4, 17, 24, 20, 18, 25,
    -- filter=26 channel=25
    -13, -18, 8, -21, -15, -11, -10, -14, -16,
    -- filter=26 channel=26
    -17, -2, -16, -1, -14, -10, -3, -18, -18,
    -- filter=26 channel=27
    11, 0, 9, -5, -5, 6, -7, 4, -10,
    -- filter=26 channel=28
    0, 8, -3, 0, -10, 0, 9, 2, 15,
    -- filter=26 channel=29
    19, 16, -8, 2, 8, 4, 15, -2, -11,
    -- filter=26 channel=30
    13, -12, -11, 5, 14, -11, 8, 9, -12,
    -- filter=26 channel=31
    -19, -5, -2, -14, -11, 0, -5, -7, 7,
    -- filter=27 channel=0
    -9, 12, -2, -14, 11, -12, 13, 15, -1,
    -- filter=27 channel=1
    -10, 3, 4, -3, -7, 13, 2, 2, -8,
    -- filter=27 channel=2
    14, 8, -3, -5, -2, -12, -2, -11, 0,
    -- filter=27 channel=3
    -6, -10, 10, -6, -12, -2, 13, -11, 11,
    -- filter=27 channel=4
    -1, -13, 8, -11, 11, 0, 13, 4, 1,
    -- filter=27 channel=5
    -5, -11, -12, 10, 12, 11, -11, 9, 9,
    -- filter=27 channel=6
    6, -4, 4, 0, 0, -8, -9, -13, 4,
    -- filter=27 channel=7
    15, -9, -14, 2, 8, 0, 9, -12, -2,
    -- filter=27 channel=8
    8, 7, 4, 7, 13, 14, 11, 6, -12,
    -- filter=27 channel=9
    -11, 4, 9, 6, 11, -9, 12, 14, 10,
    -- filter=27 channel=10
    15, 9, 8, -3, -6, 11, 0, -1, -8,
    -- filter=27 channel=11
    -6, 12, -4, 5, -11, -12, 2, -3, 15,
    -- filter=27 channel=12
    9, 0, -14, 7, 3, 0, 9, 14, -4,
    -- filter=27 channel=13
    10, -10, -9, -2, 10, 4, -1, -3, -3,
    -- filter=27 channel=14
    8, 3, -11, -5, 6, 9, -8, -8, -3,
    -- filter=27 channel=15
    -1, 4, 4, 1, 7, 14, -11, -5, 6,
    -- filter=27 channel=16
    -10, -10, 0, 14, 6, -13, 0, 1, 7,
    -- filter=27 channel=17
    -3, -7, 9, 5, 10, 3, -11, -9, -11,
    -- filter=27 channel=18
    0, 5, -7, -10, -2, -13, 2, 2, 12,
    -- filter=27 channel=19
    5, 6, 4, -2, 3, 0, 13, -4, 1,
    -- filter=27 channel=20
    2, 5, -15, -12, -10, -15, -13, -6, 6,
    -- filter=27 channel=21
    12, 12, -7, 14, -9, -8, -14, 11, 3,
    -- filter=27 channel=22
    3, 10, 7, 0, -8, 14, -4, 3, -11,
    -- filter=27 channel=23
    13, -5, 10, 2, 7, -3, -10, 14, -12,
    -- filter=27 channel=24
    1, -6, -8, -5, 3, -15, -2, 12, 12,
    -- filter=27 channel=25
    6, 6, -9, -6, -5, -7, 6, -12, 11,
    -- filter=27 channel=26
    16, 13, 0, -11, -4, -7, 11, 14, -1,
    -- filter=27 channel=27
    14, -7, 15, -10, -10, 6, 0, -3, 2,
    -- filter=27 channel=28
    -3, -9, -4, -10, 10, 2, -4, 0, -11,
    -- filter=27 channel=29
    -9, 9, -12, -5, 1, 15, -5, -3, 2,
    -- filter=27 channel=30
    12, -2, 0, -13, -5, -11, 7, 1, -3,
    -- filter=27 channel=31
    -7, -9, -9, -7, 10, 3, 6, -14, 1,
    -- filter=28 channel=0
    -8, -1, 3, -9, 0, 6, -1, -13, 3,
    -- filter=28 channel=1
    -7, -8, 0, -4, -10, -2, -5, -1, -11,
    -- filter=28 channel=2
    14, 2, -3, 3, 9, -5, -14, 4, -7,
    -- filter=28 channel=3
    8, 0, 5, 13, -5, 12, 2, -11, -12,
    -- filter=28 channel=4
    6, 7, -13, 0, 3, 14, -1, 11, -7,
    -- filter=28 channel=5
    -4, -11, -4, 0, 1, 14, 8, 15, 11,
    -- filter=28 channel=6
    3, 7, 4, 14, 4, -6, 13, -6, -13,
    -- filter=28 channel=7
    -6, 1, -15, 16, -5, -4, 5, 12, -3,
    -- filter=28 channel=8
    -10, 1, -3, -8, 2, -13, 8, 9, 14,
    -- filter=28 channel=9
    -14, 8, 2, -4, -7, -7, -6, 2, -8,
    -- filter=28 channel=10
    1, -2, 5, 10, 5, 13, -1, -9, -9,
    -- filter=28 channel=11
    6, 11, 15, 2, -12, -9, 4, -7, -1,
    -- filter=28 channel=12
    -13, -12, 1, 12, 8, -6, 10, 11, -9,
    -- filter=28 channel=13
    -14, -12, 2, 11, 6, 7, -8, 3, 3,
    -- filter=28 channel=14
    -15, 1, 7, -6, -9, -10, -2, -1, -14,
    -- filter=28 channel=15
    10, 3, -10, -7, 10, -5, -9, -4, -4,
    -- filter=28 channel=16
    -8, -1, 4, 1, -7, 5, 0, 13, 6,
    -- filter=28 channel=17
    12, 2, -5, -7, -9, -11, 16, 10, -6,
    -- filter=28 channel=18
    3, 13, -1, 0, 13, 9, 0, 4, 6,
    -- filter=28 channel=19
    5, -9, 3, 3, 14, -5, 7, 3, -13,
    -- filter=28 channel=20
    -11, -10, -7, 5, 12, -2, 0, 1, -6,
    -- filter=28 channel=21
    8, -9, -17, 8, 14, -2, 15, 8, 9,
    -- filter=28 channel=22
    13, 6, 0, 1, 3, -14, 14, 6, 7,
    -- filter=28 channel=23
    8, -5, 12, 9, -7, -15, -12, -2, 2,
    -- filter=28 channel=24
    -1, -14, 6, -9, 11, 2, -2, -2, 9,
    -- filter=28 channel=25
    0, 6, -10, 6, -6, 7, -13, 10, 1,
    -- filter=28 channel=26
    -8, -11, 6, 6, -10, 11, -9, 13, 1,
    -- filter=28 channel=27
    -4, -14, -7, 12, 8, 1, 4, 9, 14,
    -- filter=28 channel=28
    2, -2, 13, 1, -10, 6, 17, 6, 5,
    -- filter=28 channel=29
    -7, 2, 0, 14, 3, 4, 4, 1, 13,
    -- filter=28 channel=30
    -11, 0, -6, 7, -1, -2, -1, -10, -1,
    -- filter=28 channel=31
    6, 8, -17, -10, -7, 2, 16, 3, -8,
    -- filter=29 channel=0
    13, -10, -10, -7, 1, 6, 9, -13, 9,
    -- filter=29 channel=1
    13, -11, -4, -7, 10, 13, -7, -8, -2,
    -- filter=29 channel=2
    -6, -11, -9, 2, 11, -14, 10, -1, -13,
    -- filter=29 channel=3
    5, 6, 1, -6, 12, -2, -4, 12, -2,
    -- filter=29 channel=4
    5, -1, 14, 3, -5, -9, 7, -8, -12,
    -- filter=29 channel=5
    -4, 9, 4, -8, 0, -3, -6, -4, -9,
    -- filter=29 channel=6
    -10, -14, 13, 0, 13, -13, -1, 12, 8,
    -- filter=29 channel=7
    -8, 14, 8, -7, -7, 6, 14, -13, 12,
    -- filter=29 channel=8
    -14, -14, 7, -7, 2, 3, 10, 14, -7,
    -- filter=29 channel=9
    14, -8, 5, 7, 2, -2, -3, -2, -3,
    -- filter=29 channel=10
    -6, -1, -9, 6, -1, -7, 9, -7, -6,
    -- filter=29 channel=11
    8, -1, -10, 14, -2, -14, -10, -12, -14,
    -- filter=29 channel=12
    10, -10, -3, -6, 8, -12, -13, 11, -7,
    -- filter=29 channel=13
    -13, -2, -4, 10, 0, 0, 0, -14, 9,
    -- filter=29 channel=14
    2, 2, -4, -4, -1, 3, -8, 1, -2,
    -- filter=29 channel=15
    1, -10, -10, 12, -7, -4, 0, 11, -8,
    -- filter=29 channel=16
    13, 14, 7, 10, 10, -4, -5, 4, -11,
    -- filter=29 channel=17
    5, -9, 2, -9, -6, -9, -4, -5, -1,
    -- filter=29 channel=18
    6, -10, -10, 1, 12, 11, 0, -4, 2,
    -- filter=29 channel=19
    -5, 2, -6, 14, 2, 0, -11, 0, 0,
    -- filter=29 channel=20
    12, 14, -3, -12, 8, 14, 7, -6, 2,
    -- filter=29 channel=21
    12, 8, -12, 10, 0, -14, -14, 0, 0,
    -- filter=29 channel=22
    9, 4, -5, -9, 10, -6, -10, -4, -12,
    -- filter=29 channel=23
    -13, 13, -4, -10, -1, 11, 8, 10, 5,
    -- filter=29 channel=24
    12, -13, -4, 9, -5, 7, -9, -1, 4,
    -- filter=29 channel=25
    -3, 1, 1, 12, -11, 6, -12, -4, -15,
    -- filter=29 channel=26
    -8, 1, 10, 3, 10, 0, -5, -9, -3,
    -- filter=29 channel=27
    6, -8, 11, 7, 0, -12, -7, 5, 12,
    -- filter=29 channel=28
    1, 2, -14, -11, 9, 5, -8, -9, 4,
    -- filter=29 channel=29
    8, -4, 0, 8, 0, -10, -8, -1, 0,
    -- filter=29 channel=30
    12, -11, -1, 0, -11, -5, -9, -6, -12,
    -- filter=29 channel=31
    -14, -4, -13, 3, 14, -5, -14, -8, 1,
    -- filter=30 channel=0
    -12, -17, 3, -9, 0, -3, -6, -10, -4,
    -- filter=30 channel=1
    14, 0, 14, 14, 0, 12, 6, 11, 3,
    -- filter=30 channel=2
    -7, -4, -12, -6, 0, 12, 13, 0, -5,
    -- filter=30 channel=3
    6, 5, -11, 14, 13, -6, 10, -10, -12,
    -- filter=30 channel=4
    8, 5, -12, -16, 4, -2, -12, -8, -4,
    -- filter=30 channel=5
    -3, 0, -6, -2, -13, 0, 11, -11, -12,
    -- filter=30 channel=6
    -7, 2, 11, -2, 6, 0, 0, -7, 3,
    -- filter=30 channel=7
    2, -13, 7, -19, -10, -4, -22, -4, 0,
    -- filter=30 channel=8
    2, 5, -7, -5, 3, -2, 7, -3, 0,
    -- filter=30 channel=9
    -18, 5, -3, -12, 4, -6, 4, 7, -4,
    -- filter=30 channel=10
    -9, -2, -15, 4, 11, -4, 2, -12, 12,
    -- filter=30 channel=11
    0, 1, 0, -3, 0, 7, 8, 13, 17,
    -- filter=30 channel=12
    0, -6, 4, -4, -15, -9, -20, -15, 0,
    -- filter=30 channel=13
    -5, 18, 13, 3, 9, 9, 6, 7, 20,
    -- filter=30 channel=14
    9, 17, -2, 13, 6, 3, 8, 0, 13,
    -- filter=30 channel=15
    9, -10, 12, 5, -9, 0, -14, 11, -4,
    -- filter=30 channel=16
    9, 5, 10, 11, 7, 3, 0, 20, 10,
    -- filter=30 channel=17
    12, 0, -13, 10, -19, -7, -8, -15, -4,
    -- filter=30 channel=18
    15, 19, 21, 22, -3, 20, 17, 0, 9,
    -- filter=30 channel=19
    -11, 2, -8, 0, -9, 5, 13, 9, -6,
    -- filter=30 channel=20
    1, 21, 24, 22, 30, 12, 23, 14, 30,
    -- filter=30 channel=21
    -8, 0, -8, -15, -16, -18, -9, -32, -24,
    -- filter=30 channel=22
    -23, -12, -13, -27, -9, -10, -20, -28, -22,
    -- filter=30 channel=23
    1, -7, -16, 6, -19, -8, -19, 5, -18,
    -- filter=30 channel=24
    13, -2, 17, 0, 13, 27, 3, 24, 19,
    -- filter=30 channel=25
    -26, -22, -13, -29, -30, -26, -36, -29, -11,
    -- filter=30 channel=26
    -4, 10, 4, 2, -16, 0, 2, 9, -9,
    -- filter=30 channel=27
    -4, 11, 13, 9, -8, -6, 4, 3, -4,
    -- filter=30 channel=28
    14, 13, 14, -3, 15, -5, 9, 13, 4,
    -- filter=30 channel=29
    17, 15, -1, 6, 13, -3, 18, 2, 21,
    -- filter=30 channel=30
    2, 0, 0, 9, 6, -4, 11, 11, -14,
    -- filter=30 channel=31
    -5, 7, -15, -18, 1, -10, -2, -19, 1,
    -- filter=31 channel=0
    -5, -7, -9, -2, -2, 5, -11, -5, -6,
    -- filter=31 channel=1
    3, 3, 3, -1, -13, -14, 13, 3, 11,
    -- filter=31 channel=2
    13, 8, 0, -9, 0, 7, 15, -14, -9,
    -- filter=31 channel=3
    0, -14, -9, -2, 5, -5, 10, -7, 7,
    -- filter=31 channel=4
    1, 9, 4, 0, -2, 14, -1, 0, 0,
    -- filter=31 channel=5
    -2, -7, 2, -3, 9, -13, 7, -9, -6,
    -- filter=31 channel=6
    7, 0, 3, 9, -9, -12, -7, -13, 5,
    -- filter=31 channel=7
    6, -3, -14, -13, -6, -14, 6, -8, -2,
    -- filter=31 channel=8
    -9, -10, -11, -4, 7, 14, -7, -8, 5,
    -- filter=31 channel=9
    7, 3, 13, -3, -10, 11, -13, 9, -7,
    -- filter=31 channel=10
    -11, -7, 12, -1, 10, -9, 11, 11, -2,
    -- filter=31 channel=11
    -11, -3, 1, -1, 9, -14, 4, 2, 6,
    -- filter=31 channel=12
    5, -14, 3, -1, -14, 0, 12, -10, 9,
    -- filter=31 channel=13
    -10, 0, 9, -10, -3, 10, 3, -2, 1,
    -- filter=31 channel=14
    -9, -3, -3, -3, 4, 1, 4, -5, 2,
    -- filter=31 channel=15
    -7, -9, 10, -2, -8, -9, -9, -1, -13,
    -- filter=31 channel=16
    -12, -9, 13, -6, -11, 1, 11, 9, -13,
    -- filter=31 channel=17
    0, 3, -13, 12, 0, -9, -2, -6, -11,
    -- filter=31 channel=18
    9, 4, -2, -14, 3, -3, -5, -5, 4,
    -- filter=31 channel=19
    10, -9, 6, 0, -6, -3, 9, 10, -6,
    -- filter=31 channel=20
    -9, -8, -11, 6, 5, 13, -2, 11, 11,
    -- filter=31 channel=21
    2, 8, 5, 8, 13, 8, -7, -14, 4,
    -- filter=31 channel=22
    -9, -11, -1, 2, -5, 0, -4, 7, 8,
    -- filter=31 channel=23
    12, 7, -6, -4, 5, -7, 0, -13, -7,
    -- filter=31 channel=24
    11, 0, 8, 6, 2, 14, -2, -5, 1,
    -- filter=31 channel=25
    -7, -9, -12, 1, -11, -5, -3, 4, -9,
    -- filter=31 channel=26
    3, 14, 6, -2, -12, 9, 4, 7, -2,
    -- filter=31 channel=27
    -9, -12, 8, 2, 12, -8, -5, 7, -4,
    -- filter=31 channel=28
    1, -14, -1, 14, 1, -9, -3, 3, -11,
    -- filter=31 channel=29
    -14, -9, -8, -1, 3, -8, -9, 11, -11,
    -- filter=31 channel=30
    2, -10, -12, -4, 5, 6, 9, -2, -13,
    -- filter=31 channel=31
    -1, 8, 1, -14, -7, -1, -11, -7, -5,
    -- filter=32 channel=0
    -15, -9, 5, -17, -9, -8, 0, 1, -15,
    -- filter=32 channel=1
    4, 16, 2, -8, 17, 13, 5, -2, 15,
    -- filter=32 channel=2
    -1, -11, -3, 6, 14, 6, 8, 0, -10,
    -- filter=32 channel=3
    13, -2, 12, -8, 9, -8, 5, -2, 12,
    -- filter=32 channel=4
    -12, -13, 1, 11, 1, 0, -12, -13, 14,
    -- filter=32 channel=5
    -6, -4, 12, 12, -15, 1, 6, 0, 11,
    -- filter=32 channel=6
    14, -8, -7, -9, -13, 10, 14, 12, 0,
    -- filter=32 channel=7
    20, 6, 16, 2, 10, -6, 12, 9, 5,
    -- filter=32 channel=8
    10, -10, 0, 5, 5, 2, -9, 9, -8,
    -- filter=32 channel=9
    7, 9, 7, -5, -9, -14, 11, 4, -5,
    -- filter=32 channel=10
    -2, -4, -2, -1, -17, -4, -2, -15, -6,
    -- filter=32 channel=11
    -18, -17, -14, 2, -11, -4, -20, -3, -12,
    -- filter=32 channel=12
    -1, -7, 1, 0, 11, 14, 7, -3, -13,
    -- filter=32 channel=13
    -16, -6, -4, -12, -6, 9, -23, -22, -12,
    -- filter=32 channel=14
    6, -11, -7, 8, -15, -12, -1, 1, -3,
    -- filter=32 channel=15
    5, 0, -14, -11, -6, 4, -17, 0, -13,
    -- filter=32 channel=16
    13, 11, 0, 6, 9, 9, -13, 8, -12,
    -- filter=32 channel=17
    14, 3, 5, -11, 14, -6, -1, -7, 6,
    -- filter=32 channel=18
    5, -15, 5, 8, -6, 3, 9, 1, 15,
    -- filter=32 channel=19
    -2, 2, 7, 14, 13, 10, 14, 12, 10,
    -- filter=32 channel=20
    9, 20, 6, 0, -5, 6, -4, 14, 19,
    -- filter=32 channel=21
    20, 15, 12, -11, 10, 5, 3, -5, -12,
    -- filter=32 channel=22
    -6, -11, -17, -12, -20, 7, -16, 2, -12,
    -- filter=32 channel=23
    -15, -15, 2, 10, -2, -11, -9, -3, -7,
    -- filter=32 channel=24
    -9, -6, 12, -2, 0, 14, 9, -16, 14,
    -- filter=32 channel=25
    -5, -7, 2, 5, 11, -14, 15, 8, -3,
    -- filter=32 channel=26
    -6, -6, 3, -15, -22, -4, -4, -2, -5,
    -- filter=32 channel=27
    14, 0, 1, -5, -8, 0, -6, -6, -6,
    -- filter=32 channel=28
    -3, -1, -11, 0, -3, 6, -5, -1, -7,
    -- filter=32 channel=29
    -17, -14, -8, -21, -20, 0, -20, -16, -6,
    -- filter=32 channel=30
    8, 8, 2, 0, 13, 4, -10, -10, 1,
    -- filter=32 channel=31
    -6, 3, -1, 9, 6, 6, -11, -11, -15,
    -- filter=33 channel=0
    -7, -10, 12, 1, 13, 16, 8, -7, 4,
    -- filter=33 channel=1
    -8, 0, -10, 9, 7, -19, -6, 9, 5,
    -- filter=33 channel=2
    2, 12, 13, 1, 1, -4, 10, -10, -13,
    -- filter=33 channel=3
    -3, -8, -12, 0, -13, 12, -12, 15, -11,
    -- filter=33 channel=4
    8, 12, 9, 12, -11, 4, 3, 16, -8,
    -- filter=33 channel=5
    -13, -1, 3, -12, 0, -14, 5, 9, -12,
    -- filter=33 channel=6
    -7, 0, -2, 7, -4, -6, -3, 5, 0,
    -- filter=33 channel=7
    -15, -20, 7, -7, -17, -20, -19, -18, 0,
    -- filter=33 channel=8
    3, 0, 6, -13, -3, -2, -11, 8, 8,
    -- filter=33 channel=9
    -7, -2, -10, 1, 10, 4, 7, 13, -4,
    -- filter=33 channel=10
    -9, 12, -11, 17, 0, 1, -9, -12, -2,
    -- filter=33 channel=11
    8, 1, 4, -21, -13, -4, -1, -15, -8,
    -- filter=33 channel=12
    10, -8, -9, 8, 13, 14, -13, 5, 5,
    -- filter=33 channel=13
    -7, -11, -5, -14, -8, 5, -3, 8, -2,
    -- filter=33 channel=14
    12, -10, 3, -5, 2, 1, 11, 0, 1,
    -- filter=33 channel=15
    2, -7, -7, -3, -3, 14, 14, -3, 8,
    -- filter=33 channel=16
    -1, -10, 4, -7, 7, -16, -15, -1, 2,
    -- filter=33 channel=17
    -12, 9, -1, 10, 0, -14, -8, -9, -9,
    -- filter=33 channel=18
    13, 11, 0, 3, -10, 13, 16, -9, 8,
    -- filter=33 channel=19
    -4, -10, -3, 11, 7, 13, 0, -7, 5,
    -- filter=33 channel=20
    -6, -16, -7, -4, 0, -4, -16, -14, -12,
    -- filter=33 channel=21
    0, 3, -15, 3, -8, -10, -9, -4, 9,
    -- filter=33 channel=22
    -6, -2, 1, 14, 14, 12, 15, -9, 4,
    -- filter=33 channel=23
    -9, -7, -10, 15, 10, -10, -2, 4, -7,
    -- filter=33 channel=24
    10, -16, 2, -1, -10, -14, -9, -15, -11,
    -- filter=33 channel=25
    21, 10, 4, 24, 20, 16, 4, 12, 14,
    -- filter=33 channel=26
    -6, -5, 1, -1, -14, 11, 9, 0, -12,
    -- filter=33 channel=27
    13, 3, -7, -3, 0, -13, 13, 12, 2,
    -- filter=33 channel=28
    1, -8, 11, -3, -1, -4, 0, 4, -7,
    -- filter=33 channel=29
    3, -1, -5, -13, -7, -19, -2, 9, 5,
    -- filter=33 channel=30
    -13, -10, -12, 1, 2, -7, 1, 0, -13,
    -- filter=33 channel=31
    11, -5, -14, 6, -13, 10, 13, -13, 6,
    -- filter=34 channel=0
    12, -10, 7, 13, 3, 8, 6, 9, 12,
    -- filter=34 channel=1
    -10, -17, -2, -4, -10, -14, 3, 6, 0,
    -- filter=34 channel=2
    -2, 0, 0, 10, -1, 3, 8, -9, -2,
    -- filter=34 channel=3
    -9, 15, 5, 10, 13, 0, 6, 4, -10,
    -- filter=34 channel=4
    -9, -12, -3, 8, 13, 0, -12, 10, 0,
    -- filter=34 channel=5
    -9, 11, 6, -10, 6, -16, 0, -3, -15,
    -- filter=34 channel=6
    4, 14, -6, 13, -12, 0, -4, 9, 0,
    -- filter=34 channel=7
    -9, -2, 2, 0, 7, 10, 7, 4, -4,
    -- filter=34 channel=8
    7, 13, 8, -9, 7, -8, -4, 0, 11,
    -- filter=34 channel=9
    -5, 9, -4, 14, 18, 16, -6, 3, 2,
    -- filter=34 channel=10
    12, 5, -1, -5, 14, 0, -2, -5, -1,
    -- filter=34 channel=11
    10, -9, 1, -6, -5, -9, 8, 2, -7,
    -- filter=34 channel=12
    11, -2, 22, 1, 7, 18, -3, -5, -10,
    -- filter=34 channel=13
    -9, 5, -8, 8, -5, -11, -11, -13, -13,
    -- filter=34 channel=14
    -13, -12, -9, 10, -7, 8, -9, -1, 13,
    -- filter=34 channel=15
    -4, 0, 11, 13, 11, 8, -1, -11, -2,
    -- filter=34 channel=16
    -2, 1, 3, -9, 5, -1, 11, -6, -5,
    -- filter=34 channel=17
    -10, 14, 7, 5, -16, -17, 5, -15, -20,
    -- filter=34 channel=18
    7, -7, 7, -12, 0, -14, 8, 9, 14,
    -- filter=34 channel=19
    -10, 0, -9, -4, 14, 3, 7, 5, -11,
    -- filter=34 channel=20
    -6, 1, 1, -6, -6, 6, -8, 6, -16,
    -- filter=34 channel=21
    0, -6, -8, 8, 8, 0, 5, -12, 9,
    -- filter=34 channel=22
    21, 16, 10, 13, 28, 7, 26, 25, 19,
    -- filter=34 channel=23
    -5, -9, 4, -6, 15, -4, 0, -6, 8,
    -- filter=34 channel=24
    -4, -16, -16, -18, -14, -4, -14, 7, -5,
    -- filter=34 channel=25
    7, 11, 10, -8, 4, 14, 17, 14, 12,
    -- filter=34 channel=26
    14, 10, 5, -9, 0, 11, -9, 5, 0,
    -- filter=34 channel=27
    -14, -9, 0, 11, 2, -6, 11, 12, 3,
    -- filter=34 channel=28
    -1, 9, 14, -12, -13, 13, 6, -14, -5,
    -- filter=34 channel=29
    0, -5, -5, 10, 4, -3, 6, 9, -3,
    -- filter=34 channel=30
    6, 14, 1, -2, -12, -1, -9, 13, -6,
    -- filter=34 channel=31
    -2, 3, 14, 4, -8, 0, 12, -6, -16,
    -- filter=35 channel=0
    0, 10, -2, 0, -14, -7, 12, 14, -10,
    -- filter=35 channel=1
    -12, -15, -1, -11, 3, 0, 2, 3, -14,
    -- filter=35 channel=2
    -5, -10, 6, 8, 6, -11, 1, 10, -11,
    -- filter=35 channel=3
    14, -8, 10, 13, 2, -7, 11, 0, -13,
    -- filter=35 channel=4
    19, 7, 4, 17, 7, -11, 17, 10, 13,
    -- filter=35 channel=5
    -2, 7, 4, -14, 8, 9, -5, -12, -14,
    -- filter=35 channel=6
    14, 4, 5, 3, -2, -8, -5, 0, 10,
    -- filter=35 channel=7
    5, -15, 10, -16, -1, -17, -13, 1, 7,
    -- filter=35 channel=8
    3, 14, 3, 3, -1, -12, 4, 14, 9,
    -- filter=35 channel=9
    -4, -5, 3, 13, -13, 4, -7, -3, 5,
    -- filter=35 channel=10
    13, 16, 14, 17, -6, -1, 10, 0, -7,
    -- filter=35 channel=11
    -3, 8, 4, -3, -1, -3, 0, -14, -13,
    -- filter=35 channel=12
    0, -11, -10, -6, -6, -1, -12, 12, -12,
    -- filter=35 channel=13
    9, 13, -10, -12, -10, -2, 8, -4, 10,
    -- filter=35 channel=14
    -1, -4, -9, -4, 7, -2, -5, 0, -16,
    -- filter=35 channel=15
    -2, -14, 13, 6, -10, -6, -2, 4, 8,
    -- filter=35 channel=16
    -8, -9, 9, -11, -2, 10, -4, -2, -8,
    -- filter=35 channel=17
    -5, 7, -10, 0, 0, -13, 13, -7, 8,
    -- filter=35 channel=18
    13, 12, 7, -7, 3, -13, 15, 8, -5,
    -- filter=35 channel=19
    -6, 14, -1, 0, 12, 11, 7, 13, -10,
    -- filter=35 channel=20
    0, -3, -10, 10, -3, -20, -3, 2, -15,
    -- filter=35 channel=21
    -4, -3, -9, 7, 8, -15, 7, 15, -4,
    -- filter=35 channel=22
    10, -6, -2, 15, 12, -10, -4, -1, 9,
    -- filter=35 channel=23
    10, -12, -5, 12, -4, -1, -3, 8, 4,
    -- filter=35 channel=24
    6, -8, -1, -12, -15, -7, 7, 8, 0,
    -- filter=35 channel=25
    2, 7, 3, 19, 8, 2, 13, 0, -8,
    -- filter=35 channel=26
    3, 11, -7, 11, -7, -9, -4, -12, -4,
    -- filter=35 channel=27
    9, -1, 2, -13, 4, 9, 9, 5, 3,
    -- filter=35 channel=28
    6, -13, 7, -7, -13, -13, -6, -11, -8,
    -- filter=35 channel=29
    -6, -4, 11, -9, -11, -7, -17, -2, -4,
    -- filter=35 channel=30
    4, -1, 14, -2, 4, 7, -14, 10, 9,
    -- filter=35 channel=31
    2, -14, -11, -9, -9, 11, 4, -5, 0,
    -- filter=36 channel=0
    17, 12, 17, 15, -1, 4, 16, 8, 11,
    -- filter=36 channel=1
    2, 0, 6, 10, -10, -16, -6, -5, -15,
    -- filter=36 channel=2
    -1, 4, 2, -3, 1, 2, 6, -6, 4,
    -- filter=36 channel=3
    5, 4, -13, 9, 0, 7, -1, -8, -5,
    -- filter=36 channel=4
    -13, 7, 0, 14, 4, -11, 0, 0, 5,
    -- filter=36 channel=5
    -1, 8, -4, 8, -8, 9, -3, -12, 12,
    -- filter=36 channel=6
    -1, -9, 1, -6, -2, 1, 1, 2, -11,
    -- filter=36 channel=7
    8, -7, -10, 3, 12, -3, -9, -18, 9,
    -- filter=36 channel=8
    5, -4, 2, 1, -10, 10, 0, 12, -7,
    -- filter=36 channel=9
    7, 11, -5, 11, 2, -2, 15, -9, -5,
    -- filter=36 channel=10
    7, -10, -5, -4, -3, 1, 0, 12, -5,
    -- filter=36 channel=11
    0, 14, 20, 11, -5, 0, 11, 20, -8,
    -- filter=36 channel=12
    -4, 7, -1, -5, 0, 11, -3, 0, 6,
    -- filter=36 channel=13
    -5, -11, -9, 2, 11, -10, -5, -9, -5,
    -- filter=36 channel=14
    14, -4, 3, 12, -6, -13, -1, 14, 1,
    -- filter=36 channel=15
    -8, 7, 0, 10, 3, -4, 5, 13, 3,
    -- filter=36 channel=16
    4, -1, 7, 3, 10, 8, -9, 5, 6,
    -- filter=36 channel=17
    6, 14, -8, -16, -10, 10, -1, -12, 11,
    -- filter=36 channel=18
    -3, -12, -13, -7, -14, -9, -5, 13, -4,
    -- filter=36 channel=19
    -13, -14, -5, 0, 14, 2, 11, 5, -10,
    -- filter=36 channel=20
    0, -10, 10, 15, -10, -15, -9, -7, -14,
    -- filter=36 channel=21
    -1, -8, 7, -11, -3, -6, -17, -8, -6,
    -- filter=36 channel=22
    21, 22, 30, 27, 18, 11, 20, -2, 14,
    -- filter=36 channel=23
    5, 6, 11, 17, 1, 14, 13, -11, 10,
    -- filter=36 channel=24
    -5, 11, 0, 13, 4, 4, -6, 9, 12,
    -- filter=36 channel=25
    7, -11, -9, 8, -3, 12, 3, -4, -3,
    -- filter=36 channel=26
    -2, -7, -2, -13, -6, 11, -13, -13, -2,
    -- filter=36 channel=27
    10, -5, 8, -5, -3, 0, 0, -10, 6,
    -- filter=36 channel=28
    10, 15, 3, 0, -10, -8, 11, -8, 0,
    -- filter=36 channel=29
    -5, 9, -5, -6, -8, -7, -3, 19, -4,
    -- filter=36 channel=30
    -10, -9, 7, -11, 9, 0, -1, -11, 1,
    -- filter=36 channel=31
    15, 3, -1, -4, 9, -2, -1, -7, -9,
    -- filter=37 channel=0
    1, 8, 14, 7, 9, 6, 18, 18, 3,
    -- filter=37 channel=1
    -9, -15, 11, -7, 6, 4, 1, 0, -8,
    -- filter=37 channel=2
    13, -4, -1, 4, -14, 9, -2, -5, -12,
    -- filter=37 channel=3
    -5, 5, -4, 3, -7, -6, 5, -5, -14,
    -- filter=37 channel=4
    4, -2, -2, -13, 6, -3, -3, -21, -19,
    -- filter=37 channel=5
    -9, -14, 7, 5, 10, 8, 4, 7, 9,
    -- filter=37 channel=6
    7, -6, 6, -11, -12, 7, -1, -10, -7,
    -- filter=37 channel=7
    -8, -3, -2, 5, 3, 15, -16, 4, -7,
    -- filter=37 channel=8
    -1, 12, 15, 14, 15, -9, 0, 14, -7,
    -- filter=37 channel=9
    -3, -8, 4, 7, -10, 12, 0, 6, 14,
    -- filter=37 channel=10
    -10, 5, -6, 1, 4, 9, 8, 14, -12,
    -- filter=37 channel=11
    11, 20, 20, 22, -3, 20, 12, 4, 7,
    -- filter=37 channel=12
    21, 23, 14, -6, -5, 14, -8, 6, 0,
    -- filter=37 channel=13
    -18, -11, -18, -10, -14, 7, -10, 1, -4,
    -- filter=37 channel=14
    -1, 3, 13, -4, 1, 2, -8, -5, 14,
    -- filter=37 channel=15
    10, 9, 6, -4, 7, 5, -7, -7, 3,
    -- filter=37 channel=16
    -16, -12, -6, -11, 3, -8, -12, -1, -13,
    -- filter=37 channel=17
    0, 7, 10, -20, -7, 13, -20, -10, 0,
    -- filter=37 channel=18
    -20, -4, -1, 8, -17, 4, 1, -4, -15,
    -- filter=37 channel=19
    -10, 10, 10, 0, 0, 14, 1, 0, 14,
    -- filter=37 channel=20
    6, 10, 6, -21, 0, -8, -18, 7, -3,
    -- filter=37 channel=21
    -16, -14, 3, -19, 9, 4, -20, 3, 6,
    -- filter=37 channel=22
    22, 24, 30, 22, 29, 10, 17, 16, 16,
    -- filter=37 channel=23
    -2, -1, 14, 5, 3, -2, 13, 14, -12,
    -- filter=37 channel=24
    3, 9, 2, -12, 9, -11, 7, -6, 12,
    -- filter=37 channel=25
    -4, -4, 4, 7, -13, -9, 8, 10, -6,
    -- filter=37 channel=26
    -17, -14, -13, -15, -8, 2, 4, -11, 10,
    -- filter=37 channel=27
    -1, -6, 0, 2, -6, -1, -9, 9, -6,
    -- filter=37 channel=28
    2, -9, 2, -2, 9, -2, -11, 10, -11,
    -- filter=37 channel=29
    -8, 0, 9, 14, -5, 5, -2, 11, 5,
    -- filter=37 channel=30
    -14, 13, -11, -14, -11, -8, 1, 13, 13,
    -- filter=37 channel=31
    -2, -6, -9, -9, 6, 6, 8, -5, -14,
    -- filter=38 channel=0
    0, 7, -10, -21, 9, -10, -2, -9, 11,
    -- filter=38 channel=1
    -9, -12, -13, -5, 10, 14, 16, 11, -7,
    -- filter=38 channel=2
    13, 0, 10, 9, 7, -14, -4, -7, 5,
    -- filter=38 channel=3
    -14, -10, 0, -4, 4, -7, 4, -4, -6,
    -- filter=38 channel=4
    -1, 7, -3, -11, 2, 3, -13, -5, -9,
    -- filter=38 channel=5
    0, 6, 0, 0, -11, -11, 6, 2, -3,
    -- filter=38 channel=6
    12, 10, 6, 14, -8, 2, 1, -2, -7,
    -- filter=38 channel=7
    -8, 15, 0, -11, 10, -6, 12, -15, -11,
    -- filter=38 channel=8
    -8, -14, -14, -10, 11, -2, 9, -5, 4,
    -- filter=38 channel=9
    3, -9, -16, -10, -8, -7, 0, -3, -9,
    -- filter=38 channel=10
    0, 1, -6, 1, -5, 10, -7, 11, 5,
    -- filter=38 channel=11
    -14, 12, 5, 12, 15, -3, 3, -9, -9,
    -- filter=38 channel=12
    3, -5, 7, 6, 2, -3, -9, -18, 4,
    -- filter=38 channel=13
    18, 11, 17, 6, -6, 14, 7, 16, -8,
    -- filter=38 channel=14
    -5, 0, 13, 10, 2, 8, -1, 4, -7,
    -- filter=38 channel=15
    -6, -14, 4, 1, 9, -7, -9, 10, -8,
    -- filter=38 channel=16
    6, 7, -3, 16, 3, 2, 6, 9, 14,
    -- filter=38 channel=17
    18, 15, -7, 20, 4, 0, 9, -16, 2,
    -- filter=38 channel=18
    -11, 0, -4, 4, 3, 5, 2, -3, -9,
    -- filter=38 channel=19
    14, -11, 0, -8, 8, 7, -9, -10, 12,
    -- filter=38 channel=20
    -2, 14, -4, 8, 5, 0, 3, 0, 13,
    -- filter=38 channel=21
    12, -3, -17, 0, 1, 9, -15, -5, 7,
    -- filter=38 channel=22
    -13, -2, -22, -6, -10, -9, -15, -16, -16,
    -- filter=38 channel=23
    -14, -6, 2, 4, 13, 7, -14, 2, -2,
    -- filter=38 channel=24
    -2, 10, 11, 0, 2, 5, 14, 14, 15,
    -- filter=38 channel=25
    -4, -4, 4, -18, -6, 2, -11, -8, 0,
    -- filter=38 channel=26
    10, 11, -14, 3, -13, -2, 0, -1, -2,
    -- filter=38 channel=27
    -2, 14, 2, -14, 0, 9, -8, -6, -9,
    -- filter=38 channel=28
    13, 8, 3, 5, -6, -11, 2, -3, 8,
    -- filter=38 channel=29
    4, 15, 13, -9, -2, -4, -13, 9, 9,
    -- filter=38 channel=30
    -9, -3, 6, -10, -2, -13, 7, -5, 10,
    -- filter=38 channel=31
    -3, -8, -3, 6, -13, -9, 12, 0, 7,
    -- filter=39 channel=0
    -13, -14, -11, 6, -10, 4, 13, -14, 11,
    -- filter=39 channel=1
    3, 5, -12, 6, 10, -9, -11, -7, 3,
    -- filter=39 channel=2
    -8, -2, 0, -7, 6, -15, -9, 5, -14,
    -- filter=39 channel=3
    2, 11, -11, -7, 13, 4, 13, -9, -12,
    -- filter=39 channel=4
    -4, 0, -2, 5, -6, 11, -5, 5, 0,
    -- filter=39 channel=5
    15, -5, -5, 4, 13, -11, 0, 7, 0,
    -- filter=39 channel=6
    -14, 3, 9, 2, 0, 11, -9, -5, 4,
    -- filter=39 channel=7
    2, 9, -14, 11, 14, -6, 7, -2, 10,
    -- filter=39 channel=8
    -2, -5, 5, -2, 8, 0, -7, 5, 12,
    -- filter=39 channel=9
    -2, 10, -5, 9, -9, 9, -11, 4, -8,
    -- filter=39 channel=10
    -2, -10, 10, -1, -3, -9, -9, -2, -13,
    -- filter=39 channel=11
    2, 11, 1, 10, 16, 1, -4, 1, -10,
    -- filter=39 channel=12
    -13, -9, -10, 1, 14, 4, -9, 9, -10,
    -- filter=39 channel=13
    -12, 11, 1, 13, -4, 15, -3, -3, -13,
    -- filter=39 channel=14
    -7, 0, 9, 15, 5, 13, -8, 11, 3,
    -- filter=39 channel=15
    -4, -12, 4, 0, 11, 2, 6, -6, -5,
    -- filter=39 channel=16
    -3, 9, -4, 7, 4, -3, 12, -10, 6,
    -- filter=39 channel=17
    10, 0, 3, -1, 5, -9, -4, -9, -11,
    -- filter=39 channel=18
    -12, -10, 1, -3, -11, -7, -6, -5, -5,
    -- filter=39 channel=19
    13, -5, -1, -4, 7, -2, 1, 0, 12,
    -- filter=39 channel=20
    2, 9, 7, 17, -12, -10, -7, 9, -8,
    -- filter=39 channel=21
    15, -9, -4, 4, 0, -3, -5, -14, 3,
    -- filter=39 channel=22
    -15, -14, 4, 2, -10, 2, -3, -11, -11,
    -- filter=39 channel=23
    -3, -1, -10, 10, -6, 12, 10, -13, 12,
    -- filter=39 channel=24
    -8, -7, -5, 7, 12, -12, 6, 2, 7,
    -- filter=39 channel=25
    -9, 11, -6, -3, 10, -7, 4, -6, -9,
    -- filter=39 channel=26
    6, 12, 14, 1, 6, 8, -8, 15, -10,
    -- filter=39 channel=27
    7, 0, -4, 1, 12, 12, 1, -9, -3,
    -- filter=39 channel=28
    6, -12, -14, 11, 13, 1, 11, -11, -4,
    -- filter=39 channel=29
    -9, 11, -10, -11, 15, 4, 2, -5, 5,
    -- filter=39 channel=30
    -5, 2, 12, 14, -11, 8, 14, -10, -14,
    -- filter=39 channel=31
    -1, -12, -9, 9, 12, -7, -6, -12, 4,
    -- filter=40 channel=0
    0, 4, 0, 0, -6, 15, 10, 13, -2,
    -- filter=40 channel=1
    9, -10, 0, 4, -15, 3, 0, -12, 1,
    -- filter=40 channel=2
    1, -11, -14, -6, 14, -13, -7, -2, 11,
    -- filter=40 channel=3
    -9, 4, -6, -10, 14, 13, -10, -2, -12,
    -- filter=40 channel=4
    11, 9, 3, -5, -11, -6, 15, 0, 10,
    -- filter=40 channel=5
    10, -13, 8, -4, 9, 10, -11, 12, 4,
    -- filter=40 channel=6
    -4, 13, 9, -7, 2, -8, 4, -9, 1,
    -- filter=40 channel=7
    3, 8, -7, 0, 6, 9, 0, -13, -9,
    -- filter=40 channel=8
    -13, -14, -2, -10, -14, -3, -6, 9, -12,
    -- filter=40 channel=9
    -1, -5, 10, -9, -5, 1, -5, -8, 6,
    -- filter=40 channel=10
    13, 10, 10, 7, 5, 6, 13, 14, -3,
    -- filter=40 channel=11
    -4, -4, 13, -11, 11, -13, -5, -10, -7,
    -- filter=40 channel=12
    -12, 1, 16, -1, 11, 0, -11, 9, -6,
    -- filter=40 channel=13
    2, 5, 13, -4, 1, 9, -14, 10, -15,
    -- filter=40 channel=14
    -15, -2, -5, -8, -5, -2, 6, 2, -4,
    -- filter=40 channel=15
    10, 11, -9, 5, 12, -3, -14, -13, -8,
    -- filter=40 channel=16
    -10, -13, -3, -5, -5, 14, 4, 13, 0,
    -- filter=40 channel=17
    0, -2, 16, -3, -10, -2, -2, 11, -17,
    -- filter=40 channel=18
    -4, -7, 0, -3, -10, -6, -12, 6, 12,
    -- filter=40 channel=19
    0, -12, 4, 1, 10, 1, -13, -8, -5,
    -- filter=40 channel=20
    4, -1, 9, 1, -9, -7, -14, 12, -6,
    -- filter=40 channel=21
    15, 13, 14, -14, 6, 8, -10, 3, -2,
    -- filter=40 channel=22
    5, -1, 14, 9, 19, 5, -6, 13, 12,
    -- filter=40 channel=23
    -9, 7, 10, 15, 12, -10, 14, 0, 8,
    -- filter=40 channel=24
    -6, -2, 3, -14, -11, 2, -10, 13, 3,
    -- filter=40 channel=25
    -10, 10, -7, 0, 7, 5, -4, 6, 12,
    -- filter=40 channel=26
    3, -3, -11, -9, -1, -15, 2, 3, 2,
    -- filter=40 channel=27
    -3, -13, -14, -9, 6, -6, 14, -2, 2,
    -- filter=40 channel=28
    -12, 10, -11, 10, 1, 4, -14, -11, -9,
    -- filter=40 channel=29
    2, 6, 0, -9, -3, 0, -4, -7, 10,
    -- filter=40 channel=30
    -10, 11, -2, -1, -8, 9, 10, 10, -8,
    -- filter=40 channel=31
    -8, -13, -4, 3, 8, -4, -8, -6, -1,
    -- filter=41 channel=0
    10, 0, 2, -1, -8, -15, -10, -11, 11,
    -- filter=41 channel=1
    12, -8, -3, 7, 0, -3, 6, -8, -8,
    -- filter=41 channel=2
    12, -7, 0, -6, 9, -4, 0, 14, -6,
    -- filter=41 channel=3
    -1, 7, -6, -8, 6, 7, 7, -3, 12,
    -- filter=41 channel=4
    8, 9, -8, -16, 1, -8, 13, -7, 1,
    -- filter=41 channel=5
    0, 11, 9, -4, 4, 13, -1, -14, -11,
    -- filter=41 channel=6
    -2, 5, 3, -6, -5, 3, -2, -12, -7,
    -- filter=41 channel=7
    13, -2, -6, 17, -8, -13, -5, 13, 8,
    -- filter=41 channel=8
    -1, 9, 4, -13, -14, 10, 0, -6, -6,
    -- filter=41 channel=9
    3, -8, 11, -12, -14, -9, -11, -5, 0,
    -- filter=41 channel=10
    1, -2, 0, 2, 3, -3, 1, 0, 5,
    -- filter=41 channel=11
    5, -11, -18, 7, 0, -17, -1, 0, -1,
    -- filter=41 channel=12
    0, -12, 3, -15, -11, -3, 6, 12, 5,
    -- filter=41 channel=13
    -3, -20, -7, -18, -12, -18, -17, -4, 3,
    -- filter=41 channel=14
    1, 5, -9, -10, -10, 15, -1, 5, -10,
    -- filter=41 channel=15
    -8, -12, 5, 12, 10, 0, 0, 4, -16,
    -- filter=41 channel=16
    12, 3, 7, -2, 3, 13, 1, 2, -10,
    -- filter=41 channel=17
    12, 3, 0, 20, -1, -15, 19, 13, 1,
    -- filter=41 channel=18
    5, -4, -3, -14, 8, 13, -3, -4, 2,
    -- filter=41 channel=19
    -11, 9, 7, 0, 8, 1, 10, 1, -5,
    -- filter=41 channel=20
    15, 9, 0, -1, 0, 10, 4, 1, -5,
    -- filter=41 channel=21
    14, 0, -12, -4, 0, 5, 12, 9, 1,
    -- filter=41 channel=22
    0, -6, -9, 8, 4, 11, -14, 10, -11,
    -- filter=41 channel=23
    5, -8, 12, -8, 3, -14, 0, 15, 12,
    -- filter=41 channel=24
    -8, -12, 10, -5, -4, -8, 4, 12, 15,
    -- filter=41 channel=25
    -8, 9, 0, -11, 8, 5, -1, 0, -1,
    -- filter=41 channel=26
    -13, 4, 0, 3, -3, -15, -5, -10, -19,
    -- filter=41 channel=27
    7, -12, 1, 7, 13, 9, 11, 2, 14,
    -- filter=41 channel=28
    14, -13, 9, -7, 3, 4, 9, -10, -5,
    -- filter=41 channel=29
    -1, -10, -1, -1, -6, -18, -17, 5, 8,
    -- filter=41 channel=30
    3, -4, 0, 8, 0, 4, -6, -3, -10,
    -- filter=41 channel=31
    4, -15, 3, 0, -7, -9, -6, 2, 9,
    -- filter=42 channel=0
    15, 8, 1, 12, -7, -6, 1, -9, -10,
    -- filter=42 channel=1
    9, -3, 6, -6, 8, 3, 12, 11, 15,
    -- filter=42 channel=2
    -8, -8, 0, 12, -9, 0, -9, 14, 4,
    -- filter=42 channel=3
    -7, -14, 1, 11, -13, 10, -9, -3, 11,
    -- filter=42 channel=4
    2, -1, 14, 6, 14, 8, 12, 10, 15,
    -- filter=42 channel=5
    6, -12, 10, 0, -10, -2, -9, -3, 2,
    -- filter=42 channel=6
    5, -7, -2, 14, -10, 8, -8, 0, -5,
    -- filter=42 channel=7
    -12, -11, -6, -12, -15, 5, 21, 8, 0,
    -- filter=42 channel=8
    12, -3, -5, 10, -5, 2, 3, 0, 6,
    -- filter=42 channel=9
    1, -2, 4, 2, -5, -6, 2, 9, 0,
    -- filter=42 channel=10
    3, -11, -5, 0, 8, 13, 4, -8, -3,
    -- filter=42 channel=11
    5, 3, -8, 6, -15, -16, 10, 0, 2,
    -- filter=42 channel=12
    -8, -13, 2, -17, -17, 7, -6, 12, 8,
    -- filter=42 channel=13
    -2, 8, -8, 5, 5, -5, 0, -3, 0,
    -- filter=42 channel=14
    8, 0, 15, -8, -8, -10, 11, 3, -9,
    -- filter=42 channel=15
    8, -13, -4, 11, -10, 12, 4, 6, -5,
    -- filter=42 channel=16
    8, -7, -4, 5, -9, -12, -9, 6, -12,
    -- filter=42 channel=17
    9, 8, -8, -1, 3, 3, 14, 12, 14,
    -- filter=42 channel=18
    14, 0, 0, -1, -3, -6, -5, 13, 2,
    -- filter=42 channel=19
    -2, 3, -6, -10, 10, 2, 11, -13, -4,
    -- filter=42 channel=20
    -19, -15, -18, -12, 10, -19, 13, -3, -9,
    -- filter=42 channel=21
    2, -8, -1, 11, -3, 5, -2, 6, 15,
    -- filter=42 channel=22
    0, 6, -15, -12, 2, -8, 6, -16, -10,
    -- filter=42 channel=23
    -8, -13, 9, -9, -6, -8, -7, 1, -10,
    -- filter=42 channel=24
    -14, -5, -1, 10, -10, -6, -9, 2, -7,
    -- filter=42 channel=25
    -8, 7, 12, -5, -4, 3, -11, -3, 0,
    -- filter=42 channel=26
    1, 0, -14, 2, 0, 13, 12, -4, 0,
    -- filter=42 channel=27
    -5, 11, 9, -11, -13, -8, 8, 13, -2,
    -- filter=42 channel=28
    2, -14, 2, -9, -9, 11, 17, -7, -12,
    -- filter=42 channel=29
    14, -1, 13, -14, 8, 12, 13, -7, 8,
    -- filter=42 channel=30
    -11, -6, -6, 11, 13, -1, -7, 2, 14,
    -- filter=42 channel=31
    1, -2, 6, -10, 13, -15, 8, 7, 1,
    -- filter=43 channel=0
    -3, -3, 5, -2, -11, -3, -6, -9, -6,
    -- filter=43 channel=1
    6, -10, -17, -2, 9, -13, -12, 7, -2,
    -- filter=43 channel=2
    -2, -2, 6, -12, -1, 0, -14, 0, -7,
    -- filter=43 channel=3
    0, 5, -2, -6, -15, -6, 3, 0, 4,
    -- filter=43 channel=4
    14, 6, 0, -4, 13, 5, 7, 5, 2,
    -- filter=43 channel=5
    11, -1, 4, -17, 9, -4, -3, -16, -4,
    -- filter=43 channel=6
    -5, 7, 5, -5, -14, 5, -9, -7, 11,
    -- filter=43 channel=7
    0, 0, -5, 10, -2, -8, 2, 7, -22,
    -- filter=43 channel=8
    0, -14, -10, -8, -13, 4, -16, -13, 14,
    -- filter=43 channel=9
    9, -5, 14, -16, 6, 1, 2, -4, -5,
    -- filter=43 channel=10
    0, 1, -15, -15, -19, 4, -19, 3, 2,
    -- filter=43 channel=11
    18, -3, 18, 0, 15, 9, -1, -4, -4,
    -- filter=43 channel=12
    -2, 15, -11, -5, -15, -13, -2, -12, 5,
    -- filter=43 channel=13
    3, -20, -9, 0, -15, -16, -10, -6, -10,
    -- filter=43 channel=14
    0, 9, 12, 7, 3, 0, 20, -5, 15,
    -- filter=43 channel=15
    -3, -16, 8, -18, -14, -13, -9, -19, -15,
    -- filter=43 channel=16
    17, -7, 0, 5, 10, 8, -2, -11, -11,
    -- filter=43 channel=17
    0, 4, -6, -8, -12, -10, -7, -16, -24,
    -- filter=43 channel=18
    9, 5, 13, 13, 3, -3, 2, -6, 7,
    -- filter=43 channel=19
    11, 10, 5, -14, 12, 0, 7, -10, 7,
    -- filter=43 channel=20
    33, 23, 5, 0, 6, 6, 6, 15, 3,
    -- filter=43 channel=21
    4, -20, -3, -12, -19, -10, 2, 2, -19,
    -- filter=43 channel=22
    2, 8, 13, 2, 7, 1, -17, 3, -11,
    -- filter=43 channel=23
    3, 18, 3, 0, 15, 13, 4, 12, -11,
    -- filter=43 channel=24
    22, 1, 3, 17, 0, 11, 5, 21, 9,
    -- filter=43 channel=25
    -15, 3, -13, -15, -5, -6, -2, 4, 15,
    -- filter=43 channel=26
    -25, -21, -16, -12, -15, -25, -12, -2, -18,
    -- filter=43 channel=27
    8, 8, -5, -1, 4, -11, 2, 10, -8,
    -- filter=43 channel=28
    13, 9, -2, 0, -5, -1, 15, 4, -4,
    -- filter=43 channel=29
    4, 5, 17, -6, 0, 21, 17, -1, 18,
    -- filter=43 channel=30
    -11, 3, 11, -13, -12, 12, 2, 1, -9,
    -- filter=43 channel=31
    -12, -10, -12, 0, 1, -10, 2, -18, -2,
    -- filter=44 channel=0
    -16, -3, -15, 2, 9, -9, 7, -12, -11,
    -- filter=44 channel=1
    0, -2, -5, 13, 8, 4, 8, 12, 11,
    -- filter=44 channel=2
    1, 8, -8, 7, -12, 5, 10, -9, -6,
    -- filter=44 channel=3
    -7, -1, 6, 13, 2, 7, 5, -2, 6,
    -- filter=44 channel=4
    -2, 4, -2, -7, -7, -7, 16, -6, 15,
    -- filter=44 channel=5
    -1, -8, 12, 12, 12, 1, 0, -10, -16,
    -- filter=44 channel=6
    7, 10, 9, 0, -4, -2, -2, 6, 2,
    -- filter=44 channel=7
    -3, -10, 12, 8, -7, -15, 8, -1, 0,
    -- filter=44 channel=8
    -7, 0, 5, -9, 3, -1, -9, -14, -10,
    -- filter=44 channel=9
    -15, 9, -15, 13, -12, 10, 0, -14, 9,
    -- filter=44 channel=10
    -13, -18, 4, -9, -1, 8, -10, -2, -6,
    -- filter=44 channel=11
    3, -11, 11, 12, -5, -1, -1, -14, -3,
    -- filter=44 channel=12
    1, 9, 0, -12, -16, -17, 0, 2, -5,
    -- filter=44 channel=13
    5, -12, -17, 5, -20, 1, -4, -8, -20,
    -- filter=44 channel=14
    9, 8, -12, 14, 10, -1, -8, 4, 10,
    -- filter=44 channel=15
    6, -3, -18, 0, -16, -7, -13, -6, 0,
    -- filter=44 channel=16
    -14, -11, -6, -6, 7, 0, 3, 0, 5,
    -- filter=44 channel=17
    3, -5, 9, 6, 9, -5, -1, -1, -1,
    -- filter=44 channel=18
    -4, -8, 9, 8, -1, 14, -5, 0, 0,
    -- filter=44 channel=19
    2, 9, -11, -14, 7, -14, 13, 0, 7,
    -- filter=44 channel=20
    5, 5, -2, -4, 0, 0, -4, 8, 2,
    -- filter=44 channel=21
    -3, 7, 1, 11, 9, -1, 10, -5, 11,
    -- filter=44 channel=22
    6, -16, -15, 2, 5, -15, 2, 1, 4,
    -- filter=44 channel=23
    8, -9, 6, 11, 16, 10, 7, -8, 8,
    -- filter=44 channel=24
    -14, 13, 11, 10, 0, -4, -5, -1, -12,
    -- filter=44 channel=25
    15, 10, 14, -10, 8, 13, 17, 18, 10,
    -- filter=44 channel=26
    -3, -3, -4, -12, 1, -4, -3, -10, 0,
    -- filter=44 channel=27
    13, 12, -3, -11, -4, -10, 12, 8, 12,
    -- filter=44 channel=28
    11, 6, 1, -11, 11, -7, -2, -9, -9,
    -- filter=44 channel=29
    9, -15, 1, -12, 6, -2, -16, -2, 0,
    -- filter=44 channel=30
    2, 0, 12, -13, 5, -12, 12, -3, -5,
    -- filter=44 channel=31
    0, -14, -12, 2, -8, -17, -5, 0, -17,
    -- filter=45 channel=0
    -24, -22, -9, -23, -6, -1, 0, -19, 1,
    -- filter=45 channel=1
    6, -21, -3, -7, -4, 0, -7, -10, -23,
    -- filter=45 channel=2
    2, -6, -9, 8, 13, 8, 2, -4, -8,
    -- filter=45 channel=3
    3, 9, -6, 2, -8, 10, -13, 11, 8,
    -- filter=45 channel=4
    10, 13, -1, 5, 12, -2, 5, 0, -3,
    -- filter=45 channel=5
    6, 21, 0, -4, 3, -7, 7, 19, -3,
    -- filter=45 channel=6
    7, 6, 6, 8, -11, 14, -5, -2, 10,
    -- filter=45 channel=7
    16, -20, -31, 20, -16, -32, 26, 0, -27,
    -- filter=45 channel=8
    15, 9, 14, 17, 9, 0, 14, 0, 11,
    -- filter=45 channel=9
    -3, 5, -2, 8, 1, -7, 7, -7, -10,
    -- filter=45 channel=10
    8, 15, 0, 6, 17, -3, 0, 12, 5,
    -- filter=45 channel=11
    -7, -7, 1, 1, 8, 9, -2, 0, -6,
    -- filter=45 channel=12
    11, -17, -24, -10, 0, -5, 12, -10, -16,
    -- filter=45 channel=13
    -4, 1, -21, 2, -21, -26, 13, 2, -26,
    -- filter=45 channel=14
    -4, -16, -15, -20, -17, -4, -23, -5, -10,
    -- filter=45 channel=15
    14, 4, -9, 6, -3, -14, 23, 1, -12,
    -- filter=45 channel=16
    13, -8, 6, 0, 10, 8, 4, 13, 2,
    -- filter=45 channel=17
    25, 17, -33, 44, 0, -21, 48, 13, -8,
    -- filter=45 channel=18
    -7, 7, -11, 5, 6, -1, -7, 6, 13,
    -- filter=45 channel=19
    9, -13, 4, -1, 10, -7, 11, 10, -13,
    -- filter=45 channel=20
    2, -19, -22, 15, -21, -34, 13, 0, -32,
    -- filter=45 channel=21
    36, 1, -33, 43, 5, -31, 40, 19, -20,
    -- filter=45 channel=22
    -3, 24, 1, 17, 19, -4, 19, -4, -1,
    -- filter=45 channel=23
    5, 13, -5, 6, 9, -11, -8, 17, 5,
    -- filter=45 channel=24
    -5, -20, -16, 1, -16, 2, 12, -2, -10,
    -- filter=45 channel=25
    17, -5, -5, 16, -14, 0, -7, 4, -6,
    -- filter=45 channel=26
    29, 7, 3, 28, 13, -6, 35, 1, 4,
    -- filter=45 channel=27
    12, 7, 13, -11, -9, 10, 0, -9, -14,
    -- filter=45 channel=28
    0, 8, -9, -1, -7, -7, 9, 2, 13,
    -- filter=45 channel=29
    8, 9, 27, 13, 23, 17, 6, 12, 24,
    -- filter=45 channel=30
    -3, 12, -3, 0, 6, 1, 5, -4, 8,
    -- filter=45 channel=31
    13, 3, -10, 5, 11, 3, 15, -15, -11,
    -- filter=46 channel=0
    -12, 12, -6, -3, 9, 7, -4, 7, -1,
    -- filter=46 channel=1
    11, 0, -3, 11, -12, -13, 8, -16, -11,
    -- filter=46 channel=2
    11, -2, 2, -3, -10, 0, -6, 15, 9,
    -- filter=46 channel=3
    13, 7, 1, 4, -3, 1, -2, 0, -13,
    -- filter=46 channel=4
    12, 8, 0, -2, 0, -16, -14, 0, -15,
    -- filter=46 channel=5
    0, 15, 14, -11, -1, 12, -2, 0, -16,
    -- filter=46 channel=6
    4, 11, -12, 2, 4, 14, -4, 3, -7,
    -- filter=46 channel=7
    14, 16, -7, -10, -9, 13, -1, -16, -4,
    -- filter=46 channel=8
    -5, 9, 0, 8, 11, 6, 2, -1, -13,
    -- filter=46 channel=9
    1, 0, -3, 15, 17, -5, -5, -7, 3,
    -- filter=46 channel=10
    6, 11, 3, 9, 2, 0, 0, 0, -11,
    -- filter=46 channel=11
    6, -8, -4, 19, -9, 7, 0, 16, 5,
    -- filter=46 channel=12
    2, 13, 17, 17, 0, 7, 2, -10, 11,
    -- filter=46 channel=13
    3, -11, 5, 11, -4, -12, -10, -13, -10,
    -- filter=46 channel=14
    -4, -13, -15, 10, -12, -8, 13, -2, -10,
    -- filter=46 channel=15
    -9, -4, 2, 1, 14, -8, -9, 2, 10,
    -- filter=46 channel=16
    14, 0, 0, -7, -11, 0, -4, -10, -1,
    -- filter=46 channel=17
    8, 18, 16, -11, 6, -8, -9, -11, -20,
    -- filter=46 channel=18
    -14, 0, -13, -14, -2, -14, -2, 13, -5,
    -- filter=46 channel=19
    6, 14, -12, -1, -3, -2, 5, 5, 3,
    -- filter=46 channel=20
    -2, 16, 10, -9, 7, -1, -9, 6, -12,
    -- filter=46 channel=21
    7, 0, -6, 8, 4, -10, -13, -5, -8,
    -- filter=46 channel=22
    -1, 11, 6, 13, 26, 15, 28, 22, 25,
    -- filter=46 channel=23
    7, 12, 11, 14, 0, -9, 18, -8, 15,
    -- filter=46 channel=24
    -10, -15, 6, -8, -11, -8, -1, -1, -14,
    -- filter=46 channel=25
    0, -1, -3, 2, -12, -6, 12, -8, 13,
    -- filter=46 channel=26
    13, 6, 9, 4, -7, -9, -7, -17, -10,
    -- filter=46 channel=27
    0, 6, -6, -5, 3, 1, 3, -4, 5,
    -- filter=46 channel=28
    -12, 1, 2, 13, -14, 12, -3, -10, 13,
    -- filter=46 channel=29
    12, -6, 9, 14, 1, -6, -6, 15, -9,
    -- filter=46 channel=30
    -4, -2, -12, 9, -11, -14, -14, 10, -2,
    -- filter=46 channel=31
    11, -8, 3, 9, -12, -2, -9, -8, 11,
    -- filter=47 channel=0
    13, 13, 8, -2, 13, 14, 5, 1, -3,
    -- filter=47 channel=1
    1, -16, 3, -6, 1, -13, -14, 11, 14,
    -- filter=47 channel=2
    9, 0, -14, 11, -6, -15, 2, 0, 1,
    -- filter=47 channel=3
    9, -1, -10, 14, -1, 0, -5, 2, 13,
    -- filter=47 channel=4
    -10, 15, 12, 0, 15, -4, 17, 13, 13,
    -- filter=47 channel=5
    13, -9, 3, -1, -4, -2, -13, 7, 4,
    -- filter=47 channel=6
    -6, -5, -6, 8, -8, -12, -6, 9, 3,
    -- filter=47 channel=7
    4, -18, -15, -2, -18, -5, -13, 11, -2,
    -- filter=47 channel=8
    0, 8, 13, 14, 2, 8, -1, -7, 0,
    -- filter=47 channel=9
    -9, 0, -12, -1, -12, 8, -4, -6, 0,
    -- filter=47 channel=10
    10, 4, 6, 8, 7, 14, 7, 2, 9,
    -- filter=47 channel=11
    -7, -6, -10, 1, -11, -4, -22, -5, -11,
    -- filter=47 channel=12
    -12, -2, 6, 2, 11, 0, -1, -16, 0,
    -- filter=47 channel=13
    -9, 3, -3, 14, 2, 12, -11, -6, -8,
    -- filter=47 channel=14
    9, -12, -5, 2, 0, 13, -3, 0, 10,
    -- filter=47 channel=15
    7, -10, -9, -6, -6, -6, -1, -8, 6,
    -- filter=47 channel=16
    3, 5, -15, 1, 6, -12, -13, -14, -4,
    -- filter=47 channel=17
    14, -3, -8, 3, -13, 11, 8, 0, -16,
    -- filter=47 channel=18
    14, -1, 0, 6, 16, 7, 9, -2, 4,
    -- filter=47 channel=19
    -5, -3, -8, 12, -8, 13, 13, 11, -11,
    -- filter=47 channel=20
    -3, 8, -9, -13, -13, -2, -12, -1, 7,
    -- filter=47 channel=21
    -1, -5, -12, -2, 1, -9, 8, -3, 3,
    -- filter=47 channel=22
    -1, 0, -13, -10, 13, -5, -11, -13, 5,
    -- filter=47 channel=23
    3, -7, 1, -4, 16, 13, 11, -8, 15,
    -- filter=47 channel=24
    7, -7, 8, -13, -12, -8, 10, 12, 6,
    -- filter=47 channel=25
    21, 13, 4, 11, 24, 21, 21, 4, 17,
    -- filter=47 channel=26
    -10, 11, -6, 10, -3, -14, 8, -10, -15,
    -- filter=47 channel=27
    5, 10, 11, 3, 8, -11, 5, -11, -10,
    -- filter=47 channel=28
    1, 12, 7, -11, -3, -5, 12, -2, -6,
    -- filter=47 channel=29
    4, 0, -5, 0, -20, -15, 1, -19, -17,
    -- filter=47 channel=30
    5, 3, -6, 14, -10, 3, 0, 0, 0,
    -- filter=47 channel=31
    0, 8, 13, -3, -8, 5, 10, -8, -5,
    -- filter=48 channel=0
    13, 18, 7, 11, -6, 5, 1, 8, 2,
    -- filter=48 channel=1
    11, -4, 22, 7, -6, 18, 10, 7, 18,
    -- filter=48 channel=2
    -4, 4, -2, 8, -5, 15, 12, -5, -3,
    -- filter=48 channel=3
    11, 3, -14, 12, 9, -2, 0, 3, -6,
    -- filter=48 channel=4
    -7, -4, 9, -18, 4, 2, -11, -11, 13,
    -- filter=48 channel=5
    -11, 2, -4, -8, 5, -5, -5, 6, 0,
    -- filter=48 channel=6
    -1, 8, 13, 0, 3, -14, 4, 5, -10,
    -- filter=48 channel=7
    -9, 9, 26, -17, 0, 23, -10, -10, 20,
    -- filter=48 channel=8
    0, -10, -10, 14, 2, -16, 8, 10, 3,
    -- filter=48 channel=9
    -9, 4, -12, -4, -14, 5, 7, 4, -2,
    -- filter=48 channel=10
    -4, 13, 6, -9, 9, 2, 1, -6, 16,
    -- filter=48 channel=11
    -10, -19, -10, 0, -5, -12, 0, 9, 2,
    -- filter=48 channel=12
    6, -1, 6, 0, -4, 3, 4, -13, 17,
    -- filter=48 channel=13
    7, 5, 20, 7, -11, 17, 1, 9, 7,
    -- filter=48 channel=14
    -5, 1, 2, 11, -5, 12, -11, -7, 18,
    -- filter=48 channel=15
    0, 8, 3, -3, 1, -4, -16, -1, -15,
    -- filter=48 channel=16
    -4, 12, 7, -14, -11, 0, -15, -11, -7,
    -- filter=48 channel=17
    -9, -2, 7, -2, -7, 14, -3, -17, 0,
    -- filter=48 channel=18
    -15, 0, -3, -9, -6, 11, -3, 12, 6,
    -- filter=48 channel=19
    2, -1, -12, 2, 8, -6, -6, 13, 5,
    -- filter=48 channel=20
    -6, 5, 24, -27, 1, 21, -17, -2, 5,
    -- filter=48 channel=21
    -16, 16, 15, -9, -8, 25, 1, 12, 11,
    -- filter=48 channel=22
    3, -7, -20, -15, -3, -10, -9, -17, 5,
    -- filter=48 channel=23
    -13, 9, 11, 10, -2, -13, -12, -8, -8,
    -- filter=48 channel=24
    -3, 4, 1, 5, 12, 1, -15, 9, -12,
    -- filter=48 channel=25
    -9, -1, 9, -9, 7, 8, -15, -6, 14,
    -- filter=48 channel=26
    0, -18, 0, -6, -16, 2, -1, 0, 5,
    -- filter=48 channel=27
    -4, 10, -4, 0, -11, 13, 13, 1, 4,
    -- filter=48 channel=28
    8, -12, 5, -11, 12, -14, -5, 1, -9,
    -- filter=48 channel=29
    2, -2, -8, -15, 0, -11, -8, -20, -12,
    -- filter=48 channel=30
    -10, -10, 7, 1, -14, -4, -2, -5, 9,
    -- filter=48 channel=31
    -5, 14, 11, -17, -16, 6, 11, -1, 9,
    -- filter=49 channel=0
    12, 7, 7, 12, -9, -2, -7, 1, -5,
    -- filter=49 channel=1
    -5, 6, 9, -15, -5, 0, 1, 4, 6,
    -- filter=49 channel=2
    -10, -5, 10, -5, 5, 3, 0, 3, 1,
    -- filter=49 channel=3
    -13, 10, 14, -10, 12, 7, -10, -1, 11,
    -- filter=49 channel=4
    11, -10, 10, -3, -1, 6, -13, -7, 3,
    -- filter=49 channel=5
    -11, -10, 10, 7, -6, 5, 14, 2, -2,
    -- filter=49 channel=6
    -13, -1, 8, 2, 0, 1, 11, 0, 15,
    -- filter=49 channel=7
    -13, -4, 9, 1, 12, 2, -10, 5, 8,
    -- filter=49 channel=8
    -8, 13, 10, 6, 4, -6, -4, 9, -10,
    -- filter=49 channel=9
    0, 13, -13, 12, 2, 12, -4, 1, -2,
    -- filter=49 channel=10
    -14, 13, 13, 4, 0, -14, 10, 4, -13,
    -- filter=49 channel=11
    -11, 4, -9, -8, 6, 12, -9, -11, 8,
    -- filter=49 channel=12
    -2, 1, 11, 3, -10, -6, 3, -2, -12,
    -- filter=49 channel=13
    17, 4, 8, 7, -8, 12, 13, -12, -9,
    -- filter=49 channel=14
    0, -12, 0, 13, -1, 9, 2, 14, -12,
    -- filter=49 channel=15
    13, 15, -12, 12, 0, -13, -5, -12, 0,
    -- filter=49 channel=16
    0, 8, -11, 4, 4, 7, 10, -3, -4,
    -- filter=49 channel=17
    9, -1, -3, 10, 6, -12, -8, 9, -10,
    -- filter=49 channel=18
    -13, -4, 9, 11, -2, 4, -3, -3, -13,
    -- filter=49 channel=19
    0, 1, 12, 6, 11, 5, -11, 12, -5,
    -- filter=49 channel=20
    -8, -2, 5, -7, -1, -5, 4, -10, -2,
    -- filter=49 channel=21
    -3, -4, -8, -15, -14, -7, -13, -12, -9,
    -- filter=49 channel=22
    8, -9, -8, 2, 9, -6, -2, -6, -12,
    -- filter=49 channel=23
    9, -14, -5, 2, 1, -11, 14, 8, 13,
    -- filter=49 channel=24
    -1, 13, -11, -5, 11, -5, -4, -5, 1,
    -- filter=49 channel=25
    9, 6, -11, 6, 5, -2, -5, 7, -3,
    -- filter=49 channel=26
    -6, 15, 10, 7, -7, 13, 9, 8, -4,
    -- filter=49 channel=27
    1, -8, -11, 1, 11, -5, -7, 2, -15,
    -- filter=49 channel=28
    6, 3, 10, 13, -6, -3, -15, 13, -5,
    -- filter=49 channel=29
    -8, 10, -14, 1, 3, -10, -7, 2, 0,
    -- filter=49 channel=30
    -3, -9, 13, -9, 6, -11, 8, 11, -13,
    -- filter=49 channel=31
    8, -1, 1, -7, 1, 15, 0, 1, 10,
    -- filter=50 channel=0
    -9, 2, -12, -5, 10, -14, -11, 4, -9,
    -- filter=50 channel=1
    -9, 10, 7, 13, -10, 11, 10, 5, -8,
    -- filter=50 channel=2
    1, -13, 4, -11, -3, -3, -7, -5, -4,
    -- filter=50 channel=3
    12, -5, -3, 10, 6, 13, -5, -13, -7,
    -- filter=50 channel=4
    2, 11, 3, -11, -15, 10, -5, 7, 3,
    -- filter=50 channel=5
    7, 10, -5, -2, 9, 15, 10, -14, 8,
    -- filter=50 channel=6
    -14, 3, 0, -7, 5, 4, -6, 14, 13,
    -- filter=50 channel=7
    -2, 5, 16, -8, -11, 0, -12, 8, 14,
    -- filter=50 channel=8
    -11, 0, -13, -9, -9, -9, 3, -10, 5,
    -- filter=50 channel=9
    12, 0, 13, 1, 0, 0, 13, 3, 14,
    -- filter=50 channel=10
    -14, -10, -2, -6, 4, 14, 1, -4, -8,
    -- filter=50 channel=11
    -14, -19, -19, -8, -2, -8, -5, 5, -19,
    -- filter=50 channel=12
    1, 8, 4, -11, 15, -5, -6, 11, -2,
    -- filter=50 channel=13
    -9, -14, 1, -19, 3, 15, 9, -3, 0,
    -- filter=50 channel=14
    -15, 8, 4, -12, 7, 3, -3, -4, -5,
    -- filter=50 channel=15
    -5, -5, 7, 0, -7, 0, -10, 3, -9,
    -- filter=50 channel=16
    6, -7, 9, 8, -13, -5, 2, -5, -9,
    -- filter=50 channel=17
    -14, -7, 6, 10, -3, 3, 2, 16, 18,
    -- filter=50 channel=18
    3, 13, 0, 10, -7, 4, 11, -14, -3,
    -- filter=50 channel=19
    3, -10, 9, 10, -2, -5, -11, -5, -5,
    -- filter=50 channel=20
    -8, 4, 18, -10, 1, 8, -7, -7, 4,
    -- filter=50 channel=21
    -12, 9, 6, 8, 10, -8, 6, 6, 18,
    -- filter=50 channel=22
    0, -4, -13, -13, 5, 0, 1, 2, 1,
    -- filter=50 channel=23
    -8, -8, 11, -5, 0, 5, -12, 3, 10,
    -- filter=50 channel=24
    0, 8, -8, -7, 7, -10, -1, -12, -14,
    -- filter=50 channel=25
    3, -1, -6, -2, -1, 1, 1, 2, -12,
    -- filter=50 channel=26
    -15, -6, -5, -15, 0, -13, -8, -1, -4,
    -- filter=50 channel=27
    -8, 10, 8, 6, -2, -3, 10, 0, 0,
    -- filter=50 channel=28
    7, 4, -1, -7, -1, 9, 0, 10, 7,
    -- filter=50 channel=29
    0, 1, -11, -16, -17, -12, -13, 8, -6,
    -- filter=50 channel=30
    8, 2, 1, 1, 1, -1, -14, -7, -12,
    -- filter=50 channel=31
    -5, 10, 17, 10, 4, -10, -1, 4, 17,
    -- filter=51 channel=0
    14, -1, 12, 11, -9, 1, -12, 13, -12,
    -- filter=51 channel=1
    -8, -16, 7, -3, 4, 1, 9, -13, 0,
    -- filter=51 channel=2
    -6, 13, -11, -2, 12, -5, -13, -1, 2,
    -- filter=51 channel=3
    14, 4, 4, 5, -15, 12, 11, 12, -9,
    -- filter=51 channel=4
    14, 6, 16, -4, 16, 11, 19, 3, 11,
    -- filter=51 channel=5
    1, -1, 0, -3, 7, 1, 8, -16, 10,
    -- filter=51 channel=6
    0, -2, 9, 3, 2, 1, 3, 8, 5,
    -- filter=51 channel=7
    -7, -24, -19, -15, -3, -24, -22, -8, -7,
    -- filter=51 channel=8
    -1, 13, 10, 6, 0, 1, 0, 14, 10,
    -- filter=51 channel=9
    12, -7, 2, 9, -7, 3, 11, -13, -1,
    -- filter=51 channel=10
    -19, -5, -5, -10, -1, -6, -10, -11, 9,
    -- filter=51 channel=11
    7, -1, -5, 6, -2, 4, 7, -8, 6,
    -- filter=51 channel=12
    -4, 3, -9, -5, -20, -11, -20, -9, -2,
    -- filter=51 channel=13
    -16, 0, -26, -6, -11, -21, -26, -3, -27,
    -- filter=51 channel=14
    4, 1, 10, 16, 24, 23, 7, 18, 14,
    -- filter=51 channel=15
    -7, -9, -13, -12, -2, -3, -13, 9, 6,
    -- filter=51 channel=16
    5, 13, 11, 2, -8, 1, -4, -12, 3,
    -- filter=51 channel=17
    -10, -23, -25, -30, 0, -16, -11, -9, -8,
    -- filter=51 channel=18
    -4, -2, 3, -6, 17, 16, 16, 21, 19,
    -- filter=51 channel=19
    11, 10, 6, 10, 5, 3, -6, 8, 14,
    -- filter=51 channel=20
    -20, -10, -7, -20, -9, -22, -3, -5, -16,
    -- filter=51 channel=21
    -9, -9, -10, -6, -13, -15, -13, 6, -12,
    -- filter=51 channel=22
    -8, -9, 5, 0, -16, 0, 4, 6, 4,
    -- filter=51 channel=23
    0, 8, 3, 11, -8, 14, 3, 5, -3,
    -- filter=51 channel=24
    16, 1, 7, -5, 14, 6, 19, 9, 18,
    -- filter=51 channel=25
    14, 16, 22, 8, 17, 1, 16, 10, 20,
    -- filter=51 channel=26
    -4, -4, -15, -5, -3, -3, -10, -8, -8,
    -- filter=51 channel=27
    -10, 14, 9, 10, 0, 5, 3, 2, 12,
    -- filter=51 channel=28
    1, -8, -13, -6, -16, -12, -4, 5, 6,
    -- filter=51 channel=29
    3, -10, -9, 10, 7, -13, -5, 13, -4,
    -- filter=51 channel=30
    -12, -13, -6, 1, -4, -6, 1, 8, -5,
    -- filter=51 channel=31
    4, -19, 8, -4, -16, 6, -20, -10, 2,
    -- filter=52 channel=0
    4, 9, -8, -13, -15, -10, -8, 11, -10,
    -- filter=52 channel=1
    10, 11, 11, 7, 8, 8, -4, 15, 16,
    -- filter=52 channel=2
    1, -8, 4, 0, -9, 14, 12, -11, 2,
    -- filter=52 channel=3
    -13, 14, -3, 9, 6, -11, -13, 12, -5,
    -- filter=52 channel=4
    -1, 9, 15, 5, -12, 10, -6, 5, -3,
    -- filter=52 channel=5
    7, 4, -5, 2, -7, -12, 0, -1, -5,
    -- filter=52 channel=6
    -11, 7, 6, 0, -3, -1, -3, -6, 3,
    -- filter=52 channel=7
    -13, 8, 10, -6, -12, 13, -2, 10, -13,
    -- filter=52 channel=8
    -13, -6, 10, -1, 10, 7, -7, 0, 7,
    -- filter=52 channel=9
    -5, -14, -9, -6, -12, 12, -5, 5, 7,
    -- filter=52 channel=10
    0, 7, -5, -1, 6, 12, -3, 3, -12,
    -- filter=52 channel=11
    -4, -16, 2, -14, -12, 8, -8, 9, -9,
    -- filter=52 channel=12
    7, 8, -16, 1, -8, 10, -3, -11, -7,
    -- filter=52 channel=13
    -8, 0, 0, 2, 1, -16, -6, 7, -11,
    -- filter=52 channel=14
    -10, -11, 6, 2, 1, 14, 13, 1, 0,
    -- filter=52 channel=15
    0, -8, -5, -13, -9, -11, 12, 8, 12,
    -- filter=52 channel=16
    -9, 7, -4, 13, 14, -6, -2, 1, 11,
    -- filter=52 channel=17
    -6, -11, 16, -16, 3, -5, -12, 1, -15,
    -- filter=52 channel=18
    0, 0, -6, -5, 15, -7, 3, -3, 16,
    -- filter=52 channel=19
    -1, 7, 10, -10, -9, -10, -12, 14, -7,
    -- filter=52 channel=20
    2, 12, 22, -5, 11, 3, -11, -9, 17,
    -- filter=52 channel=21
    1, 4, 12, -18, -1, 4, -10, 3, 4,
    -- filter=52 channel=22
    -16, 0, -17, -16, 5, -15, -2, -18, -21,
    -- filter=52 channel=23
    -13, 1, -1, -13, 12, -15, -7, -16, 7,
    -- filter=52 channel=24
    16, -10, 9, -12, -9, 7, 1, -10, 14,
    -- filter=52 channel=25
    -6, 2, 0, 5, 12, 15, -8, 8, -7,
    -- filter=52 channel=26
    -16, 12, -11, 0, 3, -11, -1, 11, -14,
    -- filter=52 channel=27
    -11, -9, -8, -1, -13, 9, -12, -5, 5,
    -- filter=52 channel=28
    -7, -2, 2, -16, 6, -8, -10, 0, 5,
    -- filter=52 channel=29
    0, 3, -5, 7, 11, 6, -9, 2, -11,
    -- filter=52 channel=30
    -4, -1, 7, 15, 9, -4, -14, -12, 6,
    -- filter=52 channel=31
    -4, -6, -15, -15, -11, -3, -1, -7, -11,
    -- filter=53 channel=0
    -5, 13, 4, -6, -10, 13, -7, -7, 7,
    -- filter=53 channel=1
    6, -15, -9, -8, 6, 10, 7, 0, 3,
    -- filter=53 channel=2
    -1, 8, 0, 12, 11, 8, 0, -10, 5,
    -- filter=53 channel=3
    14, 0, -11, -11, 9, 11, 1, 12, -1,
    -- filter=53 channel=4
    -9, 10, -15, -9, 0, 12, 5, -12, -13,
    -- filter=53 channel=5
    0, 12, 7, -1, -4, 8, 5, -5, 10,
    -- filter=53 channel=6
    5, 0, 13, -10, -2, -8, 14, -7, 0,
    -- filter=53 channel=7
    11, -11, -5, 0, -12, -14, 10, 8, 0,
    -- filter=53 channel=8
    -11, 3, 6, -11, 10, 7, 5, -10, 2,
    -- filter=53 channel=9
    -6, -3, 10, -2, -9, -2, -14, 5, -1,
    -- filter=53 channel=10
    -9, 12, 9, 6, 10, 6, 0, -11, 4,
    -- filter=53 channel=11
    -16, -13, -12, -17, -16, -7, 0, -3, -2,
    -- filter=53 channel=12
    10, -10, 10, -7, -9, -7, -2, 1, 10,
    -- filter=53 channel=13
    6, -9, 7, -1, 7, -5, -7, 11, 0,
    -- filter=53 channel=14
    -15, -4, -14, -14, 3, 4, 5, 4, 2,
    -- filter=53 channel=15
    -4, -9, 13, 15, 8, -12, -6, -8, 5,
    -- filter=53 channel=16
    -11, -3, -6, -13, -5, -10, 0, 0, -11,
    -- filter=53 channel=17
    -13, -8, 6, 5, 11, 5, 7, -5, 3,
    -- filter=53 channel=18
    -3, -5, -7, 8, -7, 2, 5, -6, -14,
    -- filter=53 channel=19
    10, -2, 0, 6, -8, 0, 9, 9, -2,
    -- filter=53 channel=20
    -11, 5, -14, 8, 11, 1, -6, 2, 10,
    -- filter=53 channel=21
    10, 15, -1, 15, -2, 9, 6, -5, 7,
    -- filter=53 channel=22
    7, -5, 4, -2, -2, -10, -9, -12, 2,
    -- filter=53 channel=23
    0, 6, 12, -8, -15, -13, -16, -14, 1,
    -- filter=53 channel=24
    -4, -11, -13, -12, -4, -6, -6, 9, 0,
    -- filter=53 channel=25
    -2, 2, -9, -12, 2, -12, -6, -13, -8,
    -- filter=53 channel=26
    1, 3, 7, 9, 15, -11, 5, 0, 3,
    -- filter=53 channel=27
    -2, -10, -2, 4, 4, 8, -3, 3, 0,
    -- filter=53 channel=28
    0, -9, -11, -5, -5, -1, -12, -9, -9,
    -- filter=53 channel=29
    5, -15, 8, 0, -12, -8, 6, 0, 9,
    -- filter=53 channel=30
    4, -5, -14, 6, 7, -9, -2, -14, -2,
    -- filter=53 channel=31
    12, 11, 6, 9, 16, -7, -12, -5, 7,
    -- filter=54 channel=0
    -2, -7, -5, 11, -11, -13, 4, 12, -8,
    -- filter=54 channel=1
    -12, 11, -7, 2, -6, 6, -13, -4, 0,
    -- filter=54 channel=2
    -4, 10, 10, -9, -5, 4, -14, 3, 4,
    -- filter=54 channel=3
    -9, -5, -5, -4, 0, 0, 4, 13, 14,
    -- filter=54 channel=4
    1, -4, -5, -2, 8, 14, 0, -14, 4,
    -- filter=54 channel=5
    -1, 14, 3, 5, 1, 12, -2, -3, -11,
    -- filter=54 channel=6
    1, -13, 8, 5, -12, 13, -10, -1, -8,
    -- filter=54 channel=7
    -11, -4, 10, -3, 9, 16, -12, 13, -8,
    -- filter=54 channel=8
    6, 12, 9, 3, -2, -1, -3, 5, -15,
    -- filter=54 channel=9
    2, -15, 8, 1, -5, -9, -1, 0, -13,
    -- filter=54 channel=10
    0, 14, -8, 9, 5, 0, 1, 4, -8,
    -- filter=54 channel=11
    4, 1, -6, 7, 8, -7, 4, 2, 5,
    -- filter=54 channel=12
    15, -3, 9, 0, 8, -9, 14, -8, -5,
    -- filter=54 channel=13
    4, 9, -9, 6, 11, -1, -3, 16, 17,
    -- filter=54 channel=14
    -2, 12, -11, 11, 2, -4, -9, 0, 3,
    -- filter=54 channel=15
    -14, 1, -8, 7, 12, 4, -7, 11, -3,
    -- filter=54 channel=16
    8, 13, 8, 0, 3, -9, -15, -2, 4,
    -- filter=54 channel=17
    -14, 9, 17, -3, -9, 3, -6, -7, 8,
    -- filter=54 channel=18
    -5, 6, -4, 13, -11, 13, 13, 1, 13,
    -- filter=54 channel=19
    4, 4, 13, -1, 4, -6, 0, -4, 12,
    -- filter=54 channel=20
    -11, -9, 5, 8, 13, 1, -6, 2, 3,
    -- filter=54 channel=21
    2, -12, -1, 5, 3, -8, -3, -5, 11,
    -- filter=54 channel=22
    0, -8, -8, -2, 0, 0, -8, -14, -4,
    -- filter=54 channel=23
    8, -13, -6, -6, 0, -12, 13, 3, 4,
    -- filter=54 channel=24
    2, -12, 0, -2, 2, -2, -14, 8, 6,
    -- filter=54 channel=25
    -8, -12, 1, -13, 8, -2, -3, -3, 7,
    -- filter=54 channel=26
    -4, 1, -7, -1, -1, 4, 11, -13, 0,
    -- filter=54 channel=27
    1, -6, -1, 11, 1, 9, 12, 11, -12,
    -- filter=54 channel=28
    5, -11, 11, -14, -14, -4, 7, 0, -1,
    -- filter=54 channel=29
    -12, -2, -10, -15, -9, 12, 0, -7, 6,
    -- filter=54 channel=30
    -14, 7, -12, 3, -10, 3, 12, 1, 3,
    -- filter=54 channel=31
    4, 0, 17, -10, 15, 12, -5, -14, 4,
    -- filter=55 channel=0
    -8, 1, -14, 9, 4, -10, -17, 6, 9,
    -- filter=55 channel=1
    -7, -15, 12, 0, 7, -13, -13, 1, -3,
    -- filter=55 channel=2
    -8, 12, 4, -12, 11, 6, -4, 1, -9,
    -- filter=55 channel=3
    13, -8, 9, 14, -9, 10, 11, -7, 7,
    -- filter=55 channel=4
    7, -5, 13, -1, 11, 5, -16, -1, -10,
    -- filter=55 channel=5
    6, 12, -1, -4, 11, -15, -2, -10, -5,
    -- filter=55 channel=6
    9, 12, 14, -10, -14, 11, -3, -13, -13,
    -- filter=55 channel=7
    6, -5, 3, 20, 4, -8, 4, -10, 1,
    -- filter=55 channel=8
    -8, -6, -15, 8, 9, -12, -7, -12, 11,
    -- filter=55 channel=9
    -3, -2, -4, 0, 1, -10, 5, -11, 9,
    -- filter=55 channel=10
    12, -2, -12, 4, -3, -13, 1, -10, -2,
    -- filter=55 channel=11
    10, 14, 8, 17, 1, -12, 11, 0, -7,
    -- filter=55 channel=12
    -11, -13, 0, 12, 11, -4, 6, -14, -11,
    -- filter=55 channel=13
    14, -16, -8, 0, 1, 4, 6, -8, 8,
    -- filter=55 channel=14
    -18, -4, -4, -11, -15, -5, -15, -14, 12,
    -- filter=55 channel=15
    -3, -3, -13, -4, 10, 9, -9, -13, 8,
    -- filter=55 channel=16
    10, -4, 11, -12, -13, -6, -2, -15, 6,
    -- filter=55 channel=17
    22, 3, 8, 17, -16, -14, 12, -17, -13,
    -- filter=55 channel=18
    0, -6, -1, -16, 12, 0, -16, -6, 4,
    -- filter=55 channel=19
    11, -3, -10, -11, -11, 0, -1, -5, -6,
    -- filter=55 channel=20
    11, 18, 2, 18, 11, 15, -3, 11, -6,
    -- filter=55 channel=21
    11, 4, -1, 18, 5, 9, 13, -8, -11,
    -- filter=55 channel=22
    7, 13, -3, 10, -3, -11, 8, 12, -11,
    -- filter=55 channel=23
    -12, -4, 9, -5, 13, -5, -8, -8, -1,
    -- filter=55 channel=24
    -2, 4, -13, -12, 9, -4, 2, 2, -3,
    -- filter=55 channel=25
    9, 4, 2, 0, -15, -13, 5, 4, 11,
    -- filter=55 channel=26
    9, -11, -16, -10, -1, -21, 1, 1, -14,
    -- filter=55 channel=27
    1, 14, 10, -11, -14, 7, -6, -6, -3,
    -- filter=55 channel=28
    9, 0, -1, 15, 9, -11, 8, -10, 9,
    -- filter=55 channel=29
    11, -9, -8, -14, 14, 2, 2, 1, 5,
    -- filter=55 channel=30
    -2, -2, -13, 0, 13, 11, -13, -4, 13,
    -- filter=55 channel=31
    4, -7, 0, 0, -9, -14, -16, -17, 6,
    -- filter=56 channel=0
    3, -8, 8, -8, 9, 5, 6, -13, -9,
    -- filter=56 channel=1
    16, -4, 7, 7, 9, -5, 4, 10, -10,
    -- filter=56 channel=2
    -4, 5, 13, -6, 6, -1, -14, 3, 0,
    -- filter=56 channel=3
    5, -3, 6, 9, -2, -5, -2, 0, 2,
    -- filter=56 channel=4
    -6, -3, 0, -8, 11, 8, 10, 3, 0,
    -- filter=56 channel=5
    0, 0, 7, 12, 10, -5, 0, 10, -7,
    -- filter=56 channel=6
    -5, -9, -5, 5, -1, -7, -12, 13, 5,
    -- filter=56 channel=7
    12, 16, -6, -10, 7, 7, 2, -15, 6,
    -- filter=56 channel=8
    -12, 8, 8, -2, 6, 6, 12, -14, -14,
    -- filter=56 channel=9
    -17, -13, 2, -4, 0, -5, -11, 8, 1,
    -- filter=56 channel=10
    2, 3, -14, -5, -6, -1, -15, -11, 8,
    -- filter=56 channel=11
    -1, -14, 6, 5, 2, 8, -5, 15, -12,
    -- filter=56 channel=12
    -9, 3, 1, 9, -2, -3, 2, -18, -2,
    -- filter=56 channel=13
    0, 2, 8, 12, 9, 14, 11, 0, -10,
    -- filter=56 channel=14
    5, 9, 12, -11, 11, -10, 3, 15, 13,
    -- filter=56 channel=15
    16, 0, 9, 3, 0, -5, 14, -15, 3,
    -- filter=56 channel=16
    10, -5, -3, -1, 10, 1, 9, -2, 4,
    -- filter=56 channel=17
    -2, 3, 15, -2, -7, -10, 4, 8, 0,
    -- filter=56 channel=18
    17, 8, 16, 19, 1, 17, 14, -9, -8,
    -- filter=56 channel=19
    -10, 6, -11, 10, 7, 6, -10, 1, 8,
    -- filter=56 channel=20
    13, 14, 14, 4, 23, 22, 4, 21, -5,
    -- filter=56 channel=21
    1, -13, -19, -4, -15, -22, -9, -20, -20,
    -- filter=56 channel=22
    -7, -16, 0, -11, -12, -6, -6, -25, -21,
    -- filter=56 channel=23
    -8, 3, -14, -11, 8, -7, 10, -16, -7,
    -- filter=56 channel=24
    -6, 9, 18, -9, 20, -5, 11, -3, 18,
    -- filter=56 channel=25
    -10, -20, -16, -1, -7, -19, -7, -7, -15,
    -- filter=56 channel=26
    8, 10, -11, -6, -13, 1, 13, -12, 12,
    -- filter=56 channel=27
    -9, -3, -1, -3, 9, -8, 8, 10, -14,
    -- filter=56 channel=28
    10, -9, 12, -13, -11, 0, -14, 3, -11,
    -- filter=56 channel=29
    1, 12, -4, 6, 13, -1, 8, 13, -4,
    -- filter=56 channel=30
    -12, 10, -9, -1, 7, -11, 14, -2, 13,
    -- filter=56 channel=31
    0, 4, 2, -15, -8, 1, 10, -14, 8,
    -- filter=57 channel=0
    -12, 14, 13, 12, 0, 11, -9, -10, 0,
    -- filter=57 channel=1
    9, 9, -17, -13, -1, -11, -9, 0, -17,
    -- filter=57 channel=2
    5, 0, -1, 7, -13, 4, 7, 8, 0,
    -- filter=57 channel=3
    0, -9, 2, 14, 6, -7, 7, -1, 5,
    -- filter=57 channel=4
    -19, -5, -17, -12, 0, -24, -12, -3, -24,
    -- filter=57 channel=5
    4, 12, 11, 14, -2, -12, -2, -15, -7,
    -- filter=57 channel=6
    5, -11, 10, 5, -11, 2, 15, 8, 15,
    -- filter=57 channel=7
    4, -12, -13, -13, -2, -1, -6, 7, -7,
    -- filter=57 channel=8
    6, -4, -11, -5, -14, 4, 0, 8, 14,
    -- filter=57 channel=9
    -4, 12, 10, 0, -5, 6, 10, -12, -11,
    -- filter=57 channel=10
    -2, 11, 0, -12, 9, 2, 8, -15, 1,
    -- filter=57 channel=11
    8, 2, 13, -8, 1, 19, 14, -8, 18,
    -- filter=57 channel=12
    9, 16, 7, 13, 9, 8, 7, 16, 5,
    -- filter=57 channel=13
    5, 23, 1, 20, 25, 19, 15, 11, 9,
    -- filter=57 channel=14
    -18, -16, 8, 6, -7, -13, 10, -1, 5,
    -- filter=57 channel=15
    15, 13, 4, 20, 1, 0, 13, 14, 13,
    -- filter=57 channel=16
    -9, -11, -1, 15, 0, 4, 1, 0, 12,
    -- filter=57 channel=17
    7, -3, -3, -13, -10, -1, -13, 4, 5,
    -- filter=57 channel=18
    6, -16, -19, -9, -2, -14, 11, -9, -13,
    -- filter=57 channel=19
    0, 6, 5, 2, -14, 10, 10, 10, 14,
    -- filter=57 channel=20
    5, 6, 8, -9, 11, -13, 2, -13, -9,
    -- filter=57 channel=21
    10, -10, 5, 0, -20, -9, 7, -16, -16,
    -- filter=57 channel=22
    3, 5, 8, 9, -15, -10, -10, -5, 1,
    -- filter=57 channel=23
    -2, -15, 0, 1, -3, 1, 1, -8, 1,
    -- filter=57 channel=24
    1, -5, 2, 0, -13, 7, 3, -9, -12,
    -- filter=57 channel=25
    -8, -8, -23, -6, -19, -10, -7, -28, -26,
    -- filter=57 channel=26
    19, 17, 13, 4, 12, 19, -2, -3, 17,
    -- filter=57 channel=27
    7, 0, 9, -14, 11, -7, -12, -12, 11,
    -- filter=57 channel=28
    9, -14, 0, 7, -13, -2, 4, -8, 6,
    -- filter=57 channel=29
    9, 11, 6, 7, 0, -9, 15, -11, -9,
    -- filter=57 channel=30
    2, -12, 3, 0, -10, 10, 14, -7, 10,
    -- filter=57 channel=31
    -8, -7, 9, -5, 11, -10, 6, 3, 6,
    -- filter=58 channel=0
    0, 9, 10, 8, 10, 10, 10, 1, -12,
    -- filter=58 channel=1
    -7, 2, -14, 0, -7, 1, 1, -8, -14,
    -- filter=58 channel=2
    -2, 14, -12, -7, 2, 13, 9, -14, -7,
    -- filter=58 channel=3
    -11, -5, 14, 6, -1, -9, -2, 5, -13,
    -- filter=58 channel=4
    -8, -6, 4, -11, 6, 1, -7, -1, 3,
    -- filter=58 channel=5
    -5, 9, -4, -13, 3, -7, -3, 4, 9,
    -- filter=58 channel=6
    -6, -7, -13, -3, -4, -13, -8, -1, 2,
    -- filter=58 channel=7
    -5, -3, 13, -7, -11, -6, 11, 3, 5,
    -- filter=58 channel=8
    -14, -10, -1, 11, -12, -9, 14, -7, 7,
    -- filter=58 channel=9
    -9, 8, -14, 2, 5, 13, 15, -9, -12,
    -- filter=58 channel=10
    -9, -6, 1, -9, 1, 1, 2, 2, 9,
    -- filter=58 channel=11
    4, -10, -13, 10, -12, 3, -9, -1, 9,
    -- filter=58 channel=12
    13, -9, -9, 8, 5, -3, -6, 0, -4,
    -- filter=58 channel=13
    0, 0, 14, 0, 10, 8, 6, 6, 2,
    -- filter=58 channel=14
    7, 6, -6, -14, -10, 0, -2, 1, 7,
    -- filter=58 channel=15
    -4, -6, -14, -5, -6, -4, -5, 9, -6,
    -- filter=58 channel=16
    -13, -13, 6, -12, 14, 10, -6, -14, -13,
    -- filter=58 channel=17
    0, -1, 3, 12, -5, 10, -13, -3, -3,
    -- filter=58 channel=18
    6, 1, 10, 5, -8, 1, -10, 2, -13,
    -- filter=58 channel=19
    11, -1, 2, -1, -10, 13, 12, 1, -2,
    -- filter=58 channel=20
    -1, 10, -4, -9, -11, -6, 11, 8, -11,
    -- filter=58 channel=21
    2, 2, 13, 4, -5, 1, 11, -11, 1,
    -- filter=58 channel=22
    -5, 14, 3, 0, 11, -3, 1, 8, 6,
    -- filter=58 channel=23
    0, -8, -5, 5, -10, 4, 9, -5, 8,
    -- filter=58 channel=24
    8, 9, 3, -12, -10, -13, -5, -4, 13,
    -- filter=58 channel=25
    -5, 0, -6, 15, 6, -13, 11, 9, 7,
    -- filter=58 channel=26
    -11, 2, -2, 13, 7, 7, -11, -5, -14,
    -- filter=58 channel=27
    -14, 6, -6, 4, 4, 13, 0, 8, -4,
    -- filter=58 channel=28
    -13, 0, -4, -7, -6, -9, -12, -10, 2,
    -- filter=58 channel=29
    -10, -9, -1, -14, -12, -4, -6, 8, -13,
    -- filter=58 channel=30
    -12, 7, 1, -10, -14, -7, -9, 3, 9,
    -- filter=58 channel=31
    -10, 9, 10, -13, -2, -11, -8, -1, -1,
    -- filter=59 channel=0
    1, -5, -2, 12, 7, -14, -1, 6, 12,
    -- filter=59 channel=1
    5, 10, 9, 0, -14, -9, -1, 10, 6,
    -- filter=59 channel=2
    10, 8, 7, -8, 0, -3, -3, -13, 0,
    -- filter=59 channel=3
    -11, 1, 6, -10, 9, -13, 0, 9, 8,
    -- filter=59 channel=4
    11, 3, -1, 17, 3, 1, 0, 5, -8,
    -- filter=59 channel=5
    9, -5, 14, -5, 12, -6, 6, 3, 3,
    -- filter=59 channel=6
    7, 4, 4, 2, 2, -3, 5, 2, 0,
    -- filter=59 channel=7
    0, -5, -11, 4, -10, -9, 8, -9, -17,
    -- filter=59 channel=8
    14, 5, 2, 7, 11, 12, -8, 7, 14,
    -- filter=59 channel=9
    0, 6, -3, 10, -6, 9, 6, 2, -1,
    -- filter=59 channel=10
    -11, -7, 11, -7, -8, -2, 13, 9, 16,
    -- filter=59 channel=11
    4, -4, 5, -19, -10, -17, -14, 1, -17,
    -- filter=59 channel=12
    -2, -5, 0, -8, -15, -7, 11, 7, -1,
    -- filter=59 channel=13
    0, 6, -5, -9, -10, 3, -7, 3, 13,
    -- filter=59 channel=14
    11, 5, -11, -12, -17, 2, -7, -6, -7,
    -- filter=59 channel=15
    -6, -1, -13, 10, -12, -8, 0, -2, 0,
    -- filter=59 channel=16
    8, -7, -8, 10, -14, 8, -7, 8, 9,
    -- filter=59 channel=17
    8, 6, 6, 15, -6, -11, 13, -6, 0,
    -- filter=59 channel=18
    9, -1, -9, -3, 9, 0, -9, -3, 10,
    -- filter=59 channel=19
    -7, 6, -8, 11, 9, 12, -1, -12, 8,
    -- filter=59 channel=20
    -14, 3, -13, -19, -7, -2, 6, -12, -4,
    -- filter=59 channel=21
    16, 18, 0, -4, -10, 7, 6, 8, 3,
    -- filter=59 channel=22
    -3, -1, 4, -5, 14, 9, -12, -11, -9,
    -- filter=59 channel=23
    -6, 2, -12, -3, -5, -3, 14, 12, -1,
    -- filter=59 channel=24
    -12, 4, -12, -6, -16, 7, -3, -1, -15,
    -- filter=59 channel=25
    21, 15, 7, 18, 2, -1, 14, 10, 17,
    -- filter=59 channel=26
    2, -8, -2, -10, -7, -2, -9, 5, -13,
    -- filter=59 channel=27
    -2, -8, 3, -7, -8, -9, 3, 5, 8,
    -- filter=59 channel=28
    -5, 6, 12, -2, 0, -11, -3, 0, -1,
    -- filter=59 channel=29
    -11, -20, -4, -16, -11, 7, -16, -10, -14,
    -- filter=59 channel=30
    14, -13, -14, 0, -11, 12, 2, -10, 12,
    -- filter=59 channel=31
    -11, -2, 9, -2, 4, -8, -6, -10, 8,
    -- filter=60 channel=0
    6, -5, 16, -1, 14, 22, 3, -5, 23,
    -- filter=60 channel=1
    -2, -11, -15, -4, -11, 1, -5, -19, -21,
    -- filter=60 channel=2
    13, -6, 2, -2, 14, -1, 8, -11, -6,
    -- filter=60 channel=3
    13, 8, -13, -12, -4, 3, -6, -2, 8,
    -- filter=60 channel=4
    -24, -27, -27, 3, -10, -18, 3, -13, -28,
    -- filter=60 channel=5
    -7, -15, 1, -9, 7, 0, -15, 11, 8,
    -- filter=60 channel=6
    9, 0, -1, 2, -14, -8, -9, 4, -7,
    -- filter=60 channel=7
    -13, -9, -11, -11, 10, -4, 6, -2, 0,
    -- filter=60 channel=8
    15, 9, 17, 20, 19, 21, 15, 11, 20,
    -- filter=60 channel=9
    -7, -6, 1, 5, -9, 7, 7, -14, -7,
    -- filter=60 channel=10
    -7, -8, -12, -3, -15, -7, 13, -5, -5,
    -- filter=60 channel=11
    17, 21, 13, 30, 26, 33, 4, 27, 37,
    -- filter=60 channel=12
    12, 13, -10, 6, -12, -11, 4, 12, -12,
    -- filter=60 channel=13
    2, 18, 23, -8, 9, 9, -4, 12, 12,
    -- filter=60 channel=14
    -12, 12, 9, 0, 0, 9, -15, -9, -10,
    -- filter=60 channel=15
    -11, 13, 1, -11, -6, -15, 4, -7, -8,
    -- filter=60 channel=16
    13, 4, -14, -13, 4, -5, 0, -16, -1,
    -- filter=60 channel=17
    9, -10, 7, 11, 11, -13, -14, 3, -15,
    -- filter=60 channel=18
    -18, 4, -15, -5, 4, -8, -16, -9, -15,
    -- filter=60 channel=19
    -2, 3, -11, 5, 3, -11, 10, -2, 13,
    -- filter=60 channel=20
    5, -18, -1, -10, 4, -6, -7, 1, 8,
    -- filter=60 channel=21
    -12, -21, -20, -9, -16, -15, -18, 0, -17,
    -- filter=60 channel=22
    7, -19, -13, -17, -12, -13, -15, -13, -19,
    -- filter=60 channel=23
    -15, -12, 0, -5, 2, -11, -2, -3, -9,
    -- filter=60 channel=24
    3, 4, -3, 4, -7, 9, 11, 14, -14,
    -- filter=60 channel=25
    -11, -18, -34, -5, -28, -4, 3, -28, -31,
    -- filter=60 channel=26
    12, -1, 19, 12, 12, -4, -2, 16, 6,
    -- filter=60 channel=27
    -12, 9, 14, -4, 3, 0, 6, 10, 0,
    -- filter=60 channel=28
    -17, 0, -15, -3, -15, -4, 7, 0, -1,
    -- filter=60 channel=29
    23, 17, 18, 18, 30, 20, 24, 17, 29,
    -- filter=60 channel=30
    -1, -5, 6, -1, 3, -2, 13, -5, 6,
    -- filter=60 channel=31
    -6, -1, -10, -2, -5, -18, -20, -3, -14,
    -- filter=61 channel=0
    -13, 10, -14, 8, -9, -14, 1, 7, -1,
    -- filter=61 channel=1
    -7, -8, 1, 13, 12, -1, -11, -2, -3,
    -- filter=61 channel=2
    2, -6, -13, 10, -7, -1, 8, 10, 9,
    -- filter=61 channel=3
    -2, -2, 5, -2, 12, 12, 5, 7, 13,
    -- filter=61 channel=4
    12, 12, 4, 4, -7, 14, -12, -13, 1,
    -- filter=61 channel=5
    0, 5, -12, -6, 8, -8, 10, -7, 14,
    -- filter=61 channel=6
    -7, -8, -10, 2, -1, -7, 12, 10, 10,
    -- filter=61 channel=7
    5, 4, -14, -8, 7, -7, 10, 1, 8,
    -- filter=61 channel=8
    6, -13, 4, -7, 6, -8, 3, 4, -1,
    -- filter=61 channel=9
    2, 0, -9, 0, 2, 13, 5, 12, 11,
    -- filter=61 channel=10
    7, -8, -6, -13, -4, 1, 10, 0, 11,
    -- filter=61 channel=11
    6, -22, 1, -9, -3, 5, -10, -9, -19,
    -- filter=61 channel=12
    7, -6, 11, -2, -2, -4, -5, -4, 5,
    -- filter=61 channel=13
    -17, -1, -6, -4, -6, 8, 7, -10, -16,
    -- filter=61 channel=14
    -5, -11, -7, 6, -11, 4, -20, -15, 12,
    -- filter=61 channel=15
    12, -11, 5, 6, 12, 5, 9, -5, 4,
    -- filter=61 channel=16
    -14, -8, -5, 0, 0, 4, 7, -15, 4,
    -- filter=61 channel=17
    -8, 5, 1, -8, -5, 4, 0, -6, 13,
    -- filter=61 channel=18
    4, -5, -14, 1, -14, -7, 0, 8, -4,
    -- filter=61 channel=19
    -5, -14, 7, -11, 12, 0, 11, -9, -2,
    -- filter=61 channel=20
    -18, -20, -9, 0, -7, 14, 1, 12, 13,
    -- filter=61 channel=21
    15, 14, 13, 12, 11, 16, 18, 7, 4,
    -- filter=61 channel=22
    9, 11, -11, 0, 6, 0, -2, -3, -2,
    -- filter=61 channel=23
    -15, -11, 4, -7, -4, 5, 2, 2, 11,
    -- filter=61 channel=24
    5, -6, 3, 4, -5, 0, 5, 0, -9,
    -- filter=61 channel=25
    5, -1, 0, 4, -1, 2, -7, 11, -11,
    -- filter=61 channel=26
    -10, -4, 6, 7, 5, -7, -4, 2, -1,
    -- filter=61 channel=27
    -7, -3, -12, -11, -13, -1, -1, 0, -1,
    -- filter=61 channel=28
    -14, -8, 9, -14, 8, 2, -3, -12, -13,
    -- filter=61 channel=29
    -4, -22, -5, -6, -9, -10, -7, -13, -6,
    -- filter=61 channel=30
    -3, -3, -13, -6, 9, -12, 5, -2, -9,
    -- filter=61 channel=31
    -8, -12, 5, -1, -6, -1, 12, -1, 16,
    -- filter=62 channel=0
    2, 10, -12, -4, -7, -9, -1, -6, -13,
    -- filter=62 channel=1
    0, -3, 1, -6, 14, 7, -1, -2, 10,
    -- filter=62 channel=2
    -9, -3, -3, 0, 13, 9, 14, 0, 13,
    -- filter=62 channel=3
    5, 3, 0, 8, -8, -4, 7, -15, -8,
    -- filter=62 channel=4
    -13, 5, -4, -1, 5, 14, -9, -3, 4,
    -- filter=62 channel=5
    9, -2, -15, 0, 4, -5, -13, 7, -10,
    -- filter=62 channel=6
    11, -5, 7, -1, 11, 8, 9, -13, 6,
    -- filter=62 channel=7
    -7, -9, -6, 6, 9, 4, -10, 13, 14,
    -- filter=62 channel=8
    -3, -1, -9, -4, 0, -7, -1, 3, -4,
    -- filter=62 channel=9
    -7, 4, -1, 0, 7, -8, -6, 6, 2,
    -- filter=62 channel=10
    -13, 4, 3, -16, -7, -17, -8, -13, -8,
    -- filter=62 channel=11
    2, 7, 3, 17, -9, 0, 1, -8, 7,
    -- filter=62 channel=12
    -1, 7, 8, -13, -6, -14, 5, 0, 8,
    -- filter=62 channel=13
    -4, -21, -11, -20, -5, 2, -23, -24, -7,
    -- filter=62 channel=14
    -8, 0, 18, 15, 16, 11, 4, 10, 0,
    -- filter=62 channel=15
    -19, -13, -17, 3, -1, 0, -3, -10, -8,
    -- filter=62 channel=16
    1, 2, -1, 11, 11, 3, 2, -10, -9,
    -- filter=62 channel=17
    8, -9, 4, -18, 12, 5, 8, 4, 9,
    -- filter=62 channel=18
    -11, 7, 0, 4, 11, -11, -2, 6, 9,
    -- filter=62 channel=19
    -13, -1, -5, 8, -9, 3, -5, 0, -6,
    -- filter=62 channel=20
    5, 14, 23, 4, 12, 0, 16, -6, 15,
    -- filter=62 channel=21
    -19, -15, 1, -23, -13, 1, -9, 6, 5,
    -- filter=62 channel=22
    4, -9, -8, 2, -9, -12, -3, -14, 7,
    -- filter=62 channel=23
    -2, 9, -7, -18, 11, -2, -1, -1, 8,
    -- filter=62 channel=24
    0, 10, 1, -9, 0, 12, -2, -4, 2,
    -- filter=62 channel=25
    0, -5, -12, 6, -6, -7, -3, -8, -4,
    -- filter=62 channel=26
    -15, -13, -16, -7, -2, 1, -17, -5, -18,
    -- filter=62 channel=27
    -13, -14, 5, -6, 11, 9, -14, 7, 13,
    -- filter=62 channel=28
    0, -11, 7, 6, 14, 1, -8, 12, 15,
    -- filter=62 channel=29
    10, -7, -9, 17, -2, 13, 11, -1, -4,
    -- filter=62 channel=30
    -9, -6, 9, -7, 9, -8, -1, 11, 7,
    -- filter=62 channel=31
    -23, -8, -13, -13, -21, -4, -12, -20, -12,
    -- filter=63 channel=0
    12, -7, 9, 13, -10, 11, 11, 12, 10,
    -- filter=63 channel=1
    5, -19, -19, -7, -4, 5, -8, 5, -4,
    -- filter=63 channel=2
    1, -1, 8, 9, 12, 14, 13, -4, -4,
    -- filter=63 channel=3
    -11, -3, 0, -1, 13, -10, -10, 2, -10,
    -- filter=63 channel=4
    -4, -15, -12, -14, -11, 8, -6, 3, -3,
    -- filter=63 channel=5
    0, 6, 0, -6, 1, -3, 11, 13, 10,
    -- filter=63 channel=6
    12, -7, 4, 8, 9, 9, -14, 14, 0,
    -- filter=63 channel=7
    6, -12, -5, 9, -18, 2, 0, -13, -19,
    -- filter=63 channel=8
    6, 13, -3, 9, -6, 1, -4, -2, 8,
    -- filter=63 channel=9
    -4, 5, 12, -7, -8, 2, -14, -5, 6,
    -- filter=63 channel=10
    2, -1, 0, -6, 11, -13, -11, 9, -9,
    -- filter=63 channel=11
    -6, 12, -1, 0, -12, -9, 0, 11, 5,
    -- filter=63 channel=12
    8, 5, -5, -1, -2, 10, -4, 14, -13,
    -- filter=63 channel=13
    6, 27, 8, 21, 11, 11, 15, 18, 25,
    -- filter=63 channel=14
    5, -13, -12, -11, 0, 2, -10, -10, -3,
    -- filter=63 channel=15
    2, 10, 9, 0, 0, 5, 14, 20, 2,
    -- filter=63 channel=16
    -11, 3, -15, 5, -10, -7, 3, -11, -15,
    -- filter=63 channel=17
    14, 3, -9, -3, 9, -11, 8, 0, -5,
    -- filter=63 channel=18
    -3, 8, -3, -5, -11, 6, -13, 9, -7,
    -- filter=63 channel=19
    -9, 0, 4, 7, -12, -11, 11, 3, -5,
    -- filter=63 channel=20
    1, -2, 4, -6, -15, 0, -3, -17, -8,
    -- filter=63 channel=21
    4, -17, -19, -20, -18, 6, -8, -7, 7,
    -- filter=63 channel=22
    -15, -8, 0, -7, -4, -18, -18, -6, 0,
    -- filter=63 channel=23
    -15, -7, -12, -18, -10, -3, 0, 6, -6,
    -- filter=63 channel=24
    0, -13, -6, -20, -12, -13, 4, 5, -17,
    -- filter=63 channel=25
    -18, -25, -4, -10, -25, -18, -25, -3, -4,
    -- filter=63 channel=26
    -2, -3, 10, 25, 22, 9, 12, 18, 14,
    -- filter=63 channel=27
    2, 10, -9, 4, 3, 11, -4, 4, 11,
    -- filter=63 channel=28
    3, -8, -16, 7, -14, 10, -2, -10, 6,
    -- filter=63 channel=29
    11, -11, -10, -5, -8, -7, 0, -16, 0,
    -- filter=63 channel=30
    12, -9, 11, 4, 2, -12, 10, -8, 14,
    -- filter=63 channel=31
    20, 15, 8, 0, 8, -9, 7, 10, 12,

    others => 0);
end iwght_package;
