library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package ifmap_package is
  type mem is array(0 to 4000000) of integer;

  constant input_map : mem := (

    -- ifmap
    -- channel=0
    861, 879, 868, 823, 508, 353, 561, 
    433, 795, 649, 283, 217, 135, 174, 
    159, 741, 520, 262, 304, 149, 55, 
    51, 369, 450, 165, 292, 153, 124, 
    22, 107, 78, 114, 171, 58, 131, 
    0, 245, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    945, 985, 1021, 837, 527, 380, 603, 
    610, 1003, 805, 421, 284, 336, 237, 
    440, 787, 794, 610, 445, 380, 236, 
    328, 591, 502, 453, 404, 345, 315, 
    257, 414, 289, 304, 213, 37, 190, 
    0, 358, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=2
    0, 12, 0, 0, 0, 0, 0, 
    121, 136, 156, 53, 12, 18, 0, 
    24, 0, 0, 157, 154, 0, 103, 
    129, 50, 0, 0, 0, 0, 40, 
    70, 273, 263, 209, 0, 0, 17, 
    0, 13, 0, 0, 30, 137, 97, 
    0, 0, 25, 121, 142, 112, 134, 
    
    -- channel=3
    175, 24, 73, 642, 35, 0, 302, 
    0, 0, 0, 0, 66, 0, 181, 
    0, 638, 168, 0, 0, 84, 0, 
    0, 0, 720, 431, 308, 351, 11, 
    0, 0, 0, 0, 449, 9, 0, 
    690, 160, 1222, 935, 32, 0, 0, 
    486, 1291, 241, 0, 0, 142, 47, 
    
    -- channel=4
    0, 15, 2, 0, 1, 0, 0, 
    348, 494, 584, 292, 0, 3, 0, 
    0, 0, 18, 603, 418, 0, 389, 
    247, 121, 0, 0, 0, 0, 34, 
    38, 843, 785, 638, 0, 146, 0, 
    0, 0, 0, 0, 138, 312, 124, 
    0, 0, 5, 205, 242, 51, 113, 
    
    -- channel=5
    1372, 1421, 1219, 1124, 543, 453, 976, 
    674, 1179, 606, 70, 86, 0, 328, 
    0, 931, 146, 0, 0, 0, 0, 
    0, 387, 266, 0, 73, 0, 200, 
    0, 0, 0, 0, 0, 0, 262, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 132, 19, 0, 
    60, 0, 0, 0, 0, 25, 0, 
    134, 127, 33, 35, 0, 103, 0, 
    242, 344, 421, 373, 520, 650, 584, 
    715, 374, 644, 649, 739, 777, 855, 
    
    -- channel=7
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=8
    7, 0, 7, 0, 105, 0, 0, 
    283, 136, 99, 8, 184, 0, 43, 
    71, 147, 81, 0, 464, 0, 26, 
    0, 108, 36, 0, 139, 0, 59, 
    0, 370, 220, 76, 0, 174, 90, 
    49, 252, 0, 0, 81, 98, 24, 
    77, 0, 106, 23, 60, 26, 62, 
    
    -- channel=9
    429, 451, 387, 255, 125, 98, 292, 
    185, 387, 132, 51, 144, 66, 96, 
    253, 242, 260, 23, 46, 64, 77, 
    87, 159, 192, 113, 131, 77, 234, 
    97, 24, 36, 50, 4, 0, 196, 
    171, 14, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 0, 
    
    -- channel=10
    330, 322, 327, 404, 212, 222, 300, 
    148, 201, 111, 137, 183, 204, 207, 
    356, 354, 299, 157, 58, 294, 113, 
    304, 249, 473, 419, 345, 332, 207, 
    410, 97, 43, 165, 355, 119, 214, 
    531, 426, 584, 476, 180, 85, 212, 
    347, 770, 213, 109, 92, 178, 173, 
    
    -- channel=11
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 64, 46, 0, 
    0, 0, 0, 0, 23, 56, 138, 
    141, 0, 0, 0, 0, 98, 9, 
    294, 133, 125, 215, 127, 318, 92, 
    627, 316, 670, 811, 1032, 1202, 1182, 
    1217, 742, 1145, 1197, 1321, 1411, 1495, 
    
    -- channel=12
    0, 0, 267, 98, 96, 14, 0, 
    0, 0, 126, 0, 199, 52, 0, 
    315, 0, 55, 149, 338, 0, 84, 
    461, 53, 497, 54, 374, 0, 74, 
    519, 265, 0, 378, 178, 0, 138, 
    201, 961, 0, 138, 0, 62, 68, 
    0, 787, 32, 0, 59, 22, 174, 
    
    -- channel=13
    42, 19, 235, 239, 129, 93, 60, 
    0, 0, 93, 244, 209, 316, 50, 
    504, 49, 441, 477, 275, 404, 275, 
    605, 233, 508, 495, 383, 453, 186, 
    810, 359, 45, 447, 363, 167, 210, 
    717, 964, 577, 468, 379, 333, 391, 
    293, 1075, 411, 342, 353, 386, 486, 
    
    -- channel=14
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 14, 283, 191, 22, 
    343, 0, 362, 147, 327, 266, 157, 
    490, 23, 296, 328, 264, 278, 133, 
    712, 533, 263, 285, 243, 340, 137, 
    1153, 805, 1123, 1068, 969, 1102, 1139, 
    1321, 1198, 1168, 1163, 1237, 1404, 1447, 
    
    -- channel=16
    871, 875, 835, 767, 418, 313, 672, 
    431, 755, 358, 142, 175, 13, 273, 
    132, 540, 208, 0, 85, 4, 95, 
    0, 360, 313, 110, 205, 69, 264, 
    0, 0, 0, 0, 103, 0, 286, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=18
    0, 0, 0, 0, 0, 12, 0, 
    0, 0, 0, 194, 121, 398, 17, 
    628, 0, 449, 590, 271, 537, 224, 
    998, 123, 284, 456, 313, 463, 84, 
    1157, 665, 408, 598, 358, 194, 55, 
    1026, 1212, 1292, 1045, 914, 1021, 1075, 
    1217, 1396, 1131, 1150, 1228, 1328, 1499, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 0, 
    0, 0, 0, 0, 48, 58, 39, 
    0, 0, 12, 43, 45, 37, 24, 
    
    -- channel=20
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 161, 53, 0, 
    0, 0, 0, 0, 193, 54, 217, 
    259, 0, 0, 0, 0, 123, 24, 
    478, 324, 30, 212, 195, 541, 181, 
    1173, 669, 1247, 1509, 1771, 2135, 2100, 
    2254, 1525, 2062, 2157, 2365, 2576, 2687, 
    
    -- channel=21
    1204, 1317, 1178, 964, 655, 635, 932, 
    790, 1118, 831, 505, 432, 431, 554, 
    504, 788, 541, 448, 326, 379, 432, 
    214, 626, 542, 495, 496, 362, 634, 
    208, 110, 283, 298, 348, 123, 561, 
    0, 55, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=22
    0, 0, 0, 0, 0, 0, 10, 
    41, 0, 0, 0, 124, 0, 58, 
    109, 107, 101, 0, 196, 0, 0, 
    0, 60, 122, 62, 91, 48, 56, 
    14, 169, 0, 0, 11, 109, 14, 
    353, 180, 282, 240, 176, 164, 142, 
    382, 232, 248, 199, 202, 269, 258, 
    
    -- channel=23
    187, 0, 75, 228, 178, 31, 304, 
    69, 0, 0, 0, 798, 74, 248, 
    521, 889, 600, 0, 757, 178, 0, 
    202, 210, 1195, 454, 910, 364, 444, 
    532, 347, 0, 52, 372, 302, 467, 
    1507, 1264, 1225, 1139, 668, 869, 885, 
    1518, 1424, 1015, 841, 943, 1178, 1138, 
    
    -- channel=24
    134, 133, 111, 57, 18, 8, 64, 
    67, 119, 34, 0, 0, 0, 0, 
    0, 44, 0, 0, 0, 0, 0, 
    0, 26, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=25
    463, 492, 621, 311, 122, 197, 295, 
    323, 423, 358, 201, 257, 300, 33, 
    821, 173, 664, 542, 362, 294, 277, 
    779, 401, 515, 407, 429, 253, 390, 
    903, 485, 159, 578, 188, 0, 396, 
    470, 968, 0, 0, 0, 0, 0, 
    0, 493, 0, 0, 0, 0, 0, 
    
    -- channel=26
    655, 703, 563, 403, 287, 176, 429, 
    336, 650, 288, 60, 14, 0, 159, 
    0, 254, 0, 0, 0, 0, 61, 
    0, 133, 0, 0, 0, 0, 133, 
    0, 0, 0, 0, 0, 0, 149, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    568, 483, 612, 182, 326, 228, 457, 
    555, 595, 348, 115, 823, 239, 189, 
    1100, 702, 1216, 265, 1064, 252, 313, 
    867, 580, 1087, 435, 840, 222, 698, 
    1037, 960, 511, 759, 209, 82, 774, 
    1314, 1520, 236, 269, 281, 477, 493, 
    609, 645, 293, 351, 367, 421, 439, 
    
    -- channel=28
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=29
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 24, 0, 82, 
    389, 0, 0, 0, 0, 0, 0, 
    494, 305, 83, 273, 135, 350, 11, 
    998, 660, 1164, 1348, 1640, 2002, 2017, 
    2038, 1431, 1863, 1985, 2192, 2372, 2529, 
    
    -- channel=30
    622, 617, 664, 414, 286, 209, 422, 
    365, 608, 373, 168, 265, 79, 100, 
    422, 371, 466, 173, 344, 75, 153, 
    255, 312, 373, 71, 226, 52, 294, 
    247, 245, 130, 324, 41, 0, 419, 
    202, 385, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=31
    854, 825, 799, 538, 577, 379, 746, 
    470, 773, 298, 75, 698, 136, 384, 
    500, 693, 629, 0, 464, 20, 302, 
    90, 450, 845, 310, 613, 118, 746, 
    124, 64, 24, 192, 175, 73, 746, 
    536, 240, 0, 0, 0, 0, 0, 
    0, 102, 0, 0, 0, 0, 0, 
    
    -- channel=32
    152, 112, 277, 52, 29, 14, 74, 
    134, 5, 0, 8, 258, 142, 0, 
    696, 51, 509, 245, 424, 193, 163, 
    711, 203, 540, 321, 433, 237, 247, 
    857, 451, 44, 488, 156, 57, 300, 
    937, 1196, 528, 563, 440, 555, 572, 
    633, 1115, 598, 570, 633, 677, 835, 
    
    -- channel=33
    379, 305, 351, 457, 276, 201, 346, 
    81, 195, 73, 0, 397, 182, 136, 
    539, 612, 772, 44, 219, 225, 37, 
    434, 251, 882, 586, 587, 307, 337, 
    669, 199, 0, 153, 372, 70, 243, 
    956, 876, 725, 748, 70, 14, 145, 
    357, 1154, 131, 42, 11, 125, 132, 
    
    -- channel=34
    100, 0, 0, 0, 51, 0, 268, 
    760, 164, 0, 0, 713, 0, 205, 
    431, 593, 0, 0, 1322, 0, 0, 
    0, 178, 493, 0, 724, 0, 136, 
    0, 781, 103, 0, 0, 114, 363, 
    433, 778, 0, 0, 0, 115, 8, 
    617, 0, 231, 0, 9, 112, 52, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=36
    47, 60, 101, 0, 137, 159, 68, 
    202, 100, 167, 242, 186, 175, 195, 
    140, 0, 0, 267, 255, 152, 313, 
    202, 167, 0, 48, 135, 132, 208, 
    177, 271, 219, 319, 135, 225, 301, 
    50, 188, 0, 39, 279, 361, 333, 
    227, 127, 270, 290, 327, 293, 345, 
    
    -- channel=37
    1111, 1177, 1158, 884, 627, 432, 697, 
    613, 1151, 942, 421, 323, 200, 286, 
    146, 967, 682, 401, 408, 134, 174, 
    0, 536, 521, 180, 401, 180, 313, 
    0, 47, 183, 178, 67, 0, 205, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=38
    303, 269, 287, 246, 119, 94, 270, 
    101, 99, 0, 0, 220, 36, 116, 
    386, 288, 318, 0, 130, 10, 22, 
    154, 97, 497, 209, 314, 80, 258, 
    254, 0, 0, 32, 114, 0, 245, 
    487, 428, 171, 288, 7, 39, 83, 
    204, 522, 58, 61, 64, 107, 125, 
    
    -- channel=39
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 61, 61, 59, 0, 
    0, 0, 0, 50, 53, 66, 140, 
    159, 0, 0, 0, 0, 63, 9, 
    243, 100, 78, 194, 92, 233, 108, 
    419, 265, 394, 552, 740, 903, 883, 
    807, 597, 798, 873, 972, 1010, 1094, 
    
    -- channel=40
    0, 0, 0, 0, 64, 101, 19, 
    0, 0, 0, 75, 187, 172, 198, 
    32, 26, 12, 26, 74, 162, 210, 
    96, 9, 123, 144, 173, 245, 189, 
    168, 26, 31, 112, 215, 327, 185, 
    417, 184, 499, 646, 584, 679, 663, 
    801, 642, 656, 716, 754, 820, 824, 
    
    -- channel=41
    58, 310, 201, 506, 99, 226, 0, 
    0, 108, 514, 970, 0, 829, 201, 
    6, 0, 463, 1578, 0, 1427, 566, 
    773, 460, 0, 951, 0, 1311, 0, 
    731, 32, 455, 576, 575, 423, 0, 
    0, 0, 1409, 256, 373, 0, 0, 
    0, 797, 140, 49, 0, 0, 0, 
    
    -- channel=42
    442, 504, 498, 372, 271, 181, 251, 
    127, 440, 407, 248, 136, 170, 57, 
    59, 413, 416, 234, 91, 158, 101, 
    76, 181, 278, 180, 161, 160, 146, 
    171, 0, 158, 192, 64, 0, 81, 
    0, 145, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=43
    0, 0, 0, 238, 0, 0, 81, 
    0, 0, 0, 0, 132, 0, 94, 
    59, 285, 29, 0, 20, 83, 0, 
    0, 0, 406, 235, 247, 206, 0, 
    71, 0, 0, 0, 306, 177, 0, 
    623, 322, 993, 884, 357, 337, 393, 
    813, 1052, 557, 412, 440, 594, 580, 
    
    -- channel=44
    978, 1019, 989, 683, 521, 422, 677, 
    682, 967, 736, 234, 394, 148, 306, 
    388, 911, 693, 170, 456, 65, 148, 
    69, 544, 630, 203, 454, 48, 460, 
    0, 107, 187, 214, 44, 0, 407, 
    0, 189, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=45
    229, 238, 189, 144, 164, 147, 215, 
    71, 228, 171, 52, 160, 92, 109, 
    54, 90, 169, 0, 30, 0, 139, 
    36, 52, 99, 45, 92, 27, 202, 
    73, 0, 67, 68, 37, 109, 174, 
    139, 0, 0, 161, 115, 180, 145, 
    140, 79, 151, 227, 233, 240, 213, 
    
    -- channel=46
    22, 20, 0, 62, 0, 53, 22, 
    57, 22, 69, 123, 0, 104, 101, 
    27, 96, 0, 151, 0, 185, 42, 
    45, 87, 0, 90, 8, 153, 0, 
    0, 62, 159, 7, 93, 92, 0, 
    0, 0, 220, 0, 24, 0, 0, 
    66, 0, 26, 0, 0, 0, 0, 
    
    -- channel=47
    1597, 1691, 1597, 1312, 834, 732, 1170, 
    923, 1503, 1053, 474, 447, 374, 530, 
    593, 1216, 838, 408, 312, 306, 322, 
    154, 788, 792, 499, 573, 299, 645, 
    96, 9, 205, 271, 332, 0, 613, 
    0, 131, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=48
    847, 953, 944, 425, 297, 380, 524, 
    747, 903, 847, 444, 301, 296, 219, 
    638, 479, 626, 596, 504, 259, 318, 
    463, 587, 413, 172, 339, 121, 471, 
    362, 392, 488, 561, 0, 0, 397, 
    0, 361, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=49
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 150, 116, 14, 20, 0, 
    14, 0, 61, 299, 270, 10, 179, 
    345, 0, 0, 0, 0, 0, 0, 
    326, 551, 443, 428, 0, 112, 0, 
    109, 241, 0, 0, 462, 612, 528, 
    232, 0, 481, 569, 626, 576, 637, 
    
    -- channel=50
    340, 278, 302, 161, 288, 188, 330, 
    238, 365, 131, 61, 435, 114, 165, 
    459, 358, 594, 0, 389, 73, 185, 
    304, 254, 507, 230, 371, 108, 419, 
    326, 336, 186, 289, 78, 73, 420, 
    608, 426, 85, 153, 119, 178, 213, 
    268, 165, 133, 151, 130, 178, 88, 
    
    -- channel=51
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 0, 
    0, 0, 0, 0, 54, 77, 69, 
    85, 0, 70, 63, 71, 82, 69, 
    
    -- channel=52
    18, 0, 0, 0, 69, 0, 57, 
    308, 23, 0, 0, 305, 0, 110, 
    285, 123, 41, 0, 561, 0, 59, 
    100, 198, 236, 22, 316, 31, 170, 
    106, 442, 50, 83, 41, 231, 214, 
    440, 547, 135, 202, 272, 325, 288, 
    519, 355, 383, 268, 328, 372, 437, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 69, 36, 8, 
    76, 0, 0, 0, 126, 53, 82, 
    184, 0, 33, 39, 61, 52, 40, 
    289, 179, 82, 152, 46, 185, 85, 
    531, 402, 457, 538, 584, 743, 749, 
    819, 614, 680, 747, 828, 901, 967, 
    
    -- channel=54
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=55
    0, 0, 0, 0, 0, 54, 0, 
    52, 0, 0, 71, 330, 301, 95, 
    637, 0, 229, 302, 477, 397, 270, 
    874, 143, 384, 407, 377, 330, 216, 
    1070, 737, 395, 568, 428, 386, 357, 
    1352, 1266, 1296, 1301, 1215, 1432, 1522, 
    1680, 1599, 1418, 1471, 1596, 1765, 1925, 
    
    -- channel=56
    22, 0, 0, 0, 32, 0, 94, 
    276, 138, 0, 14, 111, 0, 156, 
    49, 220, 83, 0, 281, 105, 0, 
    0, 95, 0, 88, 33, 83, 14, 
    0, 311, 191, 0, 0, 223, 0, 
    88, 0, 268, 0, 120, 25, 0, 
    219, 0, 151, 17, 0, 34, 0, 
    
    -- channel=57
    0, 70, 66, 20, 0, 89, 0, 
    30, 22, 213, 216, 0, 121, 92, 
    0, 24, 0, 334, 0, 210, 103, 
    133, 100, 0, 0, 0, 157, 0, 
    42, 0, 202, 208, 37, 73, 0, 
    0, 0, 79, 0, 17, 5, 0, 
    0, 0, 0, 13, 22, 0, 48, 
    
    -- channel=58
    762, 809, 679, 639, 362, 143, 487, 
    226, 702, 325, 97, 9, 0, 89, 
    0, 521, 34, 0, 0, 0, 0, 
    0, 88, 16, 0, 4, 0, 41, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=59
    565, 640, 653, 450, 290, 376, 392, 
    414, 540, 547, 364, 155, 397, 203, 
    628, 308, 584, 612, 162, 415, 332, 
    658, 483, 384, 474, 270, 335, 349, 
    674, 339, 287, 505, 275, 0, 291, 
    183, 468, 0, 0, 0, 0, 0, 
    0, 160, 0, 0, 0, 0, 0, 
    
    -- channel=60
    28, 36, 21, 0, 7, 0, 15, 
    48, 20, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 16, 
    0, 0, 0, 0, 0, 18, 19, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=61
    66, 30, 100, 0, 83, 27, 79, 
    245, 93, 0, 0, 182, 0, 21, 
    263, 0, 0, 0, 367, 0, 77, 
    144, 110, 102, 5, 181, 0, 113, 
    156, 350, 0, 105, 58, 79, 227, 
    191, 419, 0, 72, 179, 206, 209, 
    182, 174, 199, 158, 189, 190, 268, 
    
    -- channel=62
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 0, 
    0, 25, 0, 0, 0, 40, 0, 
    0, 0, 25, 22, 0, 44, 0, 
    7, 0, 0, 0, 64, 14, 0, 
    82, 0, 221, 174, 75, 93, 109, 
    173, 184, 118, 116, 120, 167, 150, 
    
    -- channel=63
    878, 965, 806, 721, 337, 214, 569, 
    352, 707, 348, 119, 0, 0, 194, 
    0, 394, 0, 0, 0, 0, 0, 
    0, 112, 0, 0, 0, 0, 96, 
    0, 0, 0, 0, 0, 0, 53, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=64
    9, 0, 0, 38, 98, 96, 74, 
    68, 9, 0, 102, 71, 82, 133, 
    4, 0, 0, 46, 34, 146, 166, 
    46, 91, 0, 69, 0, 136, 92, 
    1, 102, 107, 96, 128, 268, 150, 
    195, 0, 280, 235, 351, 372, 374, 
    365, 215, 330, 364, 375, 417, 398, 
    
    -- channel=65
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=66
    0, 8, 234, 87, 25, 0, 0, 
    0, 0, 63, 16, 0, 139, 0, 
    350, 0, 96, 382, 0, 75, 228, 
    613, 125, 288, 158, 150, 93, 65, 
    639, 87, 0, 472, 277, 0, 80, 
    151, 756, 0, 201, 0, 0, 20, 
    0, 1141, 0, 0, 6, 0, 132, 
    
    -- channel=67
    0, 0, 0, 0, 21, 27, 25, 
    50, 0, 0, 31, 0, 32, 59, 
    0, 0, 0, 11, 0, 74, 32, 
    0, 0, 0, 52, 0, 68, 30, 
    0, 39, 84, 0, 0, 131, 0, 
    44, 0, 159, 99, 143, 118, 128, 
    130, 0, 166, 154, 144, 181, 126, 
    
    -- channel=68
    0, 0, 0, 0, 0, 4, 0, 
    31, 0, 126, 145, 0, 93, 0, 
    8, 0, 0, 225, 72, 55, 136, 
    169, 0, 0, 0, 0, 0, 0, 
    91, 134, 183, 244, 0, 69, 47, 
    0, 59, 0, 0, 152, 229, 192, 
    57, 0, 161, 215, 248, 182, 247, 
    
    -- channel=69
    139, 195, 204, 189, 77, 66, 74, 
    0, 88, 128, 78, 0, 81, 0, 
    46, 0, 0, 122, 0, 44, 54, 
    85, 9, 0, 92, 0, 32, 0, 
    114, 0, 0, 37, 61, 0, 0, 
    0, 8, 0, 37, 0, 0, 0, 
    0, 195, 0, 0, 0, 0, 0, 
    
    -- channel=70
    86, 0, 53, 0, 249, 103, 138, 
    293, 236, 155, 114, 685, 209, 206, 
    459, 633, 800, 131, 847, 212, 197, 
    325, 308, 770, 404, 668, 273, 429, 
    515, 750, 419, 304, 199, 290, 280, 
    832, 906, 486, 361, 247, 318, 322, 
    549, 417, 346, 250, 249, 334, 271, 
    
    -- channel=71
    125, 62, 28, 276, 177, 161, 214, 
    0, 0, 0, 0, 112, 101, 222, 
    33, 291, 176, 0, 0, 95, 16, 
    0, 65, 304, 332, 212, 198, 122, 
    8, 0, 0, 0, 249, 217, 88, 
    356, 0, 452, 534, 74, 0, 17, 
    219, 534, 90, 0, 0, 35, 1, 
    
    -- channel=72
    342, 372, 408, 293, 296, 355, 326, 
    302, 303, 334, 273, 298, 349, 224, 
    540, 179, 421, 351, 218, 322, 341, 
    565, 345, 482, 413, 339, 260, 404, 
    612, 275, 252, 492, 299, 78, 433, 
    398, 510, 165, 263, 140, 153, 251, 
    83, 428, 84, 148, 146, 136, 173, 
    
    -- channel=73
    0, 0, 0, 0, 0, 51, 0, 
    198, 8, 165, 105, 165, 83, 23, 
    301, 0, 85, 240, 445, 60, 105, 
    423, 90, 83, 0, 141, 0, 40, 
    422, 511, 394, 437, 42, 26, 205, 
    245, 728, 129, 91, 366, 598, 548, 
    539, 113, 412, 503, 603, 577, 733, 
    
    -- channel=74
    365, 243, 275, 0, 399, 114, 349, 
    650, 584, 57, 0, 764, 0, 142, 
    488, 503, 449, 0, 1078, 0, 87, 
    100, 406, 605, 0, 552, 0, 450, 
    13, 782, 143, 162, 0, 187, 587, 
    627, 718, 0, 0, 30, 248, 186, 
    384, 0, 61, 48, 84, 153, 76, 
    
    -- channel=75
    1383, 1409, 1325, 1395, 702, 498, 967, 
    519, 1157, 758, 396, 290, 356, 367, 
    407, 1281, 963, 368, 103, 489, 94, 
    103, 615, 856, 736, 571, 569, 354, 
    174, 0, 0, 0, 445, 62, 205, 
    98, 188, 315, 0, 0, 0, 0, 
    0, 384, 0, 0, 0, 0, 0, 
    
    -- channel=76
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 37, 103, 175, 81, 
    125, 0, 0, 85, 82, 219, 254, 
    367, 0, 0, 104, 61, 285, 36, 
    493, 246, 0, 242, 310, 467, 128, 
    882, 570, 1227, 1312, 1440, 1659, 1641, 
    1740, 1390, 1693, 1705, 1857, 2010, 2148, 
    
    -- channel=77
    0, 0, 10, 13, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 8, 
    0, 0, 0, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=78
    570, 617, 488, 414, 177, 93, 345, 
    210, 481, 189, 0, 53, 0, 122, 
    0, 465, 0, 0, 16, 0, 0, 
    0, 120, 93, 0, 33, 0, 83, 
    0, 0, 0, 0, 0, 0, 69, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=79
    0, 0, 7, 25, 64, 38, 0, 
    0, 0, 0, 147, 403, 327, 0, 
    772, 111, 788, 471, 536, 470, 248, 
    1017, 205, 781, 602, 560, 464, 216, 
    1284, 740, 176, 620, 448, 221, 224, 
    1336, 1567, 1209, 1070, 757, 813, 860, 
    918, 1716, 949, 854, 913, 1002, 1150, 
    
    -- channel=80
    1265, 1370, 1362, 1043, 685, 669, 928, 
    733, 1148, 881, 504, 455, 533, 396, 
    965, 695, 917, 652, 312, 463, 461, 
    753, 699, 837, 680, 605, 426, 693, 
    859, 330, 263, 657, 433, 0, 771, 
    362, 711, 0, 0, 0, 0, 0, 
    0, 315, 0, 0, 0, 0, 0, 
    
    -- channel=81
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=82
    69, 53, 43, 109, 42, 48, 74, 
    0, 0, 0, 0, 19, 0, 115, 
    0, 187, 0, 0, 0, 8, 0, 
    0, 5, 104, 39, 48, 92, 7, 
    0, 0, 0, 0, 69, 95, 21, 
    57, 0, 186, 169, 66, 40, 47, 
    220, 65, 113, 72, 71, 108, 102, 
    
    -- channel=83
    309, 385, 272, 78, 228, 241, 227, 
    414, 508, 445, 199, 133, 180, 133, 
    250, 111, 268, 260, 148, 130, 227, 
    234, 259, 0, 123, 47, 12, 222, 
    155, 357, 459, 273, 9, 128, 192, 
    0, 0, 0, 0, 69, 68, 75, 
    0, 0, 0, 26, 5, 0, 0, 
    
    -- channel=84
    0, 0, 18, 0, 49, 0, 0, 
    167, 144, 160, 79, 153, 78, 0, 
    288, 0, 201, 272, 439, 73, 197, 
    450, 108, 1, 0, 82, 3, 69, 
    444, 640, 330, 412, 0, 155, 148, 
    371, 576, 69, 160, 463, 589, 564, 
    443, 287, 460, 537, 602, 618, 702, 
    
    -- channel=85
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=86
    242, 210, 340, 157, 232, 0, 141, 
    244, 257, 100, 0, 307, 0, 0, 
    190, 144, 94, 0, 540, 0, 0, 
    41, 129, 383, 0, 326, 0, 105, 
    94, 294, 0, 71, 7, 0, 207, 
    166, 620, 0, 0, 0, 15, 0, 
    0, 281, 0, 0, 0, 0, 50, 
    
    -- channel=87
    0, 0, 0, 0, 0, 0, 0, 
    125, 0, 0, 0, 178, 0, 34, 
    217, 0, 0, 0, 393, 0, 39, 
    89, 4, 52, 2, 211, 56, 71, 
    161, 353, 0, 29, 1, 237, 92, 
    480, 538, 386, 434, 620, 709, 649, 
    803, 604, 818, 688, 801, 876, 961, 
    
    -- channel=88
    204, 195, 192, 124, 223, 232, 256, 
    390, 257, 156, 197, 352, 173, 335, 
    287, 122, 0, 105, 465, 107, 277, 
    136, 221, 132, 65, 296, 100, 323, 
    77, 349, 245, 222, 154, 236, 435, 
    141, 233, 0, 0, 227, 323, 298, 
    329, 0, 226, 245, 267, 276, 252, 
    
    -- channel=89
    1, 26, 199, 263, 0, 182, 43, 
    0, 0, 46, 268, 113, 464, 140, 
    673, 114, 502, 504, 0, 500, 209, 
    811, 135, 681, 642, 481, 561, 243, 
    1076, 81, 7, 496, 498, 0, 173, 
    744, 1109, 879, 750, 297, 245, 383, 
    415, 1316, 430, 362, 384, 400, 574, 
    
    -- channel=90
    232, 176, 135, 158, 275, 178, 329, 
    368, 274, 22, 69, 437, 103, 350, 
    119, 437, 6, 0, 478, 36, 196, 
    0, 249, 309, 155, 389, 160, 342, 
    0, 251, 117, 0, 180, 338, 311, 
    324, 167, 106, 169, 215, 251, 230, 
    444, 68, 279, 207, 220, 309, 229, 
    
    -- channel=91
    37, 29, 133, 0, 179, 36, 0, 
    272, 352, 356, 191, 420, 183, 0, 
    466, 0, 598, 382, 690, 138, 348, 
    603, 248, 216, 113, 241, 51, 304, 
    680, 900, 564, 671, 0, 173, 283, 
    580, 774, 0, 33, 425, 607, 556, 
    284, 149, 418, 511, 556, 539, 583, 
    
    -- channel=92
    16, 0, 0, 58, 0, 41, 107, 
    205, 0, 0, 0, 75, 0, 243, 
    24, 393, 0, 0, 145, 60, 0, 
    0, 94, 80, 11, 134, 50, 0, 
    0, 14, 140, 0, 80, 138, 47, 
    95, 0, 353, 129, 28, 35, 21, 
    429, 0, 98, 9, 20, 79, 37, 
    
    -- channel=93
    1316, 1446, 1436, 946, 612, 455, 802, 
    797, 1413, 1077, 488, 289, 214, 244, 
    373, 896, 695, 513, 467, 153, 218, 
    74, 605, 472, 160, 336, 103, 394, 
    0, 198, 276, 320, 0, 0, 349, 
    0, 41, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=94
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=95
    10, 6, 35, 150, 20, 66, 29, 
    0, 0, 45, 36, 0, 34, 25, 
    0, 88, 0, 6, 0, 63, 0, 
    40, 15, 130, 14, 6, 48, 0, 
    37, 0, 19, 26, 184, 18, 55, 
    74, 71, 178, 197, 37, 53, 107, 
    106, 307, 8, 34, 47, 72, 81, 
    
    -- channel=96
    74, 101, 94, 131, 110, 121, 61, 
    37, 93, 202, 188, 0, 206, 58, 
    85, 56, 225, 284, 0, 217, 119, 
    200, 62, 48, 244, 32, 191, 36, 
    266, 101, 173, 163, 142, 99, 5, 
    92, 93, 242, 167, 143, 46, 87, 
    0, 166, 84, 71, 60, 35, 77, 
    
    -- channel=97
    164, 100, 30, 352, 203, 136, 259, 
    0, 29, 0, 0, 83, 74, 173, 
    0, 374, 195, 0, 0, 72, 0, 
    0, 34, 302, 381, 181, 190, 97, 
    0, 0, 0, 0, 235, 165, 0, 
    294, 0, 617, 570, 6, 0, 0, 
    160, 500, 55, 0, 0, 0, 0, 
    
    -- channel=98
    535, 572, 716, 530, 170, 186, 352, 
    95, 290, 264, 38, 158, 122, 0, 
    643, 430, 684, 153, 77, 114, 0, 
    538, 224, 878, 363, 461, 122, 217, 
    776, 0, 0, 360, 190, 0, 339, 
    574, 1051, 29, 150, 0, 0, 0, 
    0, 763, 0, 0, 0, 0, 0, 
    
    -- channel=99
    289, 248, 287, 54, 234, 170, 322, 
    513, 300, 31, 0, 722, 135, 266, 
    770, 415, 350, 0, 897, 64, 227, 
    488, 350, 817, 230, 769, 79, 567, 
    601, 686, 234, 431, 206, 154, 695, 
    968, 1178, 260, 468, 440, 706, 751, 
    962, 718, 597, 597, 713, 814, 874, 
    
    -- channel=100
    0, 0, 0, 41, 0, 0, 0, 
    0, 0, 17, 176, 0, 90, 171, 
    0, 316, 0, 123, 0, 258, 0, 
    0, 11, 0, 98, 0, 268, 0, 
    0, 0, 221, 0, 0, 158, 0, 
    0, 0, 388, 0, 56, 0, 0, 
    169, 0, 90, 0, 0, 0, 0, 
    
    -- channel=101
    0, 0, 0, 0, 0, 0, 0, 
    253, 281, 370, 168, 0, 0, 0, 
    0, 0, 0, 344, 247, 0, 227, 
    152, 66, 0, 0, 0, 0, 1, 
    0, 490, 503, 432, 0, 78, 40, 
    0, 0, 0, 0, 73, 215, 113, 
    0, 0, 7, 131, 159, 30, 100, 
    
    -- channel=102
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=103
    1500, 1571, 1427, 1293, 769, 725, 1165, 
    854, 1274, 917, 276, 397, 262, 542, 
    529, 1221, 724, 111, 135, 127, 125, 
    37, 626, 869, 497, 598, 175, 581, 
    15, 0, 20, 8, 330, 0, 534, 
    0, 9, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=104
    844, 913, 860, 563, 499, 494, 655, 
    630, 871, 666, 290, 367, 331, 339, 
    593, 447, 554, 358, 288, 215, 361, 
    407, 505, 454, 368, 404, 175, 541, 
    414, 248, 327, 447, 219, 43, 577, 
    112, 299, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=105
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 32, 57, 36, 
    144, 0, 0, 0, 0, 78, 0, 
    272, 117, 0, 70, 126, 244, 0, 
    542, 480, 988, 950, 1067, 1300, 1251, 
    1417, 967, 1317, 1328, 1487, 1595, 1734, 
    
    -- channel=106
    0, 0, 0, 16, 0, 76, 0, 
    0, 0, 0, 196, 0, 129, 123, 
    0, 0, 0, 155, 0, 241, 126, 
    85, 16, 0, 61, 0, 218, 0, 
    45, 51, 115, 80, 173, 224, 26, 
    142, 4, 565, 380, 554, 567, 556, 
    610, 305, 610, 584, 630, 657, 704, 
    
    -- channel=107
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 146, 0, 0, 
    0, 0, 0, 0, 265, 0, 33, 
    68, 0, 27, 0, 79, 52, 0, 
    249, 222, 49, 84, 109, 286, 0, 
    599, 554, 727, 837, 936, 1191, 1101, 
    1336, 828, 1197, 1210, 1355, 1460, 1553, 
    
    -- channel=108
    233, 274, 186, 298, 43, 95, 118, 
    29, 169, 145, 252, 0, 183, 82, 
    0, 94, 4, 340, 0, 318, 90, 
    49, 82, 0, 191, 0, 311, 0, 
    38, 0, 62, 4, 138, 55, 0, 
    0, 0, 418, 36, 94, 0, 0, 
    0, 104, 93, 54, 21, 45, 29, 
    
    -- channel=109
    358, 353, 411, 14, 154, 201, 237, 
    613, 542, 401, 119, 448, 202, 92, 
    970, 296, 700, 401, 796, 204, 228, 
    893, 478, 520, 225, 477, 63, 400, 
    904, 999, 569, 708, 66, 0, 486, 
    769, 1214, 85, 25, 183, 361, 380, 
    381, 327, 209, 281, 322, 341, 433, 
    
    -- channel=110
    199, 206, 233, 236, 229, 78, 157, 
    46, 121, 48, 78, 183, 107, 71, 
    124, 281, 195, 34, 132, 116, 78, 
    109, 108, 379, 274, 277, 202, 163, 
    250, 68, 0, 93, 175, 118, 111, 
    338, 383, 375, 354, 171, 134, 187, 
    196, 545, 251, 132, 162, 215, 241, 
    
    -- channel=111
    87, 70, 36, 135, 54, 130, 120, 
    211, 102, 89, 131, 0, 132, 118, 
    188, 0, 6, 201, 0, 184, 94, 
    140, 159, 0, 149, 0, 127, 18, 
    82, 172, 147, 45, 138, 93, 57, 
    52, 0, 212, 48, 94, 8, 32, 
    6, 78, 55, 40, 11, 14, 21, 
    
    -- channel=112
    395, 326, 283, 105, 282, 103, 342, 
    399, 481, 131, 0, 458, 0, 113, 
    327, 502, 514, 0, 523, 0, 14, 
    14, 244, 442, 84, 348, 0, 345, 
    37, 334, 98, 50, 0, 64, 332, 
    488, 321, 0, 0, 0, 0, 0, 
    115, 0, 0, 0, 0, 0, 0, 
    
    -- channel=113
    314, 233, 245, 430, 249, 227, 374, 
    159, 105, 13, 3, 335, 131, 247, 
    370, 612, 475, 0, 209, 188, 3, 
    179, 300, 722, 455, 519, 286, 255, 
    332, 56, 0, 2, 368, 114, 227, 
    670, 591, 623, 600, 43, 0, 31, 
    341, 797, 107, 0, 0, 34, 50, 
    
    -- channel=114
    9, 0, 148, 0, 0, 11, 0, 
    218, 36, 169, 93, 301, 132, 0, 
    609, 136, 467, 423, 756, 180, 108, 
    793, 200, 368, 66, 350, 77, 77, 
    886, 846, 339, 592, 103, 58, 206, 
    726, 1465, 605, 465, 656, 944, 815, 
    918, 757, 837, 902, 1024, 1033, 1241, 
    
    -- channel=115
    0, 0, 6, 0, 7, 0, 0, 
    0, 0, 0, 0, 26, 0, 0, 
    0, 0, 1, 0, 56, 0, 11, 
    0, 0, 22, 0, 1, 0, 15, 
    0, 11, 0, 28, 0, 0, 0, 
    7, 63, 0, 0, 0, 29, 29, 
    0, 24, 0, 2, 23, 17, 35, 
    
    -- channel=116
    229, 299, 384, 52, 145, 258, 112, 
    409, 375, 466, 382, 133, 304, 39, 
    671, 0, 390, 652, 372, 348, 373, 
    852, 347, 84, 172, 114, 168, 223, 
    806, 709, 564, 801, 126, 24, 419, 
    365, 742, 53, 0, 376, 492, 517, 
    147, 172, 280, 398, 424, 356, 495, 
    
    -- channel=117
    27, 49, 126, 29, 30, 55, 15, 
    22, 0, 53, 168, 62, 156, 78, 
    145, 18, 170, 242, 92, 180, 155, 
    167, 55, 109, 134, 92, 206, 114, 
    211, 66, 75, 203, 61, 36, 69, 
    40, 215, 35, 0, 82, 62, 55, 
    0, 86, 68, 66, 67, 27, 53, 
    
    -- channel=118
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 
    0, 0, 0, 10, 0, 37, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 43, 32, 0, 4, 23, 0, 
    0, 0, 74, 0, 95, 79, 65, 
    13, 0, 80, 85, 77, 86, 61, 
    
    -- channel=119
    32, 0, 0, 0, 0, 0, 203, 
    631, 173, 0, 0, 219, 0, 452, 
    108, 629, 0, 0, 586, 184, 0, 
    0, 207, 0, 37, 133, 138, 21, 
    0, 567, 488, 0, 0, 336, 18, 
    156, 0, 498, 0, 147, 58, 0, 
    673, 0, 217, 34, 0, 108, 0, 
    
    -- channel=120
    185, 129, 145, 0, 218, 93, 159, 
    504, 492, 206, 0, 767, 0, 97, 
    471, 470, 476, 0, 1161, 0, 145, 
    298, 311, 556, 0, 487, 0, 407, 
    283, 851, 629, 622, 0, 213, 790, 
    873, 1065, 0, 107, 597, 1112, 977, 
    1109, 0, 623, 800, 963, 1009, 1044, 
    
    -- channel=121
    198, 173, 197, 326, 130, 163, 207, 
    176, 139, 104, 156, 73, 204, 161, 
    340, 167, 184, 258, 61, 335, 129, 
    343, 246, 230, 358, 220, 315, 109, 
    320, 205, 79, 120, 296, 117, 127, 
    310, 269, 417, 257, 28, 0, 13, 
    78, 602, 45, 0, 0, 0, 0, 
    
    -- channel=122
    2168, 2244, 2108, 1741, 1192, 1010, 1653, 
    1414, 2020, 1362, 705, 689, 517, 880, 
    796, 1494, 945, 525, 546, 426, 601, 
    89, 1166, 986, 692, 760, 463, 1028, 
    0, 67, 236, 304, 445, 46, 881, 
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=123
    59, 0, 0, 32, 36, 44, 194, 
    308, 97, 0, 0, 253, 0, 209, 
    185, 322, 0, 0, 332, 26, 0, 
    0, 123, 162, 57, 262, 13, 92, 
    0, 263, 204, 0, 72, 165, 146, 
    312, 39, 193, 140, 43, 63, 92, 
    378, 20, 88, 9, 0, 94, 0, 
    
    -- channel=124
    0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 14, 0, 0, 
    54, 0, 0, 0, 0, 0, 0, 
    176, 56, 0, 12, 48, 191, 0, 
    513, 305, 526, 708, 728, 890, 885, 
    962, 730, 858, 888, 990, 1080, 1157, 
    
    -- channel=125
    362, 427, 448, 87, 245, 224, 262, 
    382, 506, 382, 137, 374, 203, 49, 
    558, 49, 433, 303, 435, 90, 330, 
    548, 304, 359, 154, 330, 0, 426, 
    611, 526, 280, 562, 104, 0, 453, 
    348, 680, 0, 0, 83, 221, 264, 
    0, 220, 0, 113, 147, 116, 186, 
    
    -- channel=126
    201, 240, 252, 442, 13, 147, 152, 
    0, 0, 0, 195, 0, 309, 139, 
    355, 95, 274, 401, 0, 470, 61, 
    438, 106, 203, 585, 73, 541, 4, 
    565, 0, 0, 67, 338, 6, 0, 
    289, 243, 943, 562, 130, 0, 0, 
    102, 879, 226, 53, 16, 49, 162, 
    
    -- channel=127
    0, 31, 0, 100, 0, 35, 0, 
    0, 0, 32, 146, 0, 139, 52, 
    0, 43, 0, 220, 0, 246, 27, 
    56, 30, 0, 92, 0, 224, 0, 
    47, 0, 79, 40, 140, 3, 0, 
    0, 0, 217, 62, 49, 0, 23, 
    0, 186, 16, 21, 7, 24, 11, 
    
    
    others => 0);
end ifmap_package;
