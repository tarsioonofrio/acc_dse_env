library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    68, 68, 63, 65, 63, 66, 66, 68, 65, 67, 57, 53, 46, 46, 45, 
    55, 64, 67, 68, 69, 63, 54, 65, 61, 39, 19, 22, 40, 50, 46, 
    66, 66, 72, 67, 80, 134, 56, 33, 20, 58, 56, 18, 10, 33, 45, 
    2, 28, 68, 69, 64, 51, 49, 22, 21, 94, 43, 56, 19, 0, 44, 
    19, 63, 52, 80, 59, 51, 58, 21, 21, 47, 60, 19, 20, 0, 17, 
    78, 103, 50, 114, 178, 101, 67, 31, 0, 99, 85, 28, 41, 8, 0, 
    57, 102, 65, 44, 103, 104, 127, 51, 19, 124, 70, 27, 29, 40, 18, 
    85, 76, 27, 36, 77, 163, 77, 82, 34, 120, 77, 36, 44, 60, 24, 
    102, 121, 44, 70, 64, 94, 61, 54, 38, 60, 114, 20, 33, 36, 55, 
    133, 130, 45, 79, 63, 29, 48, 62, 54, 73, 12, 0, 9, 54, 59, 
    144, 124, 59, 124, 31, 39, 109, 109, 25, 0, 0, 0, 24, 60, 57, 
    140, 125, 72, 190, 185, 80, 76, 71, 39, 32, 30, 36, 36, 42, 37, 
    29, 115, 112, 205, 57, 26, 26, 24, 24, 24, 26, 34, 46, 47, 38, 
    29, 27, 149, 130, 42, 32, 21, 26, 26, 31, 42, 54, 35, 54, 75, 
    28, 30, 50, 79, 38, 50, 47, 24, 29, 31, 35, 29, 44, 54, 6, 
    
    -- channel=2
    1, 0, 0, 0, 0, 0, 0, 0, 0, 11, 24, 19, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 9, 40, 14, 0, 14, 47, 23, 0, 
    34, 46, 0, 0, 0, 68, 50, 68, 11, 0, 0, 0, 0, 42, 2, 
    0, 0, 0, 0, 0, 3, 0, 0, 0, 15, 0, 14, 14, 5, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 25, 
    11, 0, 0, 27, 108, 27, 0, 0, 0, 0, 0, 21, 0, 0, 0, 
    0, 0, 60, 0, 9, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 8, 42, 7, 0, 1, 19, 6, 0, 0, 
    0, 0, 0, 0, 0, 82, 38, 0, 0, 8, 77, 54, 35, 0, 0, 
    3, 0, 0, 0, 3, 0, 0, 0, 0, 43, 30, 23, 0, 0, 2, 
    14, 0, 3, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 43, 49, 
    96, 35, 0, 0, 82, 142, 102, 103, 47, 13, 0, 3, 0, 0, 0, 
    0, 78, 20, 0, 108, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 72, 60, 15, 0, 0, 0, 0, 0, 0, 18, 5, 0, 22, 
    0, 0, 15, 107, 32, 37, 22, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 1, 
    4, 3, 0, 0, 0, 54, 5, 0, 0, 20, 34, 17, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 4, 12, 5, 0, 0, 0, 0, 0, 
    23, 45, 0, 4, 9, 24, 18, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 14, 0, 14, 52, 13, 0, 0, 0, 12, 4, 0, 0, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 15, 4, 0, 0, 0, 0, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 6, 15, 0, 0, 0, 0, 2, 0, 0, 
    0, 0, 0, 8, 45, 14, 0, 0, 0, 19, 34, 26, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=4
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 34, 20, 11, 0, 0, 
    2, 0, 0, 0, 0, 0, 0, 8, 17, 16, 7, 16, 18, 20, 0, 
    7, 15, 0, 0, 0, 0, 8, 16, 28, 0, 8, 8, 18, 14, 3, 
    34, 33, 0, 0, 27, 0, 1, 9, 24, 11, 14, 14, 21, 15, 13, 
    28, 43, 0, 0, 0, 0, 7, 0, 21, 23, 16, 23, 24, 20, 21, 
    26, 33, 2, 0, 0, 13, 18, 18, 15, 22, 12, 30, 26, 23, 0, 
    36, 44, 37, 9, 0, 11, 11, 17, 5, 0, 26, 17, 26, 0, 0, 
    34, 47, 38, 33, 28, 1, 0, 15, 35, 2, 6, 16, 11, 0, 0, 
    37, 31, 40, 37, 5, 27, 27, 32, 23, 16, 46, 46, 54, 31, 22, 
    109, 45, 24, 30, 59, 81, 92, 92, 91, 85, 97, 103, 114, 116, 114, 
    129, 105, 32, 54, 75, 96, 98, 97, 99, 105, 111, 117, 115, 110, 121, 
    137, 116, 95, 69, 78, 101, 100, 103, 101, 110, 122, 129, 122, 137, 142, 
    135, 131, 113, 109, 100, 111, 105, 97, 99, 111, 122, 119, 116, 140, 128, 
    
    -- channel=5
    55, 63, 62, 60, 56, 58, 65, 67, 57, 53, 57, 60, 58, 50, 46, 
    55, 62, 65, 64, 61, 45, 47, 64, 57, 11, 0, 0, 16, 46, 52, 
    55, 76, 62, 62, 57, 46, 23, 0, 0, 0, 0, 0, 0, 7, 47, 
    0, 4, 46, 60, 50, 33, 6, 3, 0, 11, 6, 0, 0, 0, 28, 
    0, 0, 41, 54, 52, 31, 8, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 47, 27, 20, 29, 2, 0, 0, 4, 13, 0, 0, 0, 0, 
    0, 0, 28, 46, 21, 11, 22, 11, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 25, 10, 43, 39, 3, 7, 4, 0, 0, 0, 11, 19, 
    0, 0, 0, 0, 6, 0, 0, 0, 2, 0, 0, 12, 0, 1, 28, 
    2, 0, 0, 0, 0, 26, 5, 0, 0, 36, 19, 0, 5, 34, 47, 
    0, 0, 0, 0, 0, 0, 27, 30, 17, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=6
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 20, 35, 20, 6, 0, 0, 
    16, 0, 0, 0, 0, 0, 0, 23, 12, 23, 0, 9, 9, 0, 0, 
    64, 11, 0, 0, 21, 11, 7, 9, 4, 7, 21, 17, 13, 14, 0, 
    70, 16, 0, 0, 0, 6, 0, 16, 5, 31, 17, 12, 21, 23, 12, 
    71, 14, 0, 0, 0, 0, 28, 8, 25, 23, 23, 20, 13, 30, 8, 
    65, 45, 15, 0, 4, 45, 2, 0, 5, 0, 5, 13, 28, 3, 0, 
    68, 64, 40, 13, 0, 0, 0, 9, 15, 0, 18, 0, 0, 0, 0, 
    41, 54, 43, 38, 53, 5, 12, 39, 15, 6, 0, 30, 18, 0, 0, 
    55, 51, 37, 71, 65, 97, 79, 66, 61, 36, 80, 96, 88, 59, 67, 
    115, 70, 70, 48, 65, 78, 82, 85, 104, 113, 121, 125, 133, 131, 139, 
    142, 100, 66, 49, 92, 116, 117, 109, 116, 127, 138, 146, 142, 148, 156, 
    160, 135, 112, 54, 110, 120, 118, 120, 125, 134, 140, 146, 144, 172, 143, 
    152, 150, 113, 97, 108, 118, 122, 119, 126, 130, 138, 135, 155, 164, 148, 
    
    -- channel=7
    40, 42, 46, 45, 43, 41, 47, 49, 43, 27, 22, 26, 36, 41, 37, 
    44, 44, 43, 45, 40, 63, 53, 34, 17, 18, 25, 20, 16, 20, 32, 
    23, 12, 45, 49, 42, 12, 51, 20, 10, 3, 27, 27, 22, 0, 22, 
    41, 4, 41, 42, 46, 27, 31, 22, 13, 0, 55, 14, 25, 13, 0, 
    58, 15, 56, 9, 53, 54, 56, 45, 15, 0, 40, 42, 14, 21, 0, 
    55, 37, 73, 44, 14, 64, 79, 38, 36, 0, 64, 48, 2, 19, 23, 
    71, 47, 37, 52, 0, 45, 32, 60, 33, 0, 64, 40, 15, 12, 29, 
    74, 52, 42, 35, 0, 0, 69, 29, 36, 0, 56, 39, 0, 12, 43, 
    76, 37, 78, 18, 44, 18, 40, 26, 11, 36, 0, 33, 0, 23, 33, 
    57, 42, 72, 5, 30, 32, 29, 38, 30, 11, 21, 0, 0, 20, 37, 
    7, 46, 67, 1, 110, 28, 0, 25, 41, 20, 0, 0, 0, 0, 0, 
    0, 16, 47, 13, 57, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 23, 42, 58, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 43, 11, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=8
    0, 0, 0, 0, 0, 0, 0, 0, 5, 2, 3, 0, 0, 1, 7, 
    0, 0, 0, 0, 0, 0, 31, 0, 24, 0, 10, 1, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 61, 32, 3, 0, 8, 20, 28, 0, 0, 
    87, 0, 0, 0, 8, 0, 0, 34, 4, 0, 53, 0, 41, 23, 0, 
    120, 0, 49, 0, 0, 19, 43, 48, 12, 0, 1, 64, 0, 40, 0, 
    114, 0, 74, 9, 0, 45, 26, 38, 45, 0, 68, 94, 0, 30, 31, 
    131, 0, 13, 54, 0, 0, 0, 56, 59, 0, 93, 53, 0, 0, 22, 
    90, 10, 55, 20, 0, 0, 103, 3, 44, 0, 50, 56, 0, 0, 23, 
    70, 0, 135, 0, 40, 0, 26, 0, 0, 9, 0, 82, 0, 0, 0, 
    3, 0, 114, 0, 42, 33, 0, 0, 10, 12, 67, 11, 0, 0, 11, 
    0, 0, 99, 0, 107, 25, 0, 5, 91, 54, 0, 0, 0, 0, 20, 
    0, 0, 47, 0, 99, 101, 0, 0, 19, 0, 0, 0, 0, 0, 3, 
    12, 0, 0, 0, 194, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 0, 0, 37, 57, 0, 12, 0, 0, 0, 0, 0, 6, 0, 0, 
    36, 0, 0, 0, 14, 0, 0, 2, 0, 0, 3, 0, 0, 0, 58, 
    
    -- channel=9
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 0, 0, 0, 4, 4, 2, 2, 0, 0, 
    0, 4, 0, 0, 0, 41, 0, 0, 0, 62, 30, 21, 1, 0, 5, 
    0, 29, 0, 0, 0, 8, 15, 0, 6, 73, 13, 20, 0, 0, 31, 
    5, 73, 0, 39, 58, 63, 34, 0, 0, 60, 43, 0, 12, 0, 5, 
    27, 73, 0, 7, 103, 59, 37, 17, 0, 107, 34, 0, 26, 3, 0, 
    27, 66, 7, 0, 78, 61, 67, 24, 0, 128, 22, 0, 18, 25, 1, 
    43, 72, 17, 0, 48, 106, 32, 39, 0, 97, 24, 0, 29, 31, 3, 
    62, 99, 0, 55, 1, 58, 17, 14, 33, 34, 22, 0, 15, 25, 12, 
    73, 93, 6, 99, 16, 15, 52, 51, 24, 6, 0, 0, 24, 27, 0, 
    105, 84, 20, 136, 40, 30, 89, 71, 1, 0, 3, 17, 36, 37, 10, 
    109, 98, 58, 170, 57, 8, 50, 46, 20, 28, 34, 45, 47, 51, 38, 
    35, 93, 100, 110, 0, 37, 38, 35, 30, 32, 44, 48, 52, 52, 60, 
    34, 46, 125, 52, 8, 47, 33, 36, 41, 45, 48, 50, 44, 56, 57, 
    37, 50, 53, 56, 19, 36, 38, 37, 49, 51, 40, 46, 73, 65, 22, 
    
    -- channel=10
    11, 13, 5, 7, 9, 0, 10, 14, 9, 20, 27, 18, 6, 4, 10, 
    2, 0, 5, 12, 2, 0, 0, 14, 53, 0, 0, 0, 0, 6, 7, 
    40, 38, 5, 8, 9, 57, 24, 0, 0, 0, 0, 0, 7, 0, 7, 
    0, 0, 0, 0, 4, 0, 0, 0, 3, 0, 13, 4, 9, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 28, 16, 0, 0, 0, 0, 0, 14, 12, 0, 0, 0, 
    0, 21, 0, 26, 8, 0, 14, 0, 5, 0, 5, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 69, 32, 0, 0, 14, 0, 0, 10, 6, 
    0, 0, 0, 0, 0, 29, 0, 0, 0, 8, 0, 59, 0, 0, 0, 
    0, 0, 3, 0, 0, 0, 0, 0, 0, 50, 72, 0, 0, 0, 13, 
    0, 0, 8, 0, 0, 0, 0, 49, 31, 0, 0, 0, 0, 0, 0, 
    14, 2, 0, 0, 93, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 23, 40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 101, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 39, 
    0, 0, 0, 17, 4, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=11
    50, 54, 54, 57, 56, 54, 53, 53, 50, 41, 36, 37, 46, 44, 41, 
    53, 52, 55, 58, 59, 91, 61, 43, 28, 42, 53, 33, 24, 33, 44, 
    31, 38, 52, 56, 52, 56, 45, 28, 21, 64, 69, 69, 45, 17, 40, 
    58, 46, 53, 55, 52, 58, 68, 46, 45, 45, 79, 38, 38, 14, 23, 
    104, 94, 71, 73, 142, 109, 87, 51, 31, 43, 88, 58, 46, 38, 7, 
    90, 105, 81, 28, 66, 83, 104, 71, 50, 55, 103, 58, 45, 53, 36, 
    102, 95, 52, 46, 49, 83, 104, 93, 61, 72, 95, 55, 44, 52, 53, 
    106, 120, 74, 70, 52, 91, 112, 60, 57, 66, 86, 53, 38, 51, 57, 
    127, 116, 80, 70, 59, 52, 57, 55, 63, 67, 21, 38, 22, 50, 55, 
    119, 116, 99, 78, 66, 51, 78, 101, 58, 37, 39, 10, 35, 55, 57, 
    95, 111, 99, 108, 172, 93, 87, 98, 75, 49, 31, 42, 46, 60, 51, 
    54, 102, 118, 143, 110, 48, 37, 36, 40, 43, 48, 53, 62, 64, 61, 
    67, 47, 102, 129, 85, 54, 50, 47, 48, 50, 61, 65, 64, 64, 84, 
    68, 54, 49, 115, 60, 60, 59, 47, 49, 56, 60, 57, 62, 65, 64, 
    73, 57, 46, 53, 42, 35, 47, 58, 62, 71, 60, 60, 83, 97, 67, 
    
    -- channel=12
    61, 56, 61, 65, 66, 60, 61, 64, 65, 56, 42, 39, 49, 54, 52, 
    66, 59, 63, 65, 67, 97, 78, 47, 34, 48, 70, 50, 33, 38, 51, 
    34, 35, 61, 65, 66, 76, 53, 44, 31, 75, 82, 72, 67, 29, 39, 
    79, 60, 67, 67, 60, 67, 83, 58, 57, 58, 86, 55, 47, 30, 31, 
    118, 118, 82, 81, 134, 120, 92, 57, 43, 56, 106, 75, 56, 51, 24, 
    107, 112, 81, 53, 62, 82, 112, 86, 68, 65, 113, 64, 55, 63, 48, 
    112, 124, 54, 51, 71, 92, 115, 99, 73, 91, 108, 70, 62, 67, 66, 
    118, 126, 100, 76, 84, 90, 103, 69, 57, 83, 96, 69, 50, 58, 60, 
    139, 127, 97, 76, 74, 69, 74, 73, 72, 103, 37, 37, 28, 54, 64, 
    125, 132, 109, 103, 73, 53, 84, 120, 79, 29, 43, 21, 48, 72, 72, 
    108, 126, 115, 115, 190, 116, 93, 92, 74, 66, 52, 60, 71, 72, 64, 
    76, 98, 124, 174, 143, 61, 63, 56, 56, 59, 68, 74, 80, 91, 82, 
    99, 70, 103, 154, 83, 70, 70, 67, 72, 74, 86, 89, 89, 86, 104, 
    94, 80, 66, 113, 74, 82, 83, 68, 67, 75, 85, 80, 87, 87, 89, 
    95, 78, 79, 73, 68, 56, 62, 71, 83, 96, 87, 84, 106, 128, 94, 
    
    -- channel=13
    92, 92, 97, 100, 98, 90, 98, 102, 102, 89, 73, 70, 78, 87, 91, 
    95, 95, 99, 102, 97, 106, 103, 93, 65, 48, 54, 47, 43, 64, 89, 
    86, 53, 100, 102, 102, 52, 67, 39, 46, 23, 43, 32, 44, 34, 61, 
    79, 41, 92, 97, 103, 62, 73, 55, 36, 3, 49, 32, 33, 39, 22, 
    57, 46, 93, 62, 99, 72, 53, 53, 32, 0, 47, 61, 37, 46, 27, 
    38, 25, 90, 83, 0, 31, 65, 50, 56, 6, 58, 42, 24, 37, 42, 
    39, 34, 45, 100, 15, 46, 47, 53, 51, 0, 45, 46, 25, 31, 50, 
    44, 25, 45, 73, 43, 37, 47, 20, 45, 16, 42, 40, 17, 31, 46, 
    41, 14, 59, 19, 74, 0, 32, 49, 25, 41, 34, 28, 14, 36, 82, 
    27, 16, 53, 0, 51, 39, 16, 56, 43, 39, 27, 15, 24, 60, 81, 
    0, 23, 40, 3, 88, 72, 28, 14, 38, 24, 18, 21, 6, 7, 26, 
    0, 0, 31, 19, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 40, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 10, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=14
    100, 109, 109, 104, 105, 105, 110, 115, 104, 83, 78, 89, 92, 93, 88, 
    106, 112, 113, 108, 106, 120, 80, 97, 73, 57, 31, 39, 65, 80, 87, 
    79, 102, 109, 112, 112, 110, 61, 38, 26, 57, 11, 17, 18, 49, 92, 
    0, 98, 92, 110, 97, 71, 40, 15, 26, 55, 26, 31, 14, 22, 87, 
    0, 62, 65, 84, 54, 49, 27, 18, 26, 67, 23, 5, 28, 8, 59, 
    0, 51, 57, 104, 98, 37, 35, 11, 11, 99, 13, 0, 28, 10, 16, 
    0, 39, 54, 62, 102, 72, 30, 23, 0, 101, 0, 5, 30, 23, 15, 
    0, 6, 12, 39, 58, 63, 16, 35, 15, 96, 24, 4, 30, 40, 54, 
    0, 16, 0, 50, 34, 48, 25, 32, 35, 60, 34, 15, 47, 65, 87, 
    26, 20, 0, 53, 0, 38, 47, 16, 27, 27, 15, 8, 47, 90, 76, 
    50, 18, 0, 69, 0, 0, 35, 2, 0, 0, 0, 0, 0, 3, 0, 
    0, 19, 0, 87, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 31, 33, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=15
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 2, 0, 16, 0, 12, 3, 0, 0, 0, 
    13, 0, 0, 0, 0, 24, 25, 6, 0, 0, 39, 14, 22, 0, 0, 
    60, 0, 0, 0, 0, 0, 23, 5, 0, 0, 50, 17, 16, 0, 0, 
    80, 12, 9, 0, 59, 23, 70, 24, 10, 0, 45, 35, 0, 8, 0, 
    66, 62, 23, 0, 67, 59, 77, 35, 29, 0, 80, 46, 2, 8, 0, 
    52, 103, 23, 15, 0, 5, 104, 44, 61, 0, 92, 30, 0, 0, 8, 
    65, 101, 25, 26, 0, 48, 84, 43, 31, 0, 62, 41, 0, 10, 0, 
    95, 84, 70, 32, 0, 36, 42, 20, 0, 19, 35, 33, 0, 0, 0, 
    83, 76, 107, 9, 81, 0, 0, 68, 11, 35, 33, 0, 0, 0, 0, 
    59, 75, 108, 0, 111, 48, 32, 104, 81, 13, 0, 0, 14, 32, 43, 
    53, 64, 81, 37, 195, 91, 50, 47, 46, 22, 25, 26, 29, 34, 39, 
    41, 27, 12, 137, 120, 29, 33, 23, 22, 17, 21, 27, 44, 41, 33, 
    57, 33, 0, 167, 45, 23, 32, 27, 24, 27, 32, 44, 40, 26, 72, 
    57, 37, 30, 77, 27, 20, 32, 26, 21, 30, 40, 23, 13, 67, 68, 
    
    -- channel=16
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 4, 0, 6, 45, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 39, 1, 13, 47, 55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 59, 55, 53, 60, 61, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 38, 50, 51, 51, 51, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=17
    181, 182, 182, 182, 183, 183, 183, 182, 182, 183, 181, 182, 183, 182, 183, 
    183, 184, 184, 184, 184, 184, 184, 183, 185, 182, 187, 188, 183, 184, 185, 
    184, 184, 185, 184, 184, 185, 185, 188, 182, 138, 167, 184, 186, 186, 186, 
    184, 181, 189, 187, 185, 181, 190, 153, 126, 107, 101, 176, 188, 189, 189, 
    189, 196, 201, 186, 187, 161, 178, 172, 173, 176, 185, 187, 190, 198, 193, 
    67, 86, 163, 185, 191, 201, 201, 199, 193, 163, 120, 95, 68, 155, 190, 
    156, 174, 176, 131, 139, 36, 56, 76, 156, 185, 189, 182, 174, 174, 191, 
    22, 72, 83, 169, 146, 70, 90, 144, 162, 132, 94, 76, 81, 86, 132, 
    52, 113, 77, 121, 165, 181, 201, 131, 106, 125, 122, 126, 139, 149, 132, 
    131, 145, 155, 152, 148, 137, 116, 99, 109, 72, 90, 60, 53, 63, 80, 
    32, 39, 47, 54, 73, 87, 84, 78, 70, 51, 40, 33, 35, 44, 73, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 46, 48, 80, 
    0, 0, 0, 0, 0, 0, 86, 40, 12, 22, 46, 44, 47, 74, 115, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 50, 72, 99, 137, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 66, 74, 87, 104, 139, 
    
    -- channel=18
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 43, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 63, 42, 22, 10, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 
    180, 162, 35, 0, 0, 0, 0, 0, 0, 0, 17, 81, 126, 86, 0, 
    0, 0, 0, 45, 39, 94, 106, 83, 41, 0, 0, 0, 0, 0, 0, 
    175, 178, 104, 0, 0, 29, 29, 0, 0, 0, 35, 74, 65, 61, 82, 
    20, 0, 22, 49, 15, 0, 0, 0, 95, 99, 56, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 6, 37, 0, 0, 0, 0, 0, 35, 86, 88, 
    0, 120, 124, 129, 116, 101, 73, 60, 56, 40, 52, 51, 13, 3, 3, 
    124, 116, 132, 153, 165, 168, 155, 141, 116, 107, 83, 52, 13, 0, 0, 
    8, 1, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 22, 70, 44, 12, 2, 59, 0, 0, 0, 41, 83, 0, 0, 0, 
    0, 0, 7, 10, 1, 0, 17, 54, 90, 71, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 1, 53, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=19
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 
    0, 0, 0, 0, 0, 0, 19, 68, 0, 0, 0, 0, 0, 0, 0, 
    0, 17, 0, 0, 0, 14, 9, 0, 0, 0, 0, 18, 23, 20, 0, 
    70, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 18, 14, 5, 108, 124, 93, 88, 84, 23, 0, 0, 0, 
    29, 0, 0, 0, 11, 15, 0, 0, 0, 0, 0, 0, 4, 0, 0, 
    8, 21, 18, 20, 21, 22, 8, 9, 0, 40, 67, 9, 0, 0, 0, 
    0, 41, 37, 36, 40, 42, 31, 64, 84, 30, 0, 0, 0, 0, 0, 
    
    -- channel=20
    37, 37, 37, 37, 37, 37, 37, 37, 36, 39, 40, 36, 37, 37, 37, 
    37, 38, 38, 38, 38, 38, 38, 36, 39, 51, 48, 42, 38, 38, 38, 
    36, 37, 37, 38, 38, 39, 38, 47, 55, 61, 56, 36, 38, 37, 38, 
    44, 42, 40, 36, 36, 44, 42, 46, 50, 57, 55, 60, 42, 41, 40, 
    87, 77, 49, 34, 38, 36, 37, 37, 44, 57, 65, 67, 70, 50, 44, 
    37, 32, 49, 40, 47, 54, 51, 47, 39, 51, 55, 47, 45, 52, 46, 
    86, 71, 68, 30, 51, 60, 69, 68, 67, 54, 54, 54, 50, 54, 53, 
    48, 62, 55, 53, 54, 39, 39, 56, 59, 60, 64, 59, 54, 52, 60, 
    41, 44, 20, 22, 38, 48, 59, 45, 48, 58, 59, 65, 65, 71, 72, 
    66, 82, 93, 94, 93, 91, 90, 89, 90, 83, 92, 84, 78, 67, 59, 
    78, 79, 94, 96, 94, 94, 106, 99, 95, 90, 87, 78, 76, 68, 50, 
    26, 35, 23, 30, 30, 36, 35, 75, 80, 76, 66, 64, 40, 35, 30, 
    23, 27, 25, 21, 22, 22, 41, 0, 0, 0, 3, 12, 17, 20, 33, 
    19, 19, 16, 18, 19, 18, 0, 0, 0, 0, 0, 5, 19, 29, 39, 
    20, 13, 18, 20, 17, 19, 1, 0, 0, 0, 9, 19, 23, 29, 39, 
    
    -- channel=21
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 
    3, 1, 0, 0, 8, 26, 47, 44, 25, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 5, 25, 29, 34, 20, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 6, 8, 20, 16, 2, 3, 25, 23, 25, 27, 23, 19, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 0, 0, 0, 0, 0, 38, 101, 104, 86, 52, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 27, 110, 102, 38, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 2, 6, 7, 2, 0, 0, 0, 0, 
    
    -- channel=22
    61, 61, 61, 61, 61, 61, 61, 59, 59, 63, 65, 60, 61, 61, 61, 
    61, 61, 61, 60, 60, 60, 60, 58, 61, 57, 56, 62, 60, 61, 61, 
    59, 60, 59, 59, 60, 61, 64, 60, 69, 78, 74, 60, 60, 60, 61, 
    78, 71, 63, 60, 60, 49, 58, 62, 84, 89, 83, 82, 69, 68, 64, 
    49, 58, 55, 56, 60, 61, 63, 70, 77, 86, 81, 60, 52, 66, 64, 
    106, 95, 59, 55, 51, 75, 64, 67, 70, 69, 88, 92, 77, 80, 69, 
    53, 55, 67, 70, 68, 61, 58, 58, 88, 74, 71, 60, 67, 51, 66, 
    68, 62, 32, 39, 63, 96, 101, 66, 45, 51, 58, 68, 70, 84, 90, 
    86, 89, 94, 90, 88, 73, 83, 99, 99, 110, 105, 98, 84, 62, 63, 
    77, 80, 86, 91, 91, 94, 95, 92, 97, 94, 89, 87, 90, 81, 66, 
    28, 32, 47, 41, 39, 53, 80, 83, 80, 79, 81, 77, 74, 66, 53, 
    14, 39, 29, 20, 17, 28, 57, 75, 71, 71, 65, 74, 49, 26, 45, 
    10, 1, 0, 0, 6, 6, 3, 0, 0, 0, 0, 0, 26, 37, 52, 
    10, 5, 3, 4, 4, 5, 0, 0, 0, 0, 9, 24, 23, 41, 56, 
    6, 0, 5, 5, 4, 8, 0, 0, 0, 6, 11, 22, 35, 44, 59, 
    
    -- channel=23
    68, 65, 65, 65, 65, 65, 65, 67, 67, 65, 64, 65, 65, 65, 65, 
    68, 66, 66, 66, 66, 66, 65, 68, 65, 62, 42, 56, 67, 66, 66, 
    65, 65, 67, 66, 67, 68, 62, 64, 43, 44, 12, 39, 67, 65, 66, 
    55, 64, 61, 66, 69, 73, 49, 72, 57, 58, 58, 33, 60, 62, 63, 
    15, 10, 36, 63, 67, 69, 52, 64, 60, 60, 39, 31, 26, 17, 57, 
    44, 48, 41, 46, 49, 19, 8, 16, 28, 63, 62, 56, 69, 27, 50, 
    10, 2, 20, 48, 50, 70, 13, 34, 26, 43, 37, 34, 24, 26, 20, 
    0, 28, 34, 13, 50, 73, 46, 46, 39, 49, 52, 41, 34, 40, 27, 
    0, 26, 51, 35, 38, 48, 31, 41, 29, 13, 18, 16, 7, 13, 27, 
    0, 11, 6, 13, 19, 22, 27, 31, 17, 30, 7, 16, 6, 4, 14, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 10, 22, 17, 
    0, 0, 12, 10, 0, 0, 3, 41, 23, 23, 26, 25, 19, 36, 22, 
    3, 0, 0, 0, 0, 0, 0, 79, 83, 72, 50, 44, 31, 16, 18, 
    31, 0, 0, 0, 0, 0, 0, 98, 94, 56, 34, 12, 20, 14, 15, 
    28, 0, 0, 0, 0, 0, 0, 20, 31, 12, 19, 17, 14, 17, 21, 
    
    -- channel=24
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 1, 7, 24, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 28, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 0, 0, 0, 5, 12, 0, 27, 0, 0, 
    0, 0, 0, 0, 0, 156, 0, 0, 0, 0, 0, 7, 0, 0, 0, 
    0, 0, 12, 0, 0, 30, 0, 0, 0, 17, 26, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 49, 0, 0, 0, 0, 0, 0, 1, 
    0, 0, 0, 0, 0, 0, 2, 0, 0, 31, 0, 18, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    40, 0, 25, 34, 16, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 
    55, 0, 0, 25, 16, 0, 0, 9, 4, 7, 7, 0, 0, 0, 0, 
    118, 1, 0, 7, 2, 0, 0, 0, 23, 2, 0, 0, 0, 0, 0, 
    115, 14, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=25
    119, 121, 121, 121, 121, 122, 122, 121, 121, 118, 122, 121, 121, 121, 122, 
    121, 122, 122, 121, 122, 121, 122, 121, 116, 96, 122, 127, 122, 122, 123, 
    121, 123, 123, 122, 124, 120, 123, 105, 95, 73, 111, 136, 121, 122, 123, 
    120, 119, 122, 123, 125, 105, 123, 94, 95, 93, 96, 134, 119, 119, 123, 
    83, 97, 126, 124, 122, 107, 127, 113, 122, 106, 98, 92, 87, 125, 123, 
    85, 105, 137, 102, 105, 79, 94, 102, 123, 106, 85, 89, 77, 129, 128, 
    72, 106, 94, 95, 94, 1, 61, 89, 122, 116, 100, 89, 89, 102, 117, 
    68, 67, 63, 122, 99, 63, 102, 100, 94, 79, 59, 60, 75, 80, 94, 
    107, 117, 78, 114, 127, 109, 103, 60, 82, 84, 87, 77, 81, 85, 75, 
    132, 90, 102, 102, 105, 100, 93, 82, 88, 57, 75, 52, 54, 58, 77, 
    8, 31, 29, 32, 37, 50, 60, 62, 53, 48, 41, 48, 64, 56, 73, 
    0, 11, 0, 0, 0, 0, 60, 29, 40, 43, 59, 60, 74, 60, 68, 
    0, 0, 0, 0, 0, 0, 123, 98, 96, 78, 64, 51, 32, 60, 80, 
    0, 0, 0, 0, 0, 0, 39, 102, 58, 33, 22, 44, 43, 58, 87, 
    0, 0, 0, 0, 0, 0, 0, 40, 9, 45, 39, 30, 45, 62, 88, 
    
    -- channel=26
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 14, 2, 3, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    30, 11, 0, 0, 0, 0, 0, 0, 0, 0, 40, 62, 51, 0, 0, 
    0, 0, 0, 6, 10, 89, 107, 88, 43, 0, 0, 0, 0, 0, 0, 
    63, 39, 0, 0, 0, 0, 0, 0, 0, 2, 55, 80, 67, 80, 18, 
    0, 0, 0, 0, 0, 0, 0, 14, 22, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 19, 29, 2, 40, 37, 60, 74, 65, 13, 
    68, 64, 49, 36, 21, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 4, 15, 44, 65, 75, 70, 65, 57, 43, 19, 0, 0, 0, 0, 
    27, 0, 12, 1, 2, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    0, 10, 16, 15, 4, 3, 0, 27, 17, 42, 70, 0, 0, 0, 0, 
    18, 0, 1, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 
    20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=27
    161, 160, 160, 160, 160, 160, 161, 160, 159, 159, 160, 161, 161, 160, 161, 
    161, 160, 160, 160, 160, 160, 160, 160, 156, 136, 130, 149, 160, 160, 160, 
    158, 158, 161, 161, 160, 159, 159, 146, 126, 120, 109, 145, 160, 161, 162, 
    154, 160, 161, 162, 161, 151, 143, 159, 151, 153, 147, 145, 163, 163, 164, 
    67, 79, 136, 157, 158, 166, 156, 163, 161, 154, 133, 114, 93, 119, 162, 
    156, 159, 154, 122, 129, 96, 96, 109, 137, 163, 158, 158, 150, 129, 161, 
    44, 55, 88, 137, 147, 89, 63, 95, 114, 144, 127, 108, 104, 110, 111, 
    36, 88, 89, 85, 138, 154, 159, 135, 99, 94, 89, 88, 101, 118, 118, 
    49, 152, 145, 145, 148, 144, 130, 132, 131, 114, 119, 106, 89, 87, 87, 
    65, 68, 70, 72, 77, 86, 92, 79, 76, 71, 63, 59, 58, 63, 76, 
    0, 0, 0, 0, 0, 0, 0, 6, 16, 14, 15, 26, 49, 62, 74, 
    0, 0, 27, 7, 0, 0, 48, 59, 41, 41, 57, 64, 60, 72, 84, 
    0, 0, 0, 0, 0, 0, 0, 46, 52, 39, 24, 31, 48, 78, 103, 
    25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 57, 76, 85, 113, 
    37, 0, 0, 0, 0, 0, 0, 0, 8, 48, 69, 76, 82, 101, 122, 
    
    -- channel=28
    176, 175, 175, 175, 175, 175, 175, 175, 174, 176, 173, 175, 176, 175, 176, 
    176, 176, 176, 176, 175, 175, 175, 178, 174, 154, 146, 164, 176, 176, 177, 
    171, 172, 176, 177, 176, 174, 174, 166, 143, 128, 123, 153, 176, 177, 178, 
    175, 180, 179, 177, 176, 169, 157, 172, 169, 178, 178, 179, 182, 181, 181, 
    95, 96, 144, 171, 174, 181, 179, 177, 179, 166, 146, 129, 106, 127, 180, 
    161, 169, 181, 138, 135, 105, 87, 101, 139, 180, 179, 178, 172, 159, 181, 
    55, 71, 94, 136, 171, 110, 101, 135, 144, 154, 129, 107, 98, 116, 119, 
    42, 112, 115, 110, 152, 167, 179, 168, 124, 120, 123, 120, 135, 145, 145, 
    59, 164, 152, 155, 159, 159, 142, 123, 126, 115, 110, 105, 89, 100, 99, 
    78, 63, 72, 71, 81, 91, 103, 98, 94, 80, 78, 66, 68, 72, 87, 
    10, 12, 5, 0, 0, 0, 0, 1, 15, 16, 21, 35, 62, 77, 89, 
    0, 5, 23, 17, 0, 0, 58, 101, 75, 66, 74, 70, 66, 78, 103, 
    18, 0, 0, 0, 0, 0, 0, 0, 0, 2, 12, 35, 61, 99, 126, 
    40, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 76, 95, 106, 135, 
    50, 18, 11, 7, 3, 5, 11, 0, 12, 66, 86, 95, 102, 122, 145, 
    
    -- channel=29
    29, 28, 28, 28, 28, 28, 27, 28, 28, 28, 25, 28, 28, 28, 27, 
    28, 27, 27, 27, 26, 27, 26, 27, 30, 26, 0, 15, 27, 27, 26, 
    25, 24, 26, 27, 27, 29, 22, 30, 6, 10, 1, 0, 28, 27, 27, 
    20, 26, 26, 27, 26, 35, 13, 34, 29, 30, 27, 17, 24, 27, 26, 
    0, 0, 0, 22, 26, 30, 29, 30, 29, 33, 18, 0, 0, 0, 21, 
    51, 47, 21, 15, 17, 10, 0, 0, 0, 19, 36, 45, 48, 26, 17, 
    0, 0, 0, 18, 36, 29, 0, 0, 20, 23, 14, 1, 0, 0, 0, 
    0, 42, 3, 0, 6, 60, 59, 34, 0, 0, 0, 10, 13, 25, 32, 
    0, 22, 52, 41, 21, 18, 13, 29, 30, 20, 12, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 6, 
    22, 3, 31, 33, 19, 7, 0, 30, 4, 5, 9, 33, 15, 4, 19, 
    47, 13, 0, 15, 20, 19, 0, 6, 23, 23, 0, 0, 31, 28, 26, 
    66, 23, 18, 21, 22, 22, 0, 0, 16, 14, 48, 48, 33, 27, 20, 
    51, 42, 36, 30, 29, 29, 17, 4, 57, 50, 45, 35, 34, 31, 25, 
    
    -- channel=30
    21, 23, 23, 23, 23, 23, 23, 24, 24, 21, 22, 23, 23, 23, 23, 
    21, 23, 23, 23, 23, 23, 23, 23, 20, 11, 33, 27, 23, 23, 23, 
    23, 25, 25, 23, 25, 22, 21, 13, 2, 0, 22, 39, 21, 23, 23, 
    12, 13, 20, 24, 25, 19, 33, 0, 0, 0, 0, 25, 12, 16, 19, 
    10, 16, 42, 26, 23, 7, 30, 10, 17, 0, 0, 9, 12, 28, 20, 
    0, 13, 35, 17, 30, 0, 20, 20, 23, 2, 0, 0, 0, 41, 19, 
    14, 26, 12, 17, 2, 0, 6, 22, 28, 15, 11, 12, 11, 26, 26, 
    17, 32, 15, 58, 9, 0, 6, 8, 19, 4, 0, 0, 4, 0, 8, 
    72, 5, 0, 19, 23, 10, 8, 0, 0, 0, 0, 0, 2, 10, 2, 
    55, 5, 8, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 
    1, 23, 4, 12, 17, 15, 3, 0, 0, 0, 0, 0, 8, 4, 23, 
    3, 26, 10, 9, 12, 17, 44, 0, 0, 0, 12, 15, 30, 32, 30, 
    0, 36, 40, 22, 17, 24, 122, 107, 116, 98, 84, 58, 28, 31, 31, 
    0, 22, 27, 21, 22, 21, 106, 170, 132, 83, 41, 43, 30, 26, 27, 
    0, 15, 16, 15, 20, 17, 49, 71, 45, 58, 43, 22, 22, 24, 25, 
    
    -- channel=31
    119, 117, 117, 117, 117, 118, 118, 119, 115, 118, 118, 117, 118, 117, 117, 
    120, 118, 118, 119, 118, 118, 117, 119, 120, 141, 101, 110, 119, 118, 118, 
    119, 119, 118, 119, 118, 123, 116, 133, 124, 120, 77, 91, 119, 117, 119, 
    113, 117, 116, 119, 121, 139, 94, 125, 86, 89, 69, 65, 120, 117, 118, 
    96, 86, 93, 116, 120, 131, 94, 121, 104, 122, 128, 117, 113, 78, 114, 
    60, 55, 100, 114, 112, 137, 112, 113, 105, 124, 91, 74, 83, 36, 112, 
    92, 77, 100, 71, 123, 75, 15, 7, 40, 122, 128, 122, 112, 110, 88, 
    0, 3, 43, 42, 95, 72, 39, 103, 101, 97, 76, 51, 37, 51, 52, 
    0, 106, 67, 76, 104, 128, 124, 127, 77, 94, 90, 101, 90, 88, 86, 
    36, 106, 107, 115, 110, 112, 114, 89, 88, 77, 73, 70, 44, 40, 39, 
    4, 0, 26, 23, 25, 32, 61, 62, 64, 60, 42, 28, 19, 28, 25, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 33, 30, 17, 
    0, 0, 0, 0, 0, 0, 0, 85, 67, 65, 52, 28, 7, 11, 24, 
    18, 0, 0, 0, 0, 0, 0, 49, 54, 3, 0, 0, 18, 17, 40, 
    15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 17, 17, 23, 43, 
    
    -- channel=32
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    
    -- channel=33
    119, 125, 159, 166, 172, 170, 183, 176, 187, 194, 187, 193, 182, 189, 185, 
    132, 133, 172, 168, 179, 173, 186, 184, 186, 185, 178, 197, 186, 195, 190, 
    136, 131, 172, 163, 183, 167, 172, 182, 188, 128, 174, 198, 183, 192, 194, 
    131, 116, 161, 160, 168, 165, 151, 139, 140, 94, 101, 155, 194, 177, 181, 
    109, 102, 115, 142, 142, 152, 140, 121, 63, 52, 51, 27, 80, 104, 125, 
    30, 41, 39, 32, 53, 60, 77, 59, 52, 44, 43, 75, 64, 109, 45, 
    52, 47, 39, 63, 93, 70, 69, 44, 48, 62, 104, 145, 91, 106, 28, 
    40, 32, 37, 61, 89, 106, 111, 112, 120, 104, 117, 128, 113, 18, 9, 
    86, 86, 107, 121, 126, 130, 126, 105, 104, 57, 78, 105, 108, 94, 108, 
    33, 60, 86, 106, 96, 97, 104, 117, 112, 113, 111, 113, 107, 82, 67, 
    80, 86, 95, 89, 114, 114, 99, 56, 80, 123, 109, 82, 56, 26, 28, 
    93, 91, 74, 47, 43, 103, 79, 41, 56, 64, 57, 31, 18, 6, 0, 
    76, 84, 66, 49, 61, 62, 40, 37, 43, 34, 16, 15, 0, 0, 0, 
    24, 22, 13, 14, 18, 24, 25, 18, 6, 4, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 32, 0, 0, 0, 0, 0, 0, 
    
    -- channel=34
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 66, 0, 0, 0, 0, 
    0, 2, 0, 0, 0, 0, 0, 42, 33, 27, 47, 23, 7, 6, 0, 
    7, 7, 11, 19, 8, 0, 1, 0, 88, 148, 94, 197, 138, 36, 49, 
    120, 95, 123, 124, 131, 120, 107, 78, 20, 0, 0, 0, 0, 21, 100, 
    0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 10, 30, 0, 20, 0, 0, 0, 0, 0, 0, 4, 0, 27, 45, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 62, 31, 5, 0, 0, 
    11, 42, 49, 3, 5, 28, 36, 16, 0, 0, 0, 0, 3, 0, 27, 
    0, 0, 0, 12, 14, 0, 0, 3, 31, 1, 0, 9, 42, 78, 76, 
    0, 0, 0, 13, 41, 36, 20, 69, 42, 32, 61, 79, 45, 32, 20, 
    8, 15, 16, 43, 3, 3, 25, 0, 12, 41, 34, 34, 24, 17, 25, 
    17, 37, 49, 22, 50, 78, 40, 2, 25, 44, 21, 7, 19, 11, 0, 
    59, 67, 37, 18, 11, 23, 35, 31, 0, 0, 17, 10, 10, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 13, 16, 18, 4, 9, 1, 0, 13, 
    
    -- channel=35
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    3, 0, 0, 0, 14, 0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 26, 2, 0, 0, 0, 0, 0, 
    0, 6, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 95, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 1, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=36
    90, 78, 84, 79, 72, 61, 53, 51, 50, 51, 43, 42, 44, 47, 41, 
    80, 64, 67, 60, 55, 48, 49, 46, 44, 57, 42, 37, 40, 43, 37, 
    64, 50, 49, 41, 41, 35, 45, 45, 43, 54, 54, 37, 37, 36, 34, 
    43, 37, 33, 20, 19, 24, 28, 34, 53, 70, 71, 79, 47, 27, 18, 
    52, 41, 49, 42, 33, 32, 37, 55, 61, 68, 64, 46, 26, 36, 33, 
    57, 51, 51, 43, 46, 54, 66, 76, 63, 60, 48, 25, 29, 18, 33, 
    71, 61, 65, 62, 79, 73, 86, 75, 73, 72, 51, 35, 21, 31, 22, 
    73, 61, 57, 68, 74, 79, 84, 84, 77, 70, 45, 26, 25, 18, 28, 
    94, 78, 89, 89, 95, 92, 90, 78, 66, 45, 32, 33, 40, 39, 31, 
    89, 80, 78, 90, 89, 83, 73, 69, 52, 55, 50, 52, 47, 48, 42, 
    87, 93, 93, 82, 85, 75, 79, 72, 67, 63, 57, 61, 52, 46, 43, 
    91, 90, 92, 82, 76, 83, 68, 52, 56, 64, 59, 54, 58, 49, 42, 
    79, 80, 79, 69, 73, 74, 63, 61, 58, 59, 57, 51, 48, 46, 41, 
    69, 67, 62, 60, 55, 52, 57, 60, 47, 55, 48, 46, 46, 45, 46, 
    38, 40, 46, 46, 49, 48, 52, 49, 45, 52, 44, 44, 45, 43, 40, 
    
    -- channel=37
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 17, 3, 0, 1, 
    5, 6, 24, 31, 22, 13, 5, 0, 0, 0, 0, 0, 2, 30, 33, 
    0, 0, 0, 0, 3, 7, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 10, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=38
    111, 112, 108, 104, 93, 84, 76, 70, 73, 74, 66, 66, 72, 67, 72, 
    91, 92, 85, 79, 66, 64, 60, 61, 68, 51, 60, 63, 64, 60, 61, 
    72, 76, 62, 54, 46, 52, 45, 50, 60, 40, 72, 60, 47, 41, 53, 
    50, 56, 37, 28, 22, 35, 39, 48, 37, 49, 40, 25, 45, 26, 26, 
    37, 34, 27, 23, 16, 26, 43, 62, 81, 78, 74, 66, 37, 0, 17, 
    69, 79, 62, 59, 73, 85, 97, 94, 80, 78, 81, 65, 18, 25, 55, 
    84, 66, 69, 77, 90, 98, 109, 106, 98, 90, 65, 32, 37, 30, 21, 
    108, 94, 121, 123, 120, 119, 119, 105, 93, 54, 28, 33, 42, 31, 36, 
    114, 82, 96, 116, 119, 104, 88, 80, 84, 68, 60, 51, 52, 54, 30, 
    102, 128, 114, 97, 99, 107, 97, 81, 70, 67, 64, 62, 46, 30, 25, 
    108, 114, 109, 98, 88, 81, 69, 55, 66, 68, 51, 44, 48, 42, 34, 
    95, 100, 83, 78, 84, 90, 79, 66, 53, 54, 59, 41, 48, 38, 30, 
    87, 82, 77, 71, 52, 47, 61, 62, 54, 41, 51, 46, 40, 40, 38, 
    37, 42, 46, 53, 48, 44, 45, 42, 62, 50, 39, 40, 40, 40, 36, 
    31, 34, 38, 40, 49, 51, 50, 33, 45, 44, 38, 38, 40, 40, 19, 
    
    -- channel=39
    44, 27, 37, 48, 56, 60, 59, 67, 54, 63, 63, 64, 70, 66, 64, 
    49, 33, 39, 58, 56, 62, 59, 58, 57, 67, 40, 58, 73, 65, 68, 
    53, 34, 41, 64, 54, 62, 59, 38, 42, 78, 0, 37, 71, 59, 58, 
    51, 44, 44, 56, 58, 57, 56, 51, 34, 30, 10, 5, 0, 38, 44, 
    13, 18, 18, 8, 23, 19, 24, 20, 20, 9, 3, 22, 11, 57, 24, 
    0, 0, 16, 11, 18, 13, 8, 16, 9, 10, 10, 34, 74, 10, 35, 
    0, 15, 10, 0, 11, 32, 25, 32, 27, 23, 21, 41, 61, 17, 57, 
    14, 25, 18, 19, 25, 29, 29, 31, 22, 37, 18, 33, 46, 78, 46, 
    6, 8, 10, 20, 23, 20, 24, 31, 24, 46, 23, 36, 40, 42, 17, 
    30, 0, 8, 20, 28, 23, 20, 16, 12, 27, 34, 36, 22, 23, 11, 
    5, 16, 16, 14, 0, 10, 33, 26, 0, 1, 16, 19, 6, 1, 0, 
    0, 13, 25, 14, 9, 0, 13, 11, 4, 6, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    
    -- channel=40
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 5, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 92, 0, 0, 7, 0, 0, 
    16, 4, 0, 0, 0, 0, 0, 0, 31, 47, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 15, 30, 1, 0, 0, 0, 0, 0, 
    0, 0, 6, 0, 0, 0, 0, 16, 0, 0, 0, 0, 52, 0, 79, 
    0, 11, 13, 0, 0, 7, 0, 8, 0, 0, 0, 0, 44, 0, 136, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 1, 120, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 12, 0, 
    26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 32, 6, 
    0, 0, 0, 5, 0, 0, 19, 46, 0, 0, 5, 25, 21, 21, 0, 
    0, 0, 18, 16, 0, 0, 23, 22, 0, 0, 10, 14, 9, 6, 22, 
    0, 0, 11, 1, 0, 0, 4, 0, 0, 1, 13, 0, 26, 2, 6, 
    0, 0, 0, 0, 0, 0, 0, 1, 0, 16, 4, 2, 9, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 6, 0, 64, 0, 4, 0, 0, 22, 
    
    -- channel=41
    93, 107, 131, 128, 131, 126, 129, 118, 132, 130, 123, 129, 120, 129, 131, 
    91, 100, 130, 113, 125, 114, 120, 124, 128, 95, 114, 136, 117, 128, 130, 
    87, 92, 122, 104, 116, 104, 102, 114, 113, 49, 111, 131, 104, 119, 128, 
    80, 78, 106, 108, 104, 103, 93, 69, 61, 36, 63, 60, 102, 100, 109, 
    50, 49, 54, 73, 66, 73, 69, 53, 35, 42, 49, 36, 83, 59, 48, 
    43, 38, 34, 49, 58, 49, 64, 47, 44, 33, 64, 91, 30, 86, 18, 
    59, 32, 33, 68, 81, 65, 75, 63, 61, 65, 93, 100, 56, 61, 0, 
    62, 59, 73, 95, 100, 97, 91, 82, 88, 55, 78, 80, 72, 10, 28, 
    65, 74, 91, 102, 96, 90, 81, 69, 76, 50, 80, 78, 74, 50, 74, 
    51, 71, 94, 89, 76, 76, 76, 67, 71, 80, 82, 65, 51, 27, 27, 
    81, 81, 73, 61, 77, 84, 53, 29, 51, 68, 54, 30, 9, 3, 7, 
    89, 70, 49, 38, 45, 80, 43, 27, 39, 30, 11, 12, 0, 0, 0, 
    61, 50, 37, 32, 36, 31, 18, 18, 16, 15, 0, 8, 0, 0, 0, 
    11, 5, 1, 6, 5, 6, 9, 1, 10, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 25, 0, 0, 0, 0, 0, 0, 
    
    -- channel=42
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 5, 0, 51, 0, 11, 0, 0, 0, 
    20, 0, 11, 7, 9, 0, 1, 4, 50, 0, 0, 0, 13, 39, 21, 
    40, 26, 15, 26, 35, 38, 22, 33, 0, 4, 0, 0, 0, 1, 0, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 51, 
    0, 0, 0, 0, 0, 0, 0, 0, 2, 36, 4, 0, 0, 0, 0, 
    0, 33, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 29, 
    0, 0, 0, 0, 0, 0, 0, 28, 28, 0, 0, 1, 45, 42, 15, 
    0, 0, 0, 19, 35, 11, 10, 0, 0, 20, 49, 29, 23, 16, 29, 
    0, 0, 2, 0, 0, 0, 49, 29, 4, 0, 25, 23, 0, 12, 3, 
    11, 48, 59, 42, 35, 11, 0, 2, 34, 21, 0, 9, 20, 0, 0, 
    16, 11, 8, 4, 20, 27, 10, 0, 0, 8, 7, 1, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 6, 18, 0, 13, 1, 0, 0, 0, 27, 
    
    -- channel=43
    137, 120, 148, 153, 157, 156, 162, 165, 159, 164, 162, 166, 166, 168, 164, 
    138, 118, 146, 150, 156, 149, 148, 157, 157, 142, 120, 160, 164, 164, 160, 
    136, 114, 140, 149, 151, 146, 141, 124, 132, 131, 83, 141, 154, 151, 153, 
    119, 98, 112, 126, 134, 132, 137, 116, 79, 57, 46, 25, 63, 118, 115, 
    44, 38, 45, 43, 54, 58, 70, 80, 71, 65, 60, 71, 85, 91, 46, 
    53, 58, 72, 67, 82, 74, 80, 77, 68, 74, 89, 126, 106, 89, 71, 
    60, 53, 52, 57, 81, 99, 100, 103, 105, 104, 101, 115, 118, 71, 48, 
    86, 94, 100, 114, 120, 126, 127, 116, 108, 91, 74, 89, 102, 95, 76, 
    67, 70, 76, 103, 108, 104, 105, 106, 101, 116, 102, 104, 100, 88, 87, 
    80, 77, 102, 95, 101, 108, 110, 95, 90, 106, 104, 92, 73, 52, 38, 
    87, 96, 89, 79, 69, 93, 91, 57, 48, 72, 70, 58, 40, 36, 19, 
    64, 85, 81, 55, 60, 63, 74, 60, 54, 51, 40, 42, 24, 17, 9, 
    47, 56, 53, 43, 39, 36, 35, 39, 34, 33, 26, 25, 19, 8, 10, 
    6, 5, 13, 17, 23, 23, 25, 23, 34, 36, 18, 9, 9, 10, 9, 
    6, 6, 13, 15, 20, 24, 23, 16, 17, 29, 7, 4, 6, 11, 0, 
    
    -- channel=44
    155, 141, 168, 172, 173, 171, 176, 179, 177, 178, 176, 182, 182, 185, 178, 
    157, 138, 165, 167, 173, 166, 161, 169, 174, 167, 132, 173, 179, 178, 174, 
    153, 130, 157, 165, 169, 161, 157, 139, 143, 149, 97, 150, 165, 164, 166, 
    124, 102, 114, 121, 139, 140, 148, 132, 108, 73, 86, 59, 64, 118, 122, 
    49, 57, 62, 59, 61, 68, 78, 90, 75, 78, 76, 70, 103, 108, 65, 
    70, 74, 85, 83, 107, 98, 95, 87, 85, 91, 103, 142, 133, 101, 94, 
    81, 71, 66, 81, 103, 121, 127, 129, 135, 131, 123, 131, 120, 82, 44, 
    101, 108, 110, 129, 134, 144, 144, 132, 117, 107, 89, 102, 113, 113, 100, 
    77, 84, 92, 118, 122, 119, 128, 132, 124, 127, 121, 120, 114, 96, 95, 
    102, 93, 119, 117, 121, 131, 126, 105, 99, 119, 119, 101, 86, 62, 47, 
    97, 117, 106, 89, 79, 102, 117, 80, 71, 88, 83, 70, 54, 48, 34, 
    88, 105, 106, 79, 86, 84, 74, 64, 74, 69, 57, 61, 40, 33, 20, 
    58, 60, 52, 48, 59, 59, 50, 54, 49, 49, 39, 40, 31, 22, 23, 
    26, 21, 30, 32, 36, 39, 44, 41, 47, 56, 31, 24, 22, 24, 20, 
    19, 23, 32, 36, 39, 41, 41, 28, 34, 42, 21, 15, 20, 24, 12, 
    
    -- channel=45
    7, 0, 0, 3, 8, 12, 18, 26, 17, 22, 19, 23, 27, 25, 20, 
    12, 2, 2, 18, 16, 20, 20, 18, 19, 29, 0, 19, 29, 25, 21, 
    21, 7, 11, 28, 29, 27, 31, 5, 10, 35, 0, 2, 29, 23, 21, 
    20, 15, 18, 14, 28, 27, 28, 44, 0, 0, 0, 0, 0, 17, 9, 
    0, 0, 0, 0, 0, 0, 0, 2, 9, 9, 0, 22, 17, 28, 10, 
    1, 17, 23, 0, 18, 21, 11, 4, 4, 13, 10, 39, 70, 12, 42, 
    0, 5, 0, 0, 0, 3, 1, 7, 20, 21, 19, 16, 34, 31, 36, 
    3, 16, 21, 17, 6, 7, 8, 11, 0, 12, 0, 12, 26, 43, 51, 
    0, 0, 0, 0, 0, 0, 0, 0, 10, 31, 30, 27, 19, 34, 9, 
    0, 6, 0, 0, 0, 8, 14, 13, 0, 7, 13, 23, 10, 6, 1, 
    0, 0, 0, 0, 0, 0, 8, 0, 0, 3, 0, 0, 13, 10, 14, 
    0, 0, 0, 0, 0, 0, 4, 10, 1, 4, 13, 0, 13, 9, 11, 
    0, 0, 0, 0, 0, 0, 0, 13, 4, 0, 14, 8, 10, 9, 13, 
    0, 0, 0, 3, 8, 4, 0, 5, 9, 24, 5, 11, 11, 12, 17, 
    14, 13, 12, 12, 15, 18, 14, 11, 0, 17, 8, 10, 12, 10, 18, 
    
    -- channel=46
    0, 0, 0, 0, 5, 7, 16, 12, 23, 18, 15, 23, 11, 22, 19, 
    0, 0, 15, 3, 21, 16, 26, 26, 22, 10, 26, 32, 15, 26, 29, 
    0, 6, 28, 16, 31, 22, 24, 28, 24, 0, 38, 33, 21, 34, 37, 
    12, 24, 48, 52, 44, 42, 20, 19, 14, 0, 24, 24, 45, 46, 48, 
    19, 22, 23, 41, 39, 39, 23, 0, 0, 0, 0, 0, 41, 47, 39, 
    6, 0, 0, 8, 5, 0, 0, 0, 0, 0, 4, 24, 16, 44, 0, 
    0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 27, 39, 4, 26, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 37, 35, 22, 0, 13, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 25, 22, 15, 7, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 8, 13, 5, 8, 6, 19, 
    0, 0, 0, 0, 0, 4, 0, 0, 8, 8, 5, 0, 0, 0, 8, 
    8, 0, 0, 0, 0, 7, 0, 0, 8, 0, 0, 0, 0, 4, 0, 
    2, 0, 0, 0, 2, 0, 0, 0, 0, 2, 0, 5, 0, 2, 2, 
    7, 0, 0, 0, 0, 3, 1, 0, 0, 0, 3, 3, 0, 4, 6, 
    7, 8, 5, 3, 0, 0, 0, 2, 23, 0, 9, 4, 3, 7, 3, 
    
    -- channel=47
    114, 58, 97, 112, 117, 112, 118, 131, 108, 124, 123, 118, 122, 127, 114, 
    114, 59, 93, 111, 112, 110, 119, 123, 111, 151, 75, 113, 124, 130, 108, 
    114, 55, 83, 104, 108, 104, 121, 103, 92, 157, 34, 99, 121, 117, 104, 
    110, 47, 91, 94, 109, 95, 114, 96, 97, 93, 32, 48, 72, 104, 84, 
    67, 46, 63, 59, 77, 76, 78, 104, 57, 44, 29, 7, 9, 71, 44, 
    3, 5, 42, 5, 36, 35, 49, 65, 34, 30, 0, 36, 65, 66, 55, 
    27, 27, 39, 10, 49, 61, 60, 50, 37, 42, 23, 72, 112, 52, 48, 
    40, 36, 41, 45, 70, 79, 84, 83, 83, 95, 43, 61, 74, 68, 4, 
    69, 67, 44, 80, 98, 94, 83, 72, 55, 74, 28, 59, 70, 67, 66, 
    50, 33, 60, 77, 65, 62, 68, 80, 59, 69, 70, 87, 75, 64, 26, 
    45, 65, 69, 79, 64, 58, 93, 54, 0, 64, 71, 62, 37, 14, 14, 
    19, 59, 80, 37, 25, 30, 87, 35, 15, 34, 31, 13, 11, 0, 0, 
    20, 52, 62, 29, 24, 26, 22, 11, 14, 12, 4, 0, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 0, 0, 
    
    -- channel=48
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=49
    132, 133, 102, 115, 120, 125, 124, 123, 120, 125, 129, 126, 129, 143, 150, 
    138, 148, 124, 74, 118, 115, 113, 121, 118, 122, 126, 127, 141, 150, 156, 
    133, 147, 135, 76, 56, 70, 60, 71, 73, 80, 80, 99, 146, 151, 158, 
    126, 140, 92, 52, 81, 80, 67, 79, 87, 79, 88, 91, 131, 153, 157, 
    124, 140, 126, 112, 117, 121, 117, 119, 125, 112, 121, 132, 136, 147, 151, 
    140, 147, 142, 117, 108, 107, 111, 113, 109, 112, 114, 138, 146, 146, 152, 
    151, 100, 83, 158, 165, 139, 144, 146, 143, 141, 144, 144, 148, 151, 156, 
    163, 153, 108, 15, 65, 155, 165, 150, 150, 144, 143, 143, 142, 140, 148, 
    167, 165, 158, 134, 10, 39, 108, 175, 170, 148, 140, 141, 146, 147, 149, 
    166, 165, 161, 163, 19, 21, 24, 23, 53, 100, 158, 180, 166, 147, 144, 
    167, 155, 161, 106, 8, 0, 0, 27, 15, 0, 0, 0, 77, 106, 148, 
    176, 165, 169, 170, 172, 128, 103, 132, 144, 116, 121, 108, 121, 135, 139, 
    61, 46, 39, 37, 40, 32, 33, 57, 64, 68, 69, 79, 83, 79, 81, 
    51, 52, 46, 38, 34, 28, 26, 27, 22, 13, 12, 11, 9, 7, 25, 
    9, 5, 4, 9, 5, 0, 0, 5, 3, 0, 4, 4, 5, 50, 71, 
    
    -- channel=50
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 11, 25, 33, 38, 33, 27, 23, 29, 25, 0, 0, 0, 
    0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 6, 4, 0, 0, 17, 29, 24, 0, 18, 0, 0, 
    0, 0, 0, 0, 8, 16, 14, 7, 8, 14, 9, 1, 0, 0, 0, 
    0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 134, 98, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 110, 49, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 10, 88, 164, 99, 26, 1, 0, 0, 0, 0, 
    0, 0, 0, 2, 46, 46, 23, 0, 30, 137, 204, 167, 84, 12, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    70, 89, 103, 114, 123, 93, 18, 35, 96, 46, 41, 24, 32, 84, 77, 
    0, 0, 0, 0, 0, 0, 0, 1, 28, 39, 46, 59, 65, 66, 82, 
    65, 79, 73, 58, 50, 48, 40, 33, 25, 17, 16, 9, 9, 5, 0, 
    4, 5, 4, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    
    -- channel=51
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 33, 0, 0, 1, 5, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 44, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 91, 137, 129, 107, 90, 105, 124, 122, 58, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 40, 
    0, 0, 0, 0, 0, 20, 15, 16, 19, 19, 0, 0, 23, 1, 0, 
    
    -- channel=52
    50, 62, 61, 51, 49, 49, 48, 47, 47, 49, 49, 48, 45, 43, 45, 
    66, 76, 67, 17, 31, 33, 31, 27, 28, 30, 29, 23, 49, 52, 50, 
    68, 76, 78, 0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 54, 51, 
    68, 76, 52, 0, 4, 13, 0, 1, 12, 8, 5, 10, 26, 60, 59, 
    68, 75, 68, 55, 53, 54, 58, 53, 56, 51, 48, 48, 48, 63, 63, 
    62, 74, 68, 58, 57, 52, 52, 51, 52, 53, 51, 56, 63, 59, 64, 
    55, 61, 64, 82, 60, 56, 63, 64, 62, 61, 61, 60, 61, 62, 60, 
    57, 64, 47, 12, 47, 68, 47, 53, 58, 56, 56, 58, 60, 60, 64, 
    57, 55, 53, 46, 33, 29, 46, 67, 51, 48, 52, 59, 62, 63, 64, 
    49, 48, 50, 60, 36, 30, 21, 15, 26, 58, 76, 65, 46, 46, 56, 
    49, 51, 55, 43, 18, 13, 30, 21, 9, 21, 12, 26, 33, 40, 59, 
    50, 56, 56, 56, 56, 53, 40, 44, 66, 55, 59, 52, 60, 73, 70, 
    34, 43, 44, 39, 38, 36, 39, 50, 58, 60, 60, 65, 67, 67, 66, 
    33, 41, 44, 35, 29, 29, 31, 29, 27, 22, 23, 22, 21, 17, 27, 
    14, 22, 22, 20, 17, 20, 21, 17, 19, 21, 20, 17, 12, 42, 45, 
    
    -- channel=53
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 1, 34, 47, 40, 42, 49, 48, 39, 27, 2, 0, 0, 
    0, 0, 0, 29, 42, 47, 58, 52, 44, 48, 51, 49, 17, 0, 0, 
    0, 0, 0, 11, 3, 1, 0, 8, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 19, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 24, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 39, 28, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 47, 22, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    37, 39, 41, 39, 38, 45, 54, 35, 10, 17, 17, 19, 6, 0, 0, 
    0, 0, 0, 5, 7, 11, 12, 8, 4, 4, 4, 1, 3, 3, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=54
    86, 97, 76, 57, 67, 68, 62, 67, 63, 63, 64, 63, 71, 75, 77, 
    98, 102, 94, 11, 14, 3, 0, 6, 2, 6, 14, 33, 67, 75, 79, 
    93, 106, 73, 19, 11, 26, 7, 17, 32, 32, 26, 33, 65, 84, 83, 
    94, 106, 58, 15, 39, 44, 32, 34, 36, 24, 27, 28, 62, 84, 88, 
    91, 103, 95, 74, 69, 70, 71, 68, 75, 64, 62, 82, 86, 86, 93, 
    86, 101, 85, 85, 97, 97, 96, 94, 97, 93, 89, 90, 86, 82, 91, 
    81, 77, 43, 47, 72, 75, 87, 90, 88, 86, 86, 87, 86, 84, 87, 
    81, 91, 87, 52, 44, 50, 65, 72, 80, 82, 82, 86, 87, 87, 95, 
    75, 81, 76, 72, 41, 13, 6, 35, 53, 60, 76, 84, 86, 86, 93, 
    69, 74, 76, 64, 16, 17, 15, 14, 3, 4, 29, 40, 53, 66, 84, 
    74, 74, 77, 56, 74, 43, 34, 68, 62, 55, 54, 39, 75, 65, 80, 
    67, 57, 53, 50, 49, 65, 68, 59, 71, 87, 78, 91, 78, 83, 85, 
    55, 55, 58, 52, 47, 50, 55, 52, 49, 48, 44, 45, 45, 40, 38, 
    14, 8, 11, 6, 2, 10, 12, 10, 10, 8, 10, 11, 10, 16, 42, 
    16, 10, 13, 11, 8, 12, 12, 9, 10, 12, 13, 9, 26, 57, 17, 
    
    -- channel=55
    19, 38, 61, 47, 48, 53, 56, 51, 56, 55, 54, 53, 49, 50, 56, 
    21, 32, 57, 94, 60, 65, 73, 65, 72, 68, 70, 59, 60, 58, 55, 
    22, 33, 46, 84, 85, 75, 79, 73, 77, 75, 70, 67, 57, 57, 54, 
    28, 32, 81, 97, 76, 76, 84, 82, 86, 93, 84, 78, 56, 49, 51, 
    43, 35, 45, 56, 44, 40, 44, 46, 46, 49, 41, 39, 54, 52, 52, 
    41, 35, 28, 47, 50, 48, 50, 54, 55, 48, 47, 49, 54, 56, 53, 
    41, 75, 72, 3, 3, 46, 56, 58, 59, 58, 53, 53, 51, 52, 52, 
    37, 55, 59, 92, 26, 0, 18, 58, 61, 59, 54, 54, 53, 54, 49, 
    40, 54, 59, 62, 98, 9, 1, 0, 10, 36, 47, 59, 56, 53, 50, 
    41, 55, 59, 62, 90, 0, 2, 15, 16, 12, 0, 0, 9, 35, 53, 
    35, 60, 58, 79, 83, 88, 39, 20, 61, 62, 48, 50, 11, 48, 49, 
    0, 21, 17, 15, 13, 18, 4, 10, 24, 28, 18, 25, 25, 30, 29, 
    17, 25, 23, 16, 12, 13, 9, 7, 17, 10, 10, 8, 9, 15, 14, 
    20, 14, 14, 11, 9, 7, 8, 7, 6, 5, 1, 0, 1, 3, 0, 
    18, 5, 5, 2, 5, 9, 12, 7, 11, 9, 3, 4, 0, 0, 0, 
    
    -- channel=56
    0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 59, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 6, 18, 0, 0, 9, 0, 0, 1, 0, 0, 0, 0, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 36, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 85, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 3, 191, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 207, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 38, 57, 85, 0, 0, 0, 61, 0, 14, 0, 0, 0, 
    0, 0, 0, 0, 0, 26, 0, 0, 0, 8, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    22, 0, 0, 0, 3, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    36, 1, 0, 0, 2, 0, 0, 0, 2, 0, 1, 0, 0, 0, 0, 
    
    -- channel=57
    107, 123, 89, 96, 111, 106, 100, 102, 101, 104, 103, 102, 110, 119, 117, 
    110, 121, 105, 102, 110, 122, 112, 123, 122, 118, 123, 127, 124, 120, 121, 
    107, 113, 110, 111, 108, 107, 109, 122, 119, 115, 112, 115, 141, 118, 121, 
    104, 114, 105, 90, 102, 109, 91, 113, 107, 102, 107, 107, 123, 115, 120, 
    102, 114, 107, 102, 98, 98, 96, 107, 103, 96, 102, 118, 122, 118, 119, 
    108, 102, 101, 111, 106, 104, 114, 115, 109, 105, 108, 121, 117, 116, 120, 
    113, 90, 49, 85, 109, 124, 125, 125, 120, 115, 119, 115, 117, 118, 121, 
    120, 121, 90, 31, 43, 104, 128, 125, 119, 113, 114, 114, 116, 115, 118, 
    124, 122, 118, 107, 0, 33, 65, 86, 100, 111, 127, 122, 119, 115, 117, 
    123, 121, 118, 96, 0, 14, 20, 25, 36, 44, 74, 80, 99, 116, 122, 
    124, 124, 121, 97, 43, 13, 40, 75, 59, 26, 41, 35, 94, 111, 119, 
    98, 97, 87, 85, 88, 55, 70, 107, 97, 77, 100, 86, 111, 109, 106, 
    45, 57, 49, 44, 39, 34, 42, 62, 50, 51, 51, 55, 57, 55, 54, 
    8, 25, 17, 13, 3, 5, 6, 6, 0, 0, 0, 0, 0, 0, 0, 
    0, 2, 2, 1, 0, 6, 3, 5, 1, 0, 0, 0, 2, 0, 11, 
    
    -- channel=58
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 14, 1, 10, 11, 15, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 21, 33, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 3, 0, 13, 44, 73, 42, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 64, 0, 0, 0, 0, 17, 33, 87, 84, 27, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    75, 89, 100, 104, 105, 94, 82, 63, 43, 27, 33, 19, 23, 6, 9, 
    0, 0, 0, 1, 8, 13, 15, 22, 38, 44, 52, 51, 56, 62, 58, 
    6, 5, 5, 1, 6, 0, 0, 0, 1, 3, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 76, 
    
    -- channel=59
    114, 133, 131, 107, 112, 121, 121, 118, 123, 122, 122, 123, 128, 138, 139, 
    113, 130, 135, 89, 66, 87, 88, 81, 88, 90, 88, 89, 132, 138, 141, 
    110, 126, 132, 82, 92, 75, 75, 76, 89, 90, 94, 97, 116, 139, 141, 
    112, 126, 124, 70, 84, 86, 86, 80, 85, 84, 79, 93, 88, 135, 137, 
    123, 124, 131, 119, 99, 99, 104, 106, 104, 109, 104, 116, 128, 137, 136, 
    133, 123, 114, 134, 137, 135, 136, 138, 136, 137, 138, 131, 133, 135, 137, 
    136, 141, 95, 39, 71, 128, 135, 138, 140, 137, 134, 135, 135, 134, 133, 
    138, 146, 154, 140, 50, 40, 101, 138, 135, 132, 132, 134, 135, 136, 134, 
    139, 147, 148, 150, 93, 28, 26, 31, 72, 110, 129, 138, 135, 134, 134, 
    137, 141, 144, 128, 81, 7, 20, 34, 33, 14, 1, 32, 81, 120, 134, 
    133, 139, 142, 149, 128, 109, 61, 77, 126, 104, 96, 86, 83, 120, 116, 
    81, 80, 77, 72, 68, 72, 73, 77, 81, 77, 86, 87, 90, 81, 81, 
    64, 63, 64, 63, 61, 56, 52, 49, 44, 38, 37, 33, 35, 34, 25, 
    23, 13, 15, 18, 19, 14, 12, 15, 21, 20, 17, 21, 20, 26, 53, 
    27, 23, 21, 21, 22, 29, 29, 32, 37, 33, 27, 24, 41, 57, 61, 
    
    -- channel=60
    127, 139, 142, 116, 125, 136, 139, 135, 140, 140, 139, 136, 137, 146, 152, 
    129, 145, 148, 96, 56, 61, 67, 55, 62, 69, 67, 80, 137, 149, 149, 
    127, 144, 136, 51, 81, 65, 54, 57, 78, 79, 76, 76, 123, 154, 152, 
    130, 141, 149, 63, 92, 93, 99, 90, 98, 95, 94, 109, 97, 149, 151, 
    141, 143, 142, 130, 110, 112, 114, 115, 113, 117, 115, 128, 135, 151, 150, 
    150, 135, 119, 132, 150, 144, 144, 145, 143, 146, 147, 148, 150, 153, 153, 
    154, 163, 137, 66, 62, 128, 148, 151, 151, 149, 145, 146, 147, 146, 146, 
    155, 160, 156, 154, 86, 42, 93, 144, 148, 145, 146, 147, 149, 150, 149, 
    156, 160, 163, 158, 103, 45, 53, 37, 59, 101, 130, 147, 147, 148, 147, 
    155, 156, 158, 135, 80, 22, 25, 40, 59, 47, 18, 28, 66, 114, 140, 
    149, 150, 157, 167, 137, 146, 105, 101, 151, 131, 130, 128, 115, 148, 137, 
    79, 69, 66, 60, 58, 49, 54, 70, 73, 63, 78, 73, 90, 79, 76, 
    75, 62, 60, 57, 55, 51, 48, 48, 44, 37, 37, 34, 34, 35, 31, 
    48, 35, 34, 36, 40, 36, 34, 38, 40, 40, 36, 35, 35, 48, 77, 
    41, 37, 34, 36, 38, 44, 47, 50, 56, 51, 43, 42, 68, 81, 92, 
    
    -- channel=61
    8, 2, 17, 14, 3, 10, 15, 12, 17, 13, 15, 13, 15, 22, 22, 
    5, 0, 6, 0, 6, 0, 0, 0, 0, 2, 0, 0, 9, 9, 13, 
    0, 0, 3, 8, 26, 39, 33, 30, 35, 44, 44, 40, 6, 13, 10, 
    5, 0, 0, 17, 9, 6, 16, 7, 4, 0, 1, 9, 7, 6, 4, 
    13, 0, 3, 13, 6, 2, 4, 3, 7, 5, 7, 0, 17, 8, 7, 
    15, 13, 0, 1, 23, 21, 18, 18, 22, 22, 19, 13, 5, 8, 9, 
    14, 12, 30, 0, 0, 0, 2, 6, 9, 12, 7, 9, 6, 4, 2, 
    12, 10, 31, 78, 32, 0, 0, 1, 8, 8, 9, 10, 8, 8, 6, 
    14, 13, 15, 20, 77, 13, 0, 0, 0, 0, 0, 8, 9, 7, 4, 
    14, 13, 14, 30, 40, 6, 13, 21, 11, 0, 0, 0, 0, 0, 3, 
    9, 10, 13, 14, 57, 84, 28, 28, 68, 56, 55, 45, 24, 18, 6, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    23, 10, 19, 21, 27, 24, 17, 1, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 6, 14, 11, 11, 13, 21, 24, 23, 25, 24, 22, 43, 
    38, 24, 24, 27, 28, 26, 33, 32, 35, 36, 37, 35, 25, 60, 25, 
    
    -- channel=62
    30, 5, 0, 20, 27, 16, 16, 15, 17, 18, 18, 18, 20, 22, 14, 
    21, 1, 0, 34, 84, 90, 78, 84, 82, 84, 72, 53, 43, 18, 15, 
    20, 0, 15, 33, 62, 70, 67, 77, 55, 56, 63, 59, 45, 11, 14, 
    18, 0, 15, 54, 53, 44, 40, 59, 54, 51, 62, 63, 46, 14, 10, 
    15, 1, 0, 3, 14, 12, 11, 18, 14, 11, 19, 20, 14, 9, 5, 
    16, 0, 0, 10, 0, 0, 6, 5, 0, 1, 6, 13, 6, 8, 6, 
    24, 0, 0, 21, 31, 26, 12, 8, 6, 6, 10, 7, 8, 11, 9, 
    29, 7, 0, 0, 9, 49, 41, 24, 12, 7, 10, 7, 7, 5, 4, 
    35, 15, 11, 3, 0, 38, 59, 42, 36, 33, 26, 12, 8, 6, 4, 
    40, 19, 15, 13, 0, 24, 37, 38, 45, 37, 41, 31, 37, 31, 17, 
    40, 16, 15, 1, 0, 0, 20, 27, 12, 0, 14, 9, 36, 32, 16, 
    38, 23, 24, 25, 26, 0, 17, 44, 17, 3, 19, 5, 25, 15, 11, 
    23, 14, 12, 13, 16, 12, 15, 25, 13, 15, 17, 18, 18, 19, 18, 
    25, 27, 24, 27, 24, 25, 23, 24, 19, 19, 21, 23, 24, 17, 4, 
    17, 22, 23, 26, 22, 29, 23, 27, 23, 22, 20, 20, 15, 0, 9, 
    
    -- channel=63
    64, 101, 100, 86, 84, 94, 95, 87, 87, 88, 94, 93, 86, 101, 104, 
    67, 95, 116, 112, 82, 96, 101, 92, 106, 104, 108, 90, 102, 111, 108, 
    67, 93, 111, 109, 104, 84, 90, 83, 98, 103, 86, 75, 102, 109, 107, 
    72, 92, 132, 67, 82, 81, 83, 75, 81, 100, 86, 95, 62, 106, 108, 
    85, 91, 104, 116, 88, 89, 85, 90, 99, 95, 83, 87, 103, 109, 107, 
    94, 106, 101, 96, 94, 90, 93, 101, 100, 94, 90, 94, 108, 106, 104, 
    91, 107, 77, 63, 79, 95, 107, 114, 112, 112, 107, 110, 108, 111, 110, 
    89, 112, 115, 84, 33, 40, 82, 107, 117, 116, 105, 107, 107, 108, 105, 
    91, 110, 114, 121, 117, 0, 5, 60, 86, 97, 97, 113, 112, 108, 106, 
    93, 111, 114, 129, 134, 1, 0, 1, 3, 32, 36, 79, 81, 92, 103, 
    89, 114, 113, 134, 63, 34, 0, 0, 40, 16, 1, 2, 0, 57, 93, 
    87, 114, 110, 108, 104, 114, 74, 70, 114, 105, 95, 102, 97, 114, 112, 
    30, 44, 43, 35, 25, 25, 23, 26, 47, 39, 40, 38, 42, 49, 40, 
    12, 14, 15, 1, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    
    -- channel=64
    0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=65
    23, 0, 27, 35, 0, 11, 27, 33, 76, 78, 51, 69, 36, 38, 27, 
    41, 26, 44, 45, 0, 23, 25, 37, 46, 58, 39, 84, 27, 35, 52, 
    78, 57, 46, 41, 0, 0, 35, 60, 56, 46, 49, 94, 93, 78, 75, 
    14, 44, 50, 12, 0, 77, 94, 10, 64, 0, 69, 133, 129, 94, 71, 
    24, 108, 47, 30, 44, 83, 20, 19, 62, 79, 113, 119, 125, 106, 24, 
    15, 119, 105, 0, 93, 77, 31, 66, 84, 94, 75, 106, 122, 113, 3, 
    11, 82, 127, 101, 69, 60, 46, 74, 77, 70, 50, 86, 103, 115, 12, 
    47, 85, 101, 113, 61, 52, 81, 82, 51, 53, 77, 100, 72, 111, 27, 
    54, 88, 104, 103, 124, 38, 80, 76, 89, 106, 91, 101, 90, 83, 7, 
    98, 88, 72, 96, 86, 130, 67, 92, 99, 95, 86, 87, 51, 47, 59, 
    64, 78, 44, 63, 85, 55, 125, 110, 103, 101, 84, 82, 66, 50, 110, 
    40, 82, 67, 104, 85, 84, 114, 122, 107, 75, 80, 86, 69, 106, 113, 
    150, 187, 132, 115, 90, 121, 105, 111, 114, 81, 103, 64, 62, 85, 125, 
    52, 121, 185, 149, 113, 113, 121, 56, 75, 111, 97, 84, 38, 87, 60, 
    41, 0, 112, 189, 159, 118, 123, 125, 107, 95, 110, 59, 12, 29, 156, 
    
    -- channel=66
    0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 1, 0, 0, 22, 0, 
    0, 0, 0, 0, 2, 4, 25, 0, 0, 0, 0, 0, 0, 0, 0, 
    42, 34, 0, 9, 9, 0, 0, 0, 8, 30, 5, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 52, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 16, 
    6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 14, 0, 0, 0, 0, 0, 20, 0, 0, 0, 3, 0, 0, 
    8, 0, 0, 2, 0, 14, 4, 0, 0, 0, 0, 0, 0, 0, 44, 
    0, 0, 22, 22, 45, 0, 0, 0, 0, 19, 8, 0, 52, 19, 0, 
    0, 35, 27, 18, 3, 77, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 0, 0, 0, 0, 0, 5, 0, 0, 22, 1, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 6, 2, 0, 0, 0, 1, 0, 6, 
    66, 86, 0, 0, 0, 0, 0, 60, 69, 0, 0, 0, 0, 42, 9, 
    0, 110, 99, 0, 0, 0, 7, 0, 0, 6, 0, 15, 49, 8, 0, 
    0, 0, 63, 56, 0, 0, 0, 0, 32, 39, 50, 35, 0, 0, 0, 
    
    -- channel=67
    3, 13, 6, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 20, 0, 
    0, 0, 0, 0, 0, 41, 17, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 38, 0, 0, 21, 0, 0, 0, 0, 8, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 38, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 34, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    35, 35, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 10, 1, 0, 0, 0, 0, 0, 0, 
    0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 47, 47, 0, 
    
    -- channel=68
    20, 16, 25, 37, 36, 23, 18, 19, 24, 16, 27, 16, 19, 17, 19, 
    22, 18, 26, 37, 28, 24, 23, 24, 14, 21, 24, 15, 6, 17, 24, 
    36, 17, 30, 38, 20, 15, 20, 32, 21, 36, 21, 12, 17, 25, 35, 
    29, 17, 34, 24, 14, 20, 27, 15, 37, 8, 25, 15, 23, 25, 42, 
    29, 30, 22, 29, 2, 13, 18, 13, 12, 9, 21, 3, 19, 30, 43, 
    23, 37, 31, 12, 27, 11, 0, 2, 10, 12, 9, 4, 15, 37, 29, 
    16, 32, 34, 29, 2, 0, 0, 2, 7, 0, 0, 0, 8, 33, 20, 
    26, 29, 31, 30, 0, 0, 0, 0, 0, 0, 1, 0, 3, 28, 28, 
    19, 29, 34, 30, 17, 0, 0, 0, 0, 0, 0, 0, 16, 14, 13, 
    35, 26, 30, 33, 5, 22, 0, 0, 0, 0, 0, 0, 0, 26, 25, 
    35, 20, 24, 24, 37, 3, 9, 0, 0, 5, 0, 0, 3, 18, 36, 
    11, 0, 5, 33, 26, 30, 0, 0, 0, 0, 0, 0, 0, 6, 39, 
    36, 11, 0, 4, 18, 23, 3, 0, 0, 0, 0, 0, 0, 13, 42, 
    30, 33, 9, 0, 2, 8, 11, 0, 11, 0, 0, 0, 0, 33, 15, 
    24, 5, 29, 1, 0, 0, 8, 11, 15, 0, 0, 0, 6, 23, 19, 
    
    -- channel=69
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 19, 22, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 17, 24, 12, 0, 1, 22, 26, 6, 0, 0, 0, 
    0, 0, 0, 0, 10, 0, 14, 25, 33, 0, 0, 20, 7, 0, 0, 
    0, 0, 0, 0, 3, 30, 16, 28, 8, 3, 15, 18, 22, 29, 0, 
    0, 0, 0, 0, 0, 4, 35, 11, 20, 20, 14, 13, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 18, 10, 15, 19, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 12, 19, 16, 14, 18, 21, 25, 0, 0, 
    0, 17, 2, 0, 0, 0, 18, 33, 39, 18, 20, 16, 10, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 21, 20, 18, 4, 0, 0, 
    0, 0, 0, 11, 7, 0, 0, 0, 0, 32, 44, 9, 0, 0, 0, 
    
    -- channel=70
    16, 17, 18, 30, 15, 12, 10, 17, 0, 3, 8, 19, 0, 0, 18, 
    21, 24, 23, 31, 16, 0, 9, 14, 18, 17, 2, 15, 0, 33, 15, 
    6, 0, 24, 27, 11, 7, 22, 17, 13, 8, 0, 25, 11, 20, 24, 
    13, 14, 27, 2, 20, 5, 0, 0, 9, 9, 5, 10, 17, 29, 6, 
    23, 26, 22, 20, 11, 6, 0, 23, 9, 13, 0, 2, 11, 32, 6, 
    13, 22, 37, 19, 4, 0, 16, 7, 0, 0, 0, 10, 4, 37, 5, 
    25, 21, 36, 21, 0, 0, 0, 0, 0, 0, 0, 0, 10, 28, 20, 
    13, 24, 26, 21, 0, 0, 0, 0, 0, 0, 0, 10, 0, 18, 6, 
    32, 26, 30, 20, 7, 0, 0, 0, 0, 0, 0, 0, 0, 9, 5, 
    34, 11, 15, 10, 4, 30, 0, 0, 1, 0, 0, 0, 0, 16, 32, 
    7, 12, 14, 24, 22, 0, 14, 0, 0, 0, 0, 0, 0, 29, 38, 
    31, 15, 1, 22, 26, 17, 0, 0, 2, 0, 0, 0, 0, 25, 26, 
    1, 0, 0, 3, 0, 39, 0, 0, 0, 0, 0, 0, 0, 14, 22, 
    0, 0, 0, 0, 0, 0, 0, 7, 9, 0, 0, 0, 0, 15, 0, 
    3, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 13, 5, 13, 
    
    -- channel=71
    0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 
    0, 4, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 40, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 27, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 18, 0, 0, 5, 0, 11, 
    0, 0, 28, 0, 0, 0, 16, 0, 0, 0, 0, 0, 3, 0, 30, 
    11, 0, 0, 43, 0, 10, 27, 0, 7, 0, 3, 0, 9, 0, 35, 
    19, 0, 0, 10, 23, 31, 47, 29, 31, 27, 40, 33, 11, 0, 29, 
    8, 0, 0, 7, 41, 37, 30, 39, 52, 55, 50, 26, 63, 2, 22, 
    0, 0, 0, 0, 0, 85, 25, 45, 55, 51, 47, 41, 41, 8, 29, 
    0, 0, 0, 0, 3, 0, 60, 55, 48, 59, 50, 46, 49, 9, 0, 
    16, 0, 5, 0, 0, 30, 0, 56, 61, 48, 52, 48, 39, 9, 0, 
    21, 19, 32, 0, 0, 0, 22, 49, 52, 60, 51, 48, 40, 0, 0, 
    0, 0, 27, 17, 9, 0, 12, 34, 15, 57, 36, 65, 39, 0, 0, 
    3, 0, 0, 6, 24, 0, 0, 20, 5, 35, 53, 52, 38, 0, 0, 
    0, 0, 0, 0, 6, 23, 1, 0, 4, 14, 16, 39, 34, 0, 0, 
    
    -- channel=72
    0, 42, 0, 0, 66, 0, 0, 0, 0, 0, 33, 0, 90, 0, 4, 
    2, 35, 5, 0, 94, 0, 0, 0, 0, 0, 28, 0, 91, 0, 0, 
    2, 8, 7, 9, 95, 0, 0, 0, 0, 44, 0, 0, 22, 0, 0, 
    36, 0, 8, 35, 36, 0, 4, 89, 0, 73, 0, 0, 0, 0, 33, 
    50, 0, 63, 19, 0, 0, 90, 0, 0, 0, 0, 0, 0, 0, 111, 
    90, 0, 0, 109, 0, 0, 41, 0, 2, 0, 12, 0, 27, 0, 135, 
    74, 0, 0, 7, 21, 0, 12, 0, 0, 0, 0, 0, 21, 0, 129, 
    47, 0, 0, 0, 0, 49, 0, 0, 6, 0, 0, 0, 34, 0, 134, 
    0, 0, 6, 0, 0, 55, 0, 0, 0, 0, 6, 0, 19, 18, 95, 
    0, 26, 40, 0, 0, 0, 10, 0, 0, 0, 7, 2, 45, 0, 0, 
    63, 0, 46, 0, 0, 31, 0, 0, 0, 0, 0, 0, 20, 4, 0, 
    1, 0, 58, 0, 15, 0, 0, 0, 0, 31, 0, 0, 25, 0, 2, 
    0, 0, 23, 31, 34, 0, 0, 16, 0, 1, 0, 34, 22, 0, 0, 
    19, 0, 0, 0, 37, 9, 0, 37, 0, 0, 0, 30, 92, 0, 0, 
    45, 18, 0, 0, 0, 27, 15, 0, 14, 0, 0, 39, 60, 0, 0, 
    
    -- channel=73
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 0, 0, 
    3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 33, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 
    0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 20, 3, 11, 8, 0, 
    0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 13, 0, 
    0, 45, 11, 0, 5, 16, 0, 31, 0, 3, 0, 3, 0, 20, 0, 
    0, 28, 33, 3, 11, 31, 15, 39, 21, 35, 35, 37, 2, 9, 0, 
    0, 15, 9, 13, 43, 18, 47, 35, 43, 43, 39, 69, 17, 8, 0, 
    0, 9, 9, 12, 57, 5, 68, 57, 57, 57, 37, 53, 32, 5, 0, 
    2, 0, 0, 0, 8, 72, 46, 68, 64, 60, 45, 39, 11, 0, 0, 
    0, 0, 0, 17, 0, 0, 87, 74, 63, 53, 51, 42, 16, 6, 9, 
    7, 38, 0, 0, 0, 25, 68, 71, 67, 40, 63, 44, 0, 8, 0, 
    19, 50, 0, 0, 0, 20, 52, 32, 61, 57, 79, 37, 5, 0, 0, 
    0, 0, 32, 4, 0, 0, 0, 0, 36, 69, 53, 29, 0, 0, 0, 
    0, 0, 14, 31, 13, 0, 0, 0, 0, 37, 45, 11, 0, 1, 38, 
    
    -- channel=74
    0, 0, 0, 11, 42, 0, 26, 8, 41, 41, 38, 0, 67, 15, 0, 
    0, 0, 24, 10, 33, 23, 30, 0, 24, 6, 47, 0, 22, 0, 18, 
    48, 47, 6, 22, 26, 0, 0, 34, 38, 41, 8, 0, 18, 0, 4, 
    24, 0, 0, 14, 0, 0, 63, 62, 0, 0, 0, 0, 43, 4, 70, 
    18, 0, 14, 3, 0, 20, 43, 0, 19, 0, 34, 38, 27, 9, 74, 
    39, 10, 18, 0, 0, 0, 0, 13, 16, 21, 22, 0, 44, 21, 60, 
    0, 0, 8, 10, 21, 11, 0, 0, 0, 0, 0, 0, 22, 3, 38, 
    16, 0, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 58, 
    0, 0, 35, 32, 4, 0, 0, 0, 0, 0, 0, 0, 19, 59, 26, 
    5, 52, 27, 20, 45, 0, 0, 0, 0, 0, 0, 0, 16, 0, 0, 
    57, 0, 19, 2, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 16, 17, 32, 
    65, 60, 24, 9, 20, 12, 26, 66, 20, 0, 0, 0, 12, 10, 47, 
    38, 58, 69, 13, 14, 20, 19, 0, 0, 0, 0, 0, 70, 0, 14, 
    58, 22, 20, 70, 26, 1, 13, 15, 21, 34, 67, 18, 0, 0, 0, 
    
    -- channel=75
    51, 38, 38, 50, 33, 13, 47, 38, 56, 60, 61, 58, 74, 25, 43, 
    76, 56, 64, 54, 30, 4, 31, 35, 67, 58, 63, 58, 103, 56, 74, 
    39, 41, 58, 42, 24, 32, 62, 51, 59, 35, 50, 78, 114, 86, 86, 
    47, 58, 60, 46, 33, 63, 71, 44, 29, 68, 72, 84, 113, 100, 77, 
    56, 76, 103, 39, 52, 98, 77, 36, 91, 82, 88, 99, 112, 100, 67, 
    51, 58, 113, 105, 68, 78, 63, 95, 99, 94, 87, 81, 110, 100, 69, 
    59, 64, 87, 115, 86, 73, 69, 75, 63, 66, 78, 88, 93, 98, 86, 
    62, 69, 85, 99, 97, 56, 65, 74, 93, 89, 73, 82, 94, 87, 58, 
    80, 90, 80, 88, 80, 94, 73, 87, 86, 82, 80, 81, 75, 69, 69, 
    80, 76, 55, 56, 74, 54, 95, 93, 94, 97, 81, 82, 65, 45, 72, 
    77, 56, 76, 80, 79, 83, 77, 111, 96, 81, 80, 77, 72, 79, 90, 
    111, 134, 120, 87, 89, 86, 93, 94, 98, 88, 89, 75, 70, 67, 104, 
    63, 95, 149, 130, 106, 79, 98, 57, 59, 94, 90, 84, 57, 50, 87, 
    55, 12, 75, 142, 142, 110, 90, 92, 71, 77, 86, 71, 40, 25, 115, 
    60, 36, 20, 93, 148, 159, 134, 114, 66, 60, 52, 70, 71, 86, 81, 
    
    -- channel=76
    77, 64, 73, 83, 59, 37, 72, 65, 88, 86, 88, 84, 103, 53, 66, 
    106, 89, 97, 84, 51, 30, 54, 63, 95, 88, 92, 90, 128, 90, 110, 
    62, 57, 82, 68, 42, 62, 106, 86, 83, 71, 70, 117, 141, 126, 110, 
    82, 99, 96, 63, 55, 116, 115, 68, 62, 80, 119, 140, 138, 130, 105, 
    84, 109, 137, 66, 69, 126, 108, 65, 136, 130, 127, 131, 147, 129, 92, 
    71, 88, 139, 138, 123, 99, 59, 108, 129, 118, 109, 120, 145, 131, 93, 
    86, 102, 121, 139, 92, 82, 82, 100, 71, 67, 79, 104, 119, 140, 100, 
    88, 105, 119, 129, 104, 80, 74, 77, 99, 109, 93, 90, 103, 120, 89, 
    106, 128, 111, 118, 94, 84, 87, 91, 103, 97, 89, 95, 70, 79, 91, 
    108, 101, 86, 79, 110, 72, 89, 106, 99, 107, 87, 93, 83, 76, 96, 
    107, 80, 104, 112, 112, 110, 94, 121, 108, 90, 87, 87, 83, 105, 135, 
    131, 175, 173, 136, 119, 113, 107, 100, 107, 93, 95, 83, 84, 96, 146, 
    94, 113, 173, 182, 154, 107, 111, 64, 58, 95, 101, 90, 69, 78, 127, 
    84, 44, 98, 166, 191, 171, 144, 119, 107, 85, 92, 78, 56, 46, 145, 
    87, 64, 54, 126, 166, 201, 187, 172, 101, 58, 56, 79, 99, 136, 145, 
    
    -- channel=77
    51, 49, 56, 43, 46, 35, 54, 38, 54, 40, 62, 29, 89, 19, 50, 
    40, 66, 53, 42, 48, 28, 25, 42, 56, 56, 57, 26, 84, 58, 63, 
    45, 36, 45, 34, 42, 42, 70, 67, 23, 46, 38, 29, 79, 59, 68, 
    45, 40, 62, 45, 40, 72, 81, 29, 43, 50, 54, 67, 56, 55, 59, 
    56, 27, 72, 50, 55, 63, 62, 59, 66, 76, 84, 41, 64, 48, 61, 
    51, 18, 46, 80, 68, 41, 65, 62, 76, 55, 54, 71, 77, 39, 74, 
    67, 33, 28, 60, 56, 45, 64, 47, 46, 44, 48, 59, 59, 57, 70, 
    51, 34, 50, 49, 50, 53, 37, 60, 55, 61, 59, 30, 79, 54, 45, 
    49, 58, 36, 34, 21, 77, 37, 42, 53, 41, 53, 51, 38, 47, 66, 
    60, 33, 52, 42, 32, 3, 48, 49, 44, 52, 48, 53, 51, 53, 41, 
    48, 45, 68, 31, 61, 55, 20, 46, 47, 43, 38, 47, 61, 44, 67, 
    54, 92, 110, 63, 49, 35, 36, 40, 38, 51, 46, 54, 65, 58, 54, 
    33, 15, 91, 112, 80, 48, 35, 42, 7, 41, 37, 52, 65, 40, 67, 
    57, 24, 15, 78, 114, 89, 65, 68, 50, 34, 46, 57, 47, 68, 33, 
    66, 66, 25, 32, 77, 108, 106, 75, 56, 31, 27, 34, 79, 47, 62, 
    
    -- channel=78
    11, 0, 12, 0, 0, 30, 7, 8, 17, 13, 0, 36, 0, 39, 3, 
    1, 0, 0, 0, 0, 36, 11, 17, 0, 10, 0, 54, 0, 17, 3, 
    10, 17, 2, 0, 0, 21, 0, 0, 14, 0, 24, 43, 0, 3, 0, 
    0, 34, 0, 10, 0, 20, 0, 0, 36, 0, 35, 24, 0, 4, 0, 
    0, 46, 0, 0, 33, 15, 0, 12, 2, 6, 10, 16, 7, 3, 0, 
    0, 52, 0, 0, 26, 36, 13, 48, 17, 31, 18, 36, 0, 3, 0, 
    0, 35, 9, 2, 30, 65, 45, 62, 48, 55, 54, 62, 4, 7, 0, 
    0, 20, 11, 10, 45, 28, 74, 52, 58, 57, 55, 55, 35, 19, 0, 
    0, 9, 0, 1, 40, 42, 58, 55, 69, 66, 38, 62, 30, 22, 0, 
    4, 0, 0, 24, 20, 30, 61, 62, 49, 61, 49, 49, 27, 14, 3, 
    0, 24, 0, 14, 3, 23, 61, 56, 52, 42, 64, 51, 28, 4, 2, 
    0, 33, 0, 4, 0, 24, 68, 64, 53, 33, 74, 53, 39, 21, 0, 
    33, 42, 6, 0, 0, 9, 42, 47, 66, 52, 56, 49, 37, 13, 0, 
    5, 47, 59, 15, 0, 0, 3, 0, 40, 66, 59, 38, 12, 27, 12, 
    0, 14, 55, 56, 12, 0, 0, 10, 9, 56, 57, 29, 0, 13, 40, 
    
    -- channel=79
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 55, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 57, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 58, 0, 7, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 5, 67, 
    0, 0, 37, 0, 0, 0, 23, 0, 0, 0, 0, 0, 24, 16, 82, 
    3, 0, 16, 0, 0, 0, 14, 0, 0, 0, 18, 0, 25, 11, 71, 
    0, 0, 0, 25, 24, 8, 4, 4, 20, 18, 13, 0, 37, 0, 52, 
    0, 0, 0, 29, 32, 19, 8, 32, 26, 11, 14, 37, 43, 13, 42, 
    0, 0, 8, 9, 8, 39, 21, 43, 34, 44, 50, 16, 71, 13, 2, 
    0, 8, 0, 0, 10, 28, 20, 42, 52, 62, 37, 47, 56, 0, 0, 
    37, 0, 0, 0, 0, 0, 6, 57, 70, 65, 37, 45, 30, 0, 0, 
    0, 0, 3, 0, 21, 0, 15, 62, 58, 63, 35, 49, 28, 0, 0, 
    7, 13, 33, 0, 0, 0, 23, 68, 17, 50, 60, 50, 48, 0, 0, 
    17, 0, 0, 16, 11, 0, 0, 0, 0, 43, 47, 55, 52, 0, 0, 
    19, 0, 0, 0, 26, 5, 0, 0, 11, 22, 45, 26, 0, 0, 0, 
    
    -- channel=80
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 21, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=81
    0, 26, 31, 33, 27, 30, 18, 22, 7, 0, 0, 0, 0, 11, 0, 
    70, 57, 36, 39, 43, 31, 18, 20, 0, 0, 2, 3, 2, 1, 0, 
    69, 66, 50, 56, 55, 52, 33, 36, 26, 0, 0, 0, 4, 6, 2, 
    43, 66, 61, 64, 67, 53, 47, 34, 49, 36, 20, 10, 0, 4, 11, 
    58, 64, 59, 63, 64, 62, 42, 36, 33, 50, 49, 18, 7, 11, 11, 
    47, 51, 73, 72, 67, 84, 68, 94, 25, 37, 43, 0, 6, 3, 11, 
    57, 82, 87, 73, 60, 121, 71, 9, 31, 47, 20, 0, 0, 0, 6, 
    0, 84, 82, 79, 99, 81, 63, 98, 93, 79, 28, 0, 0, 7, 0, 
    9, 63, 79, 69, 126, 98, 86, 98, 97, 101, 37, 0, 1, 53, 0, 
    11, 90, 97, 33, 100, 91, 32, 29, 12, 0, 0, 0, 0, 72, 0, 
    27, 74, 100, 0, 1, 65, 26, 73, 16, 0, 0, 0, 0, 98, 34, 
    21, 45, 65, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 54, 55, 
    26, 34, 55, 80, 22, 9, 3, 0, 0, 0, 0, 0, 0, 0, 55, 
    35, 47, 34, 38, 35, 9, 35, 7, 0, 0, 0, 0, 0, 0, 0, 
    16, 31, 15, 20, 5, 24, 33, 25, 19, 2, 9, 20, 13, 4, 4, 
    
    -- channel=82
    0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 12, 4, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 21, 0, 0, 3, 0, 0, 
    57, 0, 0, 0, 15, 0, 0, 42, 12, 0, 13, 49, 9, 3, 3, 
    0, 22, 0, 0, 0, 0, 20, 0, 0, 0, 0, 8, 1, 0, 5, 
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 9, 15, 56, 19, 67, 58, 89, 112, 46, 4, 0, 0, 
    0, 1, 0, 11, 91, 0, 33, 0, 0, 42, 0, 0, 0, 0, 0, 
    0, 11, 19, 35, 3, 144, 99, 96, 96, 24, 48, 16, 0, 18, 0, 
    12, 0, 7, 0, 0, 0, 0, 0, 42, 33, 13, 41, 38, 42, 23, 
    0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 48, 
    6, 28, 0, 2, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 11, 0, 2, 0, 0, 0, 0, 0, 
    
    -- channel=83
    39, 33, 2, 11, 14, 12, 9, 12, 0, 0, 16, 30, 36, 10, 7, 
    0, 0, 11, 12, 13, 19, 20, 24, 34, 20, 7, 0, 7, 11, 15, 
    0, 0, 5, 0, 8, 4, 22, 10, 21, 57, 43, 23, 5, 2, 15, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 28, 18, 18, 26, 10, 
    0, 0, 0, 2, 0, 0, 16, 44, 5, 0, 0, 0, 1, 0, 6, 
    0, 18, 19, 0, 0, 19, 0, 0, 0, 13, 0, 0, 0, 2, 6, 
    0, 0, 0, 0, 17, 0, 0, 57, 64, 25, 0, 11, 15, 18, 3, 
    16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 43, 12, 
    16, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 5, 4, 
    27, 0, 0, 0, 0, 0, 0, 28, 7, 0, 42, 31, 6, 8, 12, 
    4, 0, 0, 0, 40, 0, 0, 0, 0, 0, 0, 4, 22, 0, 0, 
    0, 7, 0, 53, 32, 60, 42, 16, 22, 13, 10, 0, 6, 0, 0, 
    10, 12, 0, 0, 0, 0, 43, 43, 49, 61, 58, 56, 13, 26, 0, 
    0, 0, 0, 0, 0, 35, 7, 16, 36, 29, 46, 52, 53, 30, 0, 
    29, 23, 16, 19, 29, 17, 0, 0, 0, 16, 21, 19, 19, 19, 28, 
    
    -- channel=84
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 14, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 10, 8, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 9, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=85
    45, 33, 56, 68, 62, 59, 59, 47, 27, 26, 29, 16, 11, 26, 32, 
    54, 60, 59, 56, 61, 65, 71, 67, 34, 10, 25, 41, 50, 37, 31, 
    35, 46, 56, 64, 63, 64, 63, 68, 76, 33, 27, 41, 47, 50, 41, 
    45, 47, 57, 63, 71, 77, 78, 74, 74, 71, 46, 30, 32, 30, 39, 
    44, 42, 60, 56, 62, 64, 54, 45, 41, 68, 69, 45, 42, 45, 40, 
    38, 25, 31, 59, 56, 44, 25, 53, 67, 45, 39, 24, 26, 36, 38, 
    17, 67, 52, 45, 36, 39, 39, 11, 0, 17, 20, 8, 8, 23, 32, 
    31, 43, 50, 46, 42, 47, 59, 50, 38, 31, 18, 23, 23, 22, 18, 
    58, 50, 41, 42, 42, 30, 49, 71, 60, 56, 43, 7, 10, 26, 14, 
    47, 33, 37, 18, 53, 70, 62, 70, 38, 16, 6, 18, 26, 33, 1, 
    61, 55, 36, 14, 0, 0, 28, 39, 52, 24, 10, 28, 25, 44, 20, 
    69, 51, 34, 26, 36, 38, 42, 24, 0, 0, 0, 0, 19, 37, 43, 
    64, 58, 34, 50, 66, 68, 49, 38, 15, 0, 0, 0, 0, 11, 15, 
    51, 64, 65, 46, 36, 34, 51, 55, 40, 39, 34, 33, 29, 33, 37, 
    47, 47, 60, 60, 52, 53, 59, 68, 56, 49, 58, 58, 54, 46, 45, 
    
    -- channel=86
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=87
    76, 47, 58, 63, 68, 61, 61, 48, 52, 24, 33, 40, 36, 30, 48, 
    64, 65, 65, 67, 65, 72, 74, 67, 70, 30, 21, 31, 41, 51, 40, 
    60, 49, 66, 67, 69, 73, 79, 65, 66, 76, 40, 56, 45, 44, 48, 
    70, 44, 63, 65, 70, 78, 75, 72, 55, 71, 74, 65, 43, 42, 46, 
    41, 54, 67, 70, 73, 69, 69, 71, 68, 53, 66, 62, 29, 37, 43, 
    12, 72, 64, 65, 65, 42, 63, 28, 62, 42, 56, 47, 10, 34, 36, 
    0, 48, 65, 70, 61, 43, 69, 78, 42, 53, 62, 40, 15, 29, 33, 
    58, 18, 70, 52, 53, 72, 75, 57, 56, 61, 73, 35, 12, 31, 45, 
    69, 41, 68, 62, 37, 62, 77, 46, 46, 35, 40, 24, 0, 26, 75, 
    81, 31, 62, 85, 0, 43, 77, 47, 72, 35, 29, 23, 5, 13, 85, 
    80, 43, 57, 69, 19, 2, 34, 33, 50, 26, 5, 10, 24, 0, 74, 
    74, 67, 48, 80, 48, 48, 47, 46, 19, 0, 0, 0, 7, 15, 38, 
    77, 70, 66, 33, 73, 62, 64, 69, 47, 26, 15, 5, 0, 34, 16, 
    69, 54, 72, 60, 52, 55, 53, 83, 57, 51, 52, 42, 52, 40, 33, 
    70, 69, 81, 68, 76, 68, 70, 61, 65, 67, 62, 61, 69, 65, 50, 
    
    -- channel=88
    81, 0, 5, 0, 2, 0, 13, 0, 40, 5, 0, 6, 0, 0, 37, 
    2, 13, 14, 0, 0, 0, 16, 0, 43, 30, 0, 0, 0, 6, 5, 
    26, 0, 0, 0, 0, 3, 14, 0, 12, 58, 0, 25, 0, 0, 0, 
    62, 0, 0, 0, 0, 7, 8, 15, 0, 1, 22, 48, 1, 0, 0, 
    6, 0, 0, 0, 0, 4, 10, 0, 23, 0, 3, 75, 0, 0, 0, 
    0, 11, 0, 0, 12, 0, 25, 0, 46, 0, 9, 81, 0, 0, 0, 
    0, 0, 0, 6, 0, 0, 43, 43, 0, 0, 66, 59, 0, 0, 0, 
    18, 0, 9, 0, 0, 11, 17, 0, 0, 0, 72, 58, 0, 0, 44, 
    14, 0, 0, 49, 0, 0, 37, 0, 0, 3, 87, 40, 0, 0, 112, 
    27, 0, 0, 132, 0, 0, 86, 0, 54, 51, 24, 0, 0, 0, 118, 
    16, 0, 0, 152, 0, 0, 3, 0, 79, 38, 0, 0, 0, 0, 79, 
    29, 0, 0, 49, 41, 3, 0, 30, 43, 7, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 65, 18, 0, 41, 42, 22, 17, 0, 0, 17, 0, 
    0, 0, 26, 1, 30, 0, 0, 35, 7, 13, 14, 0, 14, 0, 0, 
    0, 0, 18, 0, 17, 0, 0, 4, 2, 12, 0, 0, 8, 16, 0, 
    
    -- channel=89
    0, 28, 34, 35, 28, 29, 17, 27, 0, 7, 20, 10, 14, 34, 2, 
    28, 22, 28, 40, 40, 30, 23, 33, 0, 0, 24, 25, 38, 25, 19, 
    24, 36, 34, 40, 40, 39, 26, 33, 25, 0, 37, 19, 37, 30, 28, 
    13, 51, 37, 44, 41, 42, 39, 25, 42, 42, 31, 0, 23, 30, 34, 
    38, 42, 40, 42, 41, 38, 37, 40, 25, 52, 33, 0, 20, 28, 33, 
    50, 51, 48, 42, 33, 46, 42, 44, 12, 51, 32, 0, 23, 16, 33, 
    69, 60, 56, 42, 40, 64, 35, 21, 52, 49, 11, 0, 10, 15, 26, 
    29, 92, 50, 52, 69, 54, 48, 74, 67, 62, 0, 0, 17, 39, 2, 
    36, 92, 56, 20, 68, 67, 33, 51, 48, 38, 0, 0, 23, 67, 0, 
    44, 92, 66, 0, 85, 65, 18, 72, 25, 0, 0, 0, 32, 89, 0, 
    46, 80, 58, 0, 16, 22, 22, 71, 0, 0, 0, 9, 21, 99, 2, 
    53, 64, 55, 5, 19, 19, 35, 15, 0, 0, 0, 0, 23, 46, 48, 
    53, 68, 45, 63, 0, 36, 52, 13, 0, 0, 0, 0, 19, 8, 46, 
    48, 73, 42, 41, 21, 42, 74, 36, 27, 22, 16, 30, 13, 25, 31, 
    55, 70, 50, 57, 42, 65, 50, 48, 43, 37, 47, 55, 42, 29, 31, 
    
    -- channel=90
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 25, 40, 0, 0, 8, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 1, 26, 0, 0, 43, 43, 67, 90, 9, 0, 0, 0, 
    0, 0, 0, 49, 28, 18, 19, 0, 0, 0, 0, 0, 0, 0, 7, 
    0, 0, 12, 35, 0, 10, 14, 0, 38, 10, 16, 0, 0, 0, 31, 
    0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 7, 1, 0, 0, 13, 
    0, 0, 0, 2, 0, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=91
    71, 53, 45, 39, 45, 35, 30, 31, 26, 10, 12, 15, 15, 15, 20, 
    61, 65, 49, 52, 49, 48, 40, 35, 28, 5, 5, 11, 23, 23, 18, 
    62, 59, 55, 53, 58, 52, 48, 35, 47, 54, 34, 26, 13, 17, 23, 
    71, 65, 57, 55, 61, 52, 47, 38, 38, 49, 47, 25, 12, 11, 20, 
    49, 56, 63, 61, 59, 53, 54, 57, 38, 26, 40, 36, 12, 17, 21, 
    17, 71, 61, 66, 56, 77, 87, 39, 47, 39, 30, 19, 5, 11, 16, 
    10, 59, 84, 74, 71, 81, 76, 83, 70, 73, 47, 12, 6, 12, 12, 
    33, 39, 79, 69, 90, 102, 80, 87, 95, 96, 62, 15, 14, 40, 22, 
    32, 56, 84, 53, 68, 73, 58, 41, 43, 28, 15, 0, 0, 45, 38, 
    36, 38, 94, 41, 15, 62, 56, 61, 44, 5, 7, 2, 4, 54, 74, 
    40, 38, 71, 46, 0, 0, 0, 0, 0, 0, 0, 0, 5, 34, 82, 
    40, 37, 58, 72, 45, 30, 29, 14, 0, 0, 0, 0, 0, 2, 52, 
    31, 46, 41, 51, 51, 35, 29, 30, 24, 13, 1, 3, 0, 4, 8, 
    26, 27, 42, 31, 33, 35, 33, 34, 31, 33, 34, 37, 39, 25, 30, 
    37, 37, 40, 40, 52, 44, 28, 28, 27, 23, 27, 37, 38, 33, 26, 
    
    -- channel=92
    65, 67, 40, 29, 37, 31, 19, 28, 26, 11, 8, 18, 16, 15, 12, 
    58, 63, 43, 51, 45, 41, 31, 27, 30, 16, 2, 1, 11, 20, 12, 
    73, 57, 53, 50, 54, 49, 41, 30, 31, 52, 34, 21, 4, 5, 17, 
    62, 69, 55, 51, 54, 40, 34, 30, 27, 37, 48, 29, 10, 8, 14, 
    52, 55, 59, 61, 55, 52, 51, 55, 42, 14, 29, 35, 4, 12, 16, 
    5, 84, 68, 67, 60, 78, 98, 34, 32, 37, 31, 16, 6, 8, 11, 
    27, 45, 84, 75, 72, 91, 72, 88, 85, 84, 51, 15, 12, 11, 10, 
    32, 38, 76, 69, 94, 101, 77, 86, 95, 100, 64, 13, 14, 42, 29, 
    15, 55, 84, 57, 71, 72, 50, 30, 31, 25, 5, 0, 4, 46, 40, 
    28, 44, 92, 46, 7, 58, 37, 43, 44, 3, 3, 0, 5, 55, 81, 
    27, 30, 76, 39, 17, 0, 0, 0, 0, 0, 0, 0, 9, 34, 80, 
    21, 27, 63, 62, 46, 15, 21, 17, 0, 0, 0, 0, 0, 5, 40, 
    19, 33, 43, 47, 39, 27, 12, 22, 24, 24, 14, 15, 8, 4, 11, 
    17, 9, 25, 26, 28, 25, 26, 17, 22, 23, 24, 33, 36, 24, 27, 
    22, 32, 22, 25, 42, 34, 20, 9, 19, 8, 15, 27, 28, 27, 17, 
    
    -- channel=93
    80, 83, 60, 69, 68, 67, 67, 57, 62, 36, 34, 43, 37, 37, 48, 
    74, 74, 67, 67, 69, 76, 79, 67, 75, 52, 25, 34, 37, 46, 40, 
    72, 60, 71, 68, 72, 73, 79, 69, 77, 87, 56, 57, 38, 38, 46, 
    60, 54, 66, 69, 74, 70, 70, 74, 60, 62, 63, 72, 36, 40, 40, 
    41, 59, 70, 69, 73, 75, 60, 70, 67, 45, 65, 78, 37, 39, 37, 
    2, 55, 67, 73, 65, 68, 73, 45, 48, 41, 54, 47, 26, 40, 34, 
    31, 37, 64, 66, 64, 68, 47, 69, 62, 62, 57, 45, 29, 40, 35, 
    47, 22, 61, 49, 58, 68, 76, 57, 51, 51, 80, 51, 19, 42, 58, 
    58, 33, 60, 69, 40, 26, 74, 36, 32, 28, 22, 27, 18, 28, 78, 
    49, 29, 53, 87, 0, 42, 48, 52, 70, 33, 38, 48, 19, 22, 87, 
    59, 30, 43, 53, 29, 0, 5, 7, 34, 40, 19, 16, 37, 7, 67, 
    38, 50, 35, 82, 60, 58, 55, 43, 37, 25, 24, 14, 8, 23, 23, 
    52, 38, 55, 25, 92, 49, 39, 68, 59, 46, 43, 32, 27, 24, 28, 
    49, 25, 54, 44, 43, 43, 34, 55, 53, 56, 54, 58, 62, 57, 34, 
    39, 51, 49, 54, 58, 48, 52, 41, 47, 42, 47, 47, 55, 55, 51, 
    
    -- channel=94
    51, 95, 99, 111, 107, 111, 99, 100, 60, 65, 73, 71, 69, 81, 55, 
    88, 91, 98, 109, 113, 110, 110, 120, 80, 54, 78, 76, 92, 82, 70, 
    71, 97, 104, 110, 112, 111, 112, 116, 100, 69, 87, 78, 94, 86, 84, 
    59, 96, 102, 110, 113, 120, 114, 111, 114, 110, 98, 68, 82, 89, 87, 
    75, 96, 105, 111, 108, 104, 91, 95, 86, 119, 100, 53, 83, 82, 86, 
    104, 91, 100, 99, 94, 82, 54, 65, 72, 98, 79, 37, 73, 76, 88, 
    118, 101, 86, 87, 80, 90, 61, 58, 66, 71, 43, 33, 62, 74, 81, 
    84, 121, 81, 75, 93, 68, 88, 91, 66, 66, 33, 32, 63, 79, 47, 
    88, 123, 75, 57, 112, 89, 71, 103, 93, 75, 39, 41, 77, 96, 23, 
    98, 113, 73, 26, 88, 98, 58, 115, 74, 50, 42, 56, 85, 104, 10, 
    97, 111, 79, 4, 87, 64, 76, 121, 41, 47, 49, 58, 82, 112, 23, 
    94, 112, 78, 50, 62, 76, 90, 71, 34, 30, 28, 51, 74, 94, 76, 
    110, 105, 95, 80, 53, 94, 101, 63, 48, 40, 31, 43, 67, 66, 95, 
    102, 111, 85, 104, 67, 96, 115, 91, 80, 73, 72, 84, 71, 84, 71, 
    99, 117, 98, 102, 91, 108, 106, 96, 101, 93, 106, 106, 94, 87, 88, 
    
    -- channel=95
    20, 0, 14, 9, 14, 5, 9, 0, 17, 0, 0, 0, 0, 0, 8, 
    21, 30, 2, 14, 17, 12, 8, 1, 15, 0, 0, 0, 0, 10, 0, 
    50, 16, 9, 19, 18, 22, 23, 2, 7, 0, 0, 0, 3, 6, 0, 
    24, 19, 21, 16, 26, 23, 33, 17, 13, 22, 6, 18, 3, 0, 4, 
    21, 17, 21, 13, 26, 25, 31, 20, 27, 13, 16, 47, 0, 2, 5, 
    0, 28, 22, 28, 29, 0, 59, 57, 36, 4, 34, 30, 0, 0, 0, 
    0, 9, 53, 45, 5, 33, 53, 34, 4, 9, 45, 9, 0, 0, 0, 
    14, 0, 59, 36, 16, 63, 31, 42, 54, 57, 63, 10, 0, 0, 15, 
    29, 0, 54, 37, 41, 30, 83, 39, 49, 58, 71, 0, 0, 0, 53, 
    40, 0, 62, 93, 8, 19, 81, 22, 46, 7, 0, 0, 0, 0, 91, 
    48, 3, 64, 87, 0, 8, 22, 15, 54, 0, 0, 0, 0, 0, 103, 
    43, 21, 36, 19, 5, 0, 0, 19, 0, 0, 0, 0, 0, 0, 41, 
    20, 36, 18, 42, 28, 20, 10, 18, 0, 0, 0, 0, 0, 0, 0, 
    45, 15, 56, 0, 56, 4, 16, 44, 5, 4, 0, 0, 0, 0, 23, 
    28, 19, 40, 18, 16, 31, 29, 32, 21, 15, 8, 15, 23, 25, 0, 
    
    -- channel=96
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 18, 14, 38, 
    0, 0, 0, 5, 24, 17, 17, 19, 32, 5, 0, 5, 53, 50, 35, 
    
    -- channel=97
    0, 0, 6, 7, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 39, 66, 124, 103, 35, 0, 3, 0, 0, 
    0, 0, 0, 0, 13, 69, 88, 43, 23, 36, 176, 0, 0, 0, 0, 
    0, 0, 0, 0, 1, 5, 0, 0, 0, 110, 158, 98, 0, 0, 0, 
    0, 0, 21, 38, 13, 18, 31, 151, 184, 179, 158, 0, 0, 0, 66, 
    0, 38, 0, 9, 0, 0, 71, 168, 155, 190, 153, 4, 65, 94, 108, 
    17, 151, 15, 0, 0, 0, 86, 145, 156, 16, 90, 187, 124, 111, 22, 
    6, 8, 37, 0, 0, 47, 111, 142, 24, 0, 0, 73, 92, 17, 0, 
    0, 11, 50, 0, 0, 20, 134, 145, 4, 0, 0, 0, 105, 0, 0, 
    0, 15, 61, 25, 97, 141, 157, 156, 27, 29, 9, 0, 10, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 2, 0, 0, 0, 0, 
    
    -- channel=98
    0, 0, 9, 24, 31, 31, 32, 26, 31, 63, 25, 15, 26, 46, 0, 
    32, 13, 25, 37, 37, 28, 25, 21, 15, 0, 0, 9, 5, 0, 0, 
    43, 65, 46, 27, 19, 4, 2, 0, 0, 0, 0, 8, 0, 0, 0, 
    20, 3, 0, 0, 0, 0, 0, 0, 0, 0, 33, 36, 0, 5, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 11, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 45, 0, 0, 67, 0, 7, 
    0, 0, 0, 1, 0, 59, 128, 167, 112, 32, 0, 0, 0, 60, 27, 
    0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 32, 0, 0, 0, 
    0, 0, 28, 70, 25, 55, 21, 0, 0, 15, 2, 86, 0, 0, 0, 
    0, 0, 0, 16, 31, 19, 0, 0, 7, 65, 77, 0, 0, 0, 25, 
    13, 96, 24, 0, 29, 0, 0, 0, 44, 157, 129, 144, 23, 60, 120, 
    24, 16, 0, 0, 0, 0, 0, 0, 20, 0, 4, 51, 29, 39, 19, 
    24, 0, 0, 0, 0, 0, 0, 10, 2, 0, 0, 8, 66, 66, 18, 
    0, 1, 41, 66, 108, 199, 218, 229, 147, 9, 48, 24, 70, 52, 3, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 40, 25, 27, 0, 0, 0, 
    
    -- channel=99
    63, 55, 48, 47, 46, 48, 46, 49, 45, 2, 33, 42, 1, 5, 42, 
    69, 65, 54, 57, 56, 54, 52, 54, 51, 50, 83, 40, 15, 37, 60, 
    17, 28, 48, 56, 57, 62, 61, 61, 59, 64, 14, 0, 53, 45, 41, 
    55, 61, 62, 63, 65, 63, 82, 79, 70, 52, 0, 0, 15, 32, 48, 
    61, 63, 60, 58, 62, 52, 38, 71, 147, 146, 72, 27, 56, 50, 52, 
    63, 65, 60, 58, 71, 114, 43, 0, 0, 0, 32, 16, 0, 47, 47, 
    65, 61, 54, 67, 31, 0, 0, 0, 0, 43, 0, 39, 23, 0, 26, 
    60, 60, 82, 59, 14, 0, 13, 180, 231, 68, 0, 0, 0, 38, 113, 
    56, 86, 28, 0, 0, 0, 14, 0, 0, 0, 0, 0, 107, 110, 0, 
    88, 126, 7, 0, 0, 0, 0, 0, 0, 0, 0, 28, 28, 0, 0, 
    27, 0, 0, 0, 2, 85, 21, 0, 0, 0, 0, 0, 0, 0, 0, 
    25, 0, 0, 0, 49, 0, 0, 0, 0, 17, 13, 0, 0, 0, 9, 
    35, 0, 0, 40, 97, 86, 0, 0, 0, 21, 40, 0, 0, 0, 7, 
    39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    31, 38, 64, 66, 43, 48, 38, 33, 30, 0, 0, 0, 25, 26, 27, 
    
    -- channel=100
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 20, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 15, 26, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 49, 59, 38, 27, 66, 24, 26, 5, 0, 
    0, 0, 0, 0, 4, 1, 14, 9, 15, 33, 64, 69, 14, 9, 0, 
    0, 0, 0, 24, 37, 27, 25, 35, 45, 55, 63, 38, 0, 13, 27, 
    0, 0, 27, 44, 34, 32, 23, 69, 67, 79, 37, 0, 26, 52, 57, 
    0, 38, 53, 47, 24, 20, 54, 68, 91, 56, 72, 68, 67, 75, 43, 
    0, 35, 62, 41, 19, 52, 55, 65, 65, 30, 38, 48, 61, 62, 16, 
    0, 34, 60, 35, 33, 51, 68, 71, 61, 29, 38, 36, 63, 42, 9, 
    0, 27, 65, 52, 72, 83, 82, 83, 55, 39, 46, 37, 47, 30, 16, 
    0, 7, 37, 36, 32, 32, 35, 33, 29, 42, 33, 23, 21, 19, 18, 
    
    -- channel=101
    163, 171, 181, 186, 177, 162, 156, 145, 127, 99, 92, 63, 33, 40, 64, 
    169, 159, 159, 156, 146, 133, 127, 118, 107, 99, 72, 46, 12, 26, 75, 
    138, 125, 121, 122, 112, 108, 104, 102, 96, 89, 58, 35, 24, 50, 83, 
    94, 101, 104, 103, 105, 104, 103, 93, 92, 77, 22, 2, 53, 78, 84, 
    96, 106, 109, 108, 107, 105, 99, 76, 28, 0, 0, 2, 60, 84, 83, 
    102, 107, 105, 104, 85, 45, 50, 103, 111, 87, 10, 0, 16, 58, 74, 
    107, 107, 102, 86, 71, 45, 0, 0, 0, 0, 0, 0, 0, 0, 51, 
    109, 101, 76, 45, 17, 8, 0, 0, 0, 0, 0, 4, 21, 0, 0, 
    106, 72, 7, 0, 0, 0, 0, 8, 12, 0, 0, 0, 0, 0, 0, 
    77, 34, 0, 0, 0, 0, 0, 0, 0, 13, 58, 16, 0, 0, 0, 
    85, 48, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    55, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    43, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 9, 0, 5, 0, 1, 8, 7, 5, 0, 0, 0, 0, 0, 0, 
    32, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 0, 
    
    -- channel=102
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 43, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 35, 42, 31, 49, 64, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 0, 0, 48, 90, 40, 25, 0, 0, 
    0, 0, 0, 0, 0, 18, 22, 23, 69, 105, 88, 63, 0, 14, 6, 
    0, 0, 0, 34, 23, 11, 67, 89, 79, 78, 46, 9, 14, 67, 57, 
    0, 22, 48, 39, 18, 32, 70, 80, 91, 82, 75, 69, 88, 70, 42, 
    0, 49, 44, 25, 12, 35, 90, 86, 52, 8, 11, 78, 75, 52, 0, 
    0, 41, 54, 27, 31, 61, 85, 96, 38, 23, 29, 40, 63, 30, 1, 
    0, 41, 58, 48, 71, 82, 87, 87, 49, 46, 35, 25, 39, 19, 0, 
    0, 30, 40, 38, 31, 27, 27, 27, 23, 20, 31, 20, 3, 10, 2, 
    0, 11, 39, 46, 42, 39, 32, 24, 14, 26, 26, 4, 10, 8, 12, 
    
    -- channel=103
    135, 133, 127, 127, 124, 116, 108, 107, 88, 86, 74, 58, 27, 16, 58, 
    125, 123, 118, 118, 108, 101, 94, 92, 85, 81, 69, 43, 23, 27, 68, 
    90, 96, 97, 97, 89, 90, 91, 85, 82, 79, 35, 33, 28, 46, 72, 
    79, 85, 88, 91, 88, 95, 94, 96, 85, 72, 30, 0, 60, 73, 72, 
    81, 90, 92, 93, 90, 85, 76, 88, 97, 93, 44, 18, 57, 67, 65, 
    89, 94, 95, 90, 84, 73, 34, 21, 6, 8, 53, 79, 0, 60, 62, 
    93, 95, 93, 81, 44, 19, 26, 19, 10, 0, 0, 130, 6, 0, 39, 
    93, 98, 71, 55, 40, 15, 21, 48, 33, 13, 49, 54, 60, 0, 24, 
    95, 83, 38, 0, 5, 0, 0, 0, 39, 56, 78, 109, 32, 30, 16, 
    90, 48, 77, 0, 17, 0, 0, 17, 43, 20, 5, 95, 33, 37, 38, 
    45, 0, 60, 5, 7, 0, 0, 28, 45, 50, 0, 0, 42, 29, 32, 
    37, 26, 0, 20, 0, 0, 0, 37, 76, 1, 2, 0, 19, 40, 13, 
    24, 2, 0, 38, 0, 24, 2, 45, 85, 0, 31, 0, 0, 41, 0, 
    29, 0, 0, 0, 0, 0, 0, 0, 20, 0, 13, 6, 0, 0, 0, 
    29, 25, 5, 3, 0, 0, 0, 0, 0, 0, 0, 9, 0, 0, 0, 
    
    -- channel=104
    0, 8, 0, 7, 17, 14, 0, 26, 1, 0, 11, 13, 17, 0, 9, 
    4, 15, 17, 14, 9, 11, 0, 13, 4, 7, 0, 25, 47, 0, 5, 
    2, 20, 12, 11, 1, 3, 0, 0, 0, 0, 0, 60, 17, 0, 10, 
    0, 0, 0, 5, 0, 0, 0, 0, 0, 1, 47, 0, 0, 2, 11, 
    0, 0, 1, 3, 0, 0, 0, 0, 0, 11, 59, 0, 0, 3, 3, 
    0, 2, 2, 1, 0, 0, 0, 0, 0, 15, 0, 181, 0, 12, 4, 
    0, 3, 7, 0, 0, 0, 4, 53, 0, 0, 0, 233, 42, 0, 1, 
    2, 8, 0, 0, 14, 0, 23, 0, 0, 0, 0, 125, 115, 0, 0, 
    4, 0, 6, 0, 34, 0, 0, 0, 0, 0, 21, 229, 0, 0, 0, 
    0, 0, 167, 0, 86, 0, 0, 0, 0, 3, 0, 95, 0, 0, 7, 
    0, 0, 115, 11, 60, 0, 0, 0, 18, 151, 0, 0, 32, 19, 125, 
    0, 25, 0, 83, 0, 0, 0, 0, 183, 0, 21, 0, 0, 115, 35, 
    0, 0, 0, 107, 0, 0, 0, 0, 202, 0, 43, 2, 0, 161, 0, 
    0, 0, 0, 42, 0, 0, 0, 0, 112, 0, 33, 55, 0, 49, 0, 
    0, 16, 8, 12, 2, 0, 0, 5, 7, 0, 11, 68, 0, 0, 0, 
    
    -- channel=105
    59, 43, 51, 39, 34, 32, 38, 22, 35, 35, 18, 16, 0, 6, 17, 
    46, 36, 45, 43, 43, 37, 42, 28, 29, 23, 30, 0, 0, 27, 25, 
    39, 41, 38, 39, 39, 39, 42, 32, 32, 36, 24, 0, 0, 39, 24, 
    35, 40, 42, 38, 43, 47, 49, 41, 37, 35, 0, 4, 31, 28, 23, 
    46, 46, 46, 43, 52, 45, 44, 57, 59, 26, 0, 10, 23, 22, 23, 
    48, 47, 43, 41, 55, 62, 59, 60, 77, 70, 61, 0, 11, 19, 21, 
    47, 48, 41, 47, 43, 64, 34, 0, 0, 69, 161, 0, 0, 21, 13, 
    49, 46, 46, 37, 12, 19, 12, 21, 61, 118, 127, 22, 0, 5, 33, 
    50, 57, 15, 23, 0, 7, 50, 143, 128, 124, 98, 0, 59, 42, 103, 
    67, 89, 0, 22, 0, 0, 87, 133, 104, 82, 106, 41, 90, 84, 48, 
    74, 110, 0, 0, 0, 12, 102, 111, 52, 0, 31, 128, 72, 41, 0, 
    52, 0, 41, 0, 0, 55, 111, 105, 0, 0, 0, 74, 67, 0, 0, 
    30, 25, 60, 0, 45, 67, 128, 96, 0, 37, 0, 0, 72, 0, 0, 
    21, 25, 33, 0, 44, 53, 51, 48, 0, 41, 9, 0, 8, 0, 0, 
    23, 2, 0, 0, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 
    
    -- channel=106
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 28, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 8, 97, 108, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 41, 39, 32, 17, 0, 0, 0, 0, 17, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 88, 31, 0, 0, 
    0, 0, 0, 0, 49, 6, 0, 0, 10, 0, 7, 0, 0, 0, 0, 
    0, 0, 0, 0, 20, 0, 0, 0, 0, 77, 86, 0, 0, 0, 20, 
    0, 97, 45, 7, 2, 0, 0, 0, 68, 58, 12, 14, 36, 45, 112, 
    0, 0, 0, 11, 0, 0, 0, 0, 77, 0, 0, 0, 0, 60, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 26, 0, 0, 0, 39, 58, 0, 
    0, 0, 69, 73, 97, 131, 141, 143, 117, 2, 7, 0, 37, 8, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 52, 20, 0, 0, 0, 
    
    -- channel=107
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 8, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 3, 10, 40, 42, 35, 11, 0, 0, 0, 
    0, 0, 0, 0, 0, 22, 58, 71, 64, 82, 140, 49, 0, 7, 0, 
    0, 0, 0, 0, 0, 16, 16, 0, 0, 31, 126, 127, 0, 0, 0, 
    0, 0, 0, 7, 26, 16, 41, 77, 109, 126, 159, 96, 30, 0, 43, 
    0, 0, 0, 11, 20, 0, 38, 127, 151, 157, 140, 58, 32, 56, 103, 
    0, 54, 73, 8, 2, 0, 43, 127, 135, 89, 107, 144, 107, 106, 70, 
    0, 45, 68, 9, 0, 19, 55, 129, 87, 29, 0, 39, 108, 71, 28, 
    0, 12, 58, 21, 2, 27, 86, 140, 99, 6, 5, 1, 76, 49, 0, 
    0, 16, 56, 39, 53, 102, 106, 128, 88, 29, 41, 0, 20, 19, 0, 
    0, 0, 17, 3, 0, 2, 5, 7, 16, 12, 22, 0, 0, 0, 0, 
    0, 4, 19, 12, 4, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=108
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 4, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 46, 56, 50, 31, 0, 0, 0, 
    0, 0, 0, 0, 0, 13, 54, 50, 41, 53, 138, 78, 0, 0, 0, 
    0, 0, 0, 0, 0, 17, 32, 8, 0, 51, 155, 124, 28, 0, 0, 
    0, 0, 0, 1, 28, 20, 58, 107, 150, 173, 181, 99, 6, 19, 54, 
    0, 0, 13, 12, 35, 20, 47, 145, 166, 165, 169, 60, 39, 67, 121, 
    0, 46, 92, 21, 10, 0, 55, 149, 147, 98, 83, 131, 131, 125, 81, 
    0, 53, 61, 25, 0, 37, 91, 150, 108, 28, 18, 42, 114, 75, 31, 
    0, 22, 72, 36, 15, 52, 99, 158, 113, 22, 16, 23, 77, 67, 0, 
    0, 26, 78, 59, 82, 135, 151, 151, 99, 41, 54, 8, 32, 17, 0, 
    0, 1, 25, 0, 7, 3, 4, 3, 0, 24, 38, 4, 0, 0, 0, 
    0, 20, 44, 37, 26, 28, 25, 16, 7, 2, 0, 0, 0, 0, 3, 
    
    -- channel=109
    101, 103, 99, 104, 100, 91, 84, 87, 70, 48, 60, 46, 49, 15, 44, 
    91, 99, 81, 76, 70, 67, 62, 67, 61, 62, 48, 67, 37, 16, 46, 
    65, 50, 53, 57, 55, 55, 54, 62, 60, 53, 68, 35, 41, 40, 57, 
    44, 48, 51, 55, 53, 53, 56, 65, 68, 64, 51, 2, 31, 45, 49, 
    43, 48, 49, 52, 46, 62, 55, 44, 48, 85, 68, 30, 41, 51, 48, 
    45, 49, 52, 52, 38, 45, 78, 77, 44, 5, 51, 81, 2, 41, 43, 
    50, 49, 52, 37, 61, 9, 0, 0, 0, 0, 0, 91, 40, 0, 25, 
    47, 48, 44, 59, 37, 25, 24, 27, 61, 74, 17, 45, 43, 10, 32, 
    46, 36, 51, 4, 19, 0, 0, 28, 18, 3, 21, 26, 0, 58, 20, 
    27, 70, 82, 2, 22, 9, 0, 0, 7, 17, 0, 61, 52, 22, 30, 
    36, 0, 30, 21, 18, 9, 0, 2, 32, 0, 0, 0, 7, 15, 0, 
    27, 23, 8, 28, 17, 5, 0, 16, 45, 13, 25, 0, 0, 25, 19, 
    27, 12, 0, 28, 14, 26, 6, 6, 61, 0, 42, 23, 0, 20, 10, 
    29, 17, 0, 3, 0, 0, 0, 0, 0, 0, 0, 27, 0, 13, 16, 
    28, 25, 13, 41, 22, 22, 23, 19, 21, 0, 13, 21, 23, 23, 22, 
    
    -- channel=110
    236, 234, 246, 245, 231, 217, 213, 192, 184, 158, 140, 109, 64, 74, 113, 
    229, 208, 211, 211, 197, 183, 183, 168, 158, 149, 138, 77, 35, 104, 130, 
    180, 173, 173, 171, 166, 163, 164, 158, 153, 145, 97, 22, 59, 119, 129, 
    152, 159, 162, 158, 163, 165, 166, 159, 147, 125, 38, 58, 120, 142, 133, 
    156, 164, 165, 162, 165, 152, 146, 138, 124, 70, 0, 46, 106, 126, 134, 
    163, 163, 161, 158, 152, 116, 60, 44, 56, 15, 24, 0, 46, 94, 122, 
    165, 162, 155, 144, 109, 81, 37, 11, 33, 48, 47, 0, 1, 49, 82, 
    163, 157, 121, 79, 43, 36, 18, 23, 14, 39, 9, 0, 14, 31, 59, 
    161, 137, 63, 18, 2, 30, 15, 58, 22, 11, 16, 0, 57, 32, 41, 
    142, 107, 0, 19, 0, 27, 56, 27, 0, 0, 12, 0, 13, 7, 12, 
    131, 49, 0, 9, 0, 31, 44, 6, 0, 0, 44, 50, 0, 0, 0, 
    111, 18, 16, 0, 15, 36, 43, 0, 0, 22, 0, 59, 19, 0, 18, 
    84, 29, 23, 0, 19, 3, 35, 0, 0, 25, 0, 20, 55, 0, 45, 
    81, 42, 21, 0, 38, 30, 29, 24, 0, 57, 0, 0, 39, 1, 32, 
    69, 35, 0, 0, 0, 1, 3, 9, 11, 38, 17, 1, 19, 20, 23, 
    
    -- channel=111
    0, 5, 13, 15, 24, 16, 12, 13, 0, 31, 0, 0, 6, 0, 0, 
    17, 23, 25, 24, 20, 15, 10, 7, 0, 0, 0, 0, 0, 0, 0, 
    24, 29, 18, 13, 3, 3, 4, 0, 0, 0, 7, 13, 0, 0, 4, 
    0, 0, 0, 2, 0, 2, 0, 1, 0, 0, 31, 0, 0, 0, 0, 
    0, 1, 3, 5, 1, 7, 7, 9, 0, 21, 13, 0, 0, 0, 0, 
    0, 4, 6, 3, 0, 0, 27, 51, 71, 101, 44, 49, 0, 4, 0, 
    3, 7, 12, 0, 0, 25, 64, 34, 5, 0, 67, 152, 0, 8, 0, 
    6, 11, 0, 2, 15, 0, 10, 0, 0, 0, 102, 196, 22, 0, 0, 
    11, 0, 6, 13, 40, 0, 0, 38, 109, 124, 152, 114, 0, 0, 41, 
    0, 0, 81, 0, 7, 0, 0, 89, 100, 142, 104, 84, 38, 70, 86, 
    0, 80, 97, 0, 0, 0, 0, 88, 149, 61, 0, 29, 115, 94, 83, 
    0, 0, 42, 22, 0, 0, 0, 94, 176, 0, 0, 0, 52, 103, 0, 
    0, 0, 28, 11, 0, 4, 19, 94, 150, 0, 11, 0, 7, 58, 0, 
    0, 0, 23, 7, 0, 51, 65, 75, 94, 0, 39, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 
    
    -- channel=112
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=113
    41, 36, 43, 47, 55, 55, 46, 29, 17, 17, 8, 0, 0, 0, 0, 
    40, 32, 43, 29, 53, 76, 58, 44, 22, 7, 0, 0, 0, 0, 0, 
    39, 34, 32, 30, 46, 52, 67, 63, 42, 26, 27, 30, 26, 23, 14, 
    30, 27, 0, 18, 43, 47, 48, 62, 74, 86, 66, 47, 27, 13, 1, 
    26, 40, 43, 0, 43, 60, 60, 55, 69, 75, 87, 65, 35, 15, 12, 
    97, 114, 61, 4, 20, 73, 89, 68, 65, 62, 73, 80, 62, 38, 32, 
    111, 105, 78, 0, 54, 84, 78, 70, 76, 62, 65, 78, 65, 57, 36, 
    92, 92, 101, 57, 0, 26, 45, 71, 93, 74, 63, 72, 68, 43, 15, 
    99, 102, 85, 82, 87, 60, 60, 64, 100, 83, 69, 66, 71, 50, 21, 
    122, 160, 200, 134, 140, 95, 87, 69, 97, 90, 82, 70, 69, 17, 0, 
    202, 201, 115, 137, 126, 107, 92, 76, 89, 91, 80, 67, 50, 5, 0, 
    208, 163, 82, 55, 36, 60, 57, 23, 75, 78, 72, 60, 34, 33, 0, 
    93, 79, 63, 56, 26, 10, 60, 40, 53, 79, 86, 77, 31, 26, 21, 
    45, 49, 58, 48, 28, 18, 20, 45, 44, 81, 98, 71, 51, 11, 24, 
    40, 29, 12, 0, 1, 26, 24, 2, 0, 7, 28, 38, 10, 0, 0, 
    
    -- channel=114
    0, 0, 0, 3, 8, 0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 
    0, 0, 0, 21, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 18, 9, 17, 1, 9, 4, 0, 0, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 6, 0, 0, 0, 0, 22, 0, 1, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 5, 0, 0, 0, 
    13, 14, 0, 0, 24, 21, 0, 0, 0, 0, 0, 0, 1, 20, 28, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 7, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    0, 0, 0, 0, 28, 0, 6, 0, 0, 0, 0, 0, 0, 14, 8, 
    0, 3, 87, 122, 65, 72, 30, 36, 0, 0, 2, 0, 0, 0, 0, 
    106, 144, 40, 0, 7, 29, 0, 0, 44, 16, 0, 0, 0, 0, 0, 
    59, 32, 30, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 6, 40, 44, 0, 0, 0, 0, 26, 47, 9, 8, 10, 11, 
    13, 44, 34, 6, 1, 0, 0, 7, 0, 0, 8, 23, 15, 7, 10, 
    
    -- channel=115
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 34, 35, 30, 20, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    0, 0, 40, 0, 0, 1, 2, 0, 0, 0, 0, 0, 0, 0, 2, 
    46, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 9, 11, 
    0, 0, 0, 0, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 36, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 54, 48, 0, 0, 0, 0, 0, 0, 0, 0, 5, 
    0, 4, 50, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 6, 8, 0, 0, 0, 7, 2, 0, 0, 0, 6, 7, 
    
    -- channel=116
    29, 28, 24, 28, 19, 3, 19, 24, 23, 24, 25, 26, 24, 20, 20, 
    29, 28, 25, 22, 7, 0, 0, 0, 14, 17, 12, 11, 8, 8, 10, 
    30, 28, 27, 8, 0, 0, 0, 0, 0, 5, 2, 3, 3, 8, 8, 
    24, 22, 18, 13, 0, 0, 0, 0, 0, 0, 1, 0, 5, 11, 0, 
    15, 14, 19, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    19, 24, 23, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    27, 27, 25, 6, 15, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 21, 22, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    14, 10, 9, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    15, 17, 33, 14, 11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 42, 30, 37, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    45, 49, 24, 6, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    36, 27, 27, 16, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    18, 14, 9, 0, 0, 0, 0, 0, 0, 0, 2, 0, 0, 0, 0, 
    7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=117
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 3, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 4, 6, 3, 
    0, 0, 0, 0, 0, 0, 0, 7, 5, 0, 0, 0, 0, 0, 2, 
    0, 0, 0, 0, 0, 4, 0, 0, 7, 3, 0, 4, 7, 9, 16, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 4, 0, 10, 27, 22, 
    0, 0, 0, 0, 0, 24, 7, 0, 0, 0, 2, 3, 9, 19, 13, 
    0, 0, 0, 19, 0, 0, 0, 3, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 10, 2, 0, 0, 0, 0, 0, 13, 29, 
    0, 11, 27, 24, 6, 8, 3, 4, 0, 0, 0, 0, 0, 3, 20, 
    0, 3, 0, 0, 0, 1, 1, 17, 5, 0, 1, 0, 0, 14, 20, 
    23, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 7, 29, 22, 
    0, 0, 0, 0, 16, 19, 12, 0, 0, 0, 0, 0, 13, 22, 29, 
    0, 0, 13, 18, 12, 7, 3, 6, 13, 3, 0, 0, 7, 34, 32, 
    17, 19, 14, 17, 29, 26, 20, 28, 27, 17, 17, 20, 23, 31, 35, 
    
    -- channel=118
    26, 22, 21, 22, 0, 0, 6, 11, 15, 12, 12, 11, 9, 8, 8, 
    25, 21, 15, 7, 0, 0, 0, 0, 3, 3, 2, 5, 10, 11, 9, 
    20, 18, 9, 0, 0, 0, 0, 0, 0, 5, 5, 0, 4, 3, 0, 
    16, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    31, 41, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 32, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 26, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 27, 20, 25, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    24, 27, 40, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    66, 63, 57, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    60, 53, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 13, 29, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    20, 11, 7, 6, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=119
    2, 3, 1, 6, 4, 4, 6, 2, 1, 0, 0, 0, 0, 0, 1, 
    2, 5, 0, 7, 0, 0, 0, 0, 0, 4, 8, 11, 8, 11, 13, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 13, 16, 15, 15, 15, 
    0, 2, 29, 0, 0, 0, 0, 0, 0, 0, 5, 14, 17, 21, 20, 
    18, 21, 35, 19, 0, 0, 0, 0, 0, 0, 0, 0, 17, 35, 31, 
    27, 29, 44, 17, 0, 0, 0, 0, 0, 0, 0, 0, 5, 37, 36, 
    24, 29, 34, 70, 0, 0, 0, 0, 0, 0, 0, 0, 2, 13, 24, 
    25, 32, 34, 29, 59, 2, 9, 0, 0, 0, 0, 0, 0, 0, 22, 
    29, 44, 64, 64, 45, 52, 18, 8, 0, 0, 0, 0, 0, 0, 24, 
    54, 57, 46, 74, 7, 33, 1, 17, 0, 0, 0, 0, 0, 13, 26, 
    68, 69, 87, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 30, 
    35, 39, 40, 11, 15, 0, 0, 15, 0, 0, 0, 0, 3, 9, 50, 
    15, 11, 19, 18, 14, 6, 0, 5, 0, 0, 0, 0, 16, 18, 22, 
    12, 12, 10, 15, 22, 21, 9, 0, 0, 0, 0, 0, 0, 19, 19, 
    10, 16, 21, 25, 17, 18, 22, 25, 21, 11, 0, 0, 17, 22, 26, 
    
    -- channel=120
    0, 2, 0, 0, 0, 0, 7, 2, 5, 0, 7, 11, 9, 0, 10, 
    0, 2, 0, 17, 0, 0, 7, 6, 12, 0, 3, 0, 0, 0, 1, 
    0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 3, 11, 
    0, 0, 35, 0, 0, 0, 0, 0, 0, 0, 0, 14, 2, 7, 5, 
    0, 0, 7, 74, 0, 0, 0, 18, 0, 0, 0, 0, 0, 2, 0, 
    0, 0, 52, 73, 0, 0, 0, 20, 0, 0, 0, 0, 0, 0, 5, 
    0, 0, 7, 116, 0, 0, 15, 0, 0, 7, 3, 0, 0, 0, 18, 
    0, 0, 0, 26, 83, 0, 3, 0, 0, 14, 12, 0, 0, 0, 5, 
    0, 0, 0, 40, 0, 28, 0, 18, 0, 5, 8, 7, 0, 2, 20, 
    0, 0, 0, 75, 0, 29, 0, 45, 0, 0, 0, 20, 0, 38, 11, 
    0, 0, 157, 0, 0, 11, 0, 7, 0, 0, 3, 17, 6, 3, 19, 
    21, 37, 62, 15, 44, 0, 0, 39, 0, 0, 0, 7, 26, 0, 46, 
    11, 0, 1, 0, 26, 14, 0, 24, 0, 0, 0, 6, 36, 0, 0, 
    0, 0, 0, 14, 10, 0, 3, 0, 1, 0, 0, 12, 11, 12, 0, 
    2, 12, 8, 11, 0, 0, 5, 22, 6, 0, 0, 0, 18, 0, 0, 
    
    -- channel=121
    6, 1, 16, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 0, 
    1, 1, 0, 0, 0, 0, 0, 0, 0, 4, 5, 7, 7, 8, 1, 
    0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 5, 0, 
    26, 37, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 12, 13, 9, 
    61, 59, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 3, 23, 16, 
    54, 51, 41, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 16, 6, 
    46, 53, 45, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    59, 80, 74, 21, 28, 0, 3, 0, 0, 0, 0, 0, 0, 0, 0, 
    103, 121, 110, 23, 44, 4, 14, 0, 0, 0, 0, 0, 0, 0, 0, 
    130, 107, 7, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    79, 56, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 
    14, 24, 23, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 
    10, 13, 7, 2, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 
    4, 1, 0, 0, 7, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=122
    1, 4, 0, 9, 17, 15, 6, 9, 4, 7, 10, 11, 6, 0, 0, 
    2, 2, 5, 0, 31, 46, 49, 26, 8, 0, 0, 0, 0, 0, 0, 
    7, 8, 25, 31, 33, 38, 49, 32, 3, 0, 0, 0, 0, 7, 9, 
    1, 0, 0, 0, 37, 20, 12, 29, 40, 32, 24, 19, 0, 0, 0, 
    0, 0, 0, 18, 32, 30, 19, 30, 38, 44, 45, 34, 0, 0, 0, 
    0, 0, 25, 0, 5, 0, 34, 46, 29, 32, 47, 38, 2, 0, 0, 
    3, 0, 0, 0, 0, 61, 66, 44, 26, 24, 42, 37, 32, 13, 15, 
    0, 0, 0, 0, 0, 0, 2, 22, 34, 40, 43, 44, 40, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 22, 38, 40, 34, 45, 34, 24, 42, 
    0, 0, 24, 74, 37, 59, 10, 37, 35, 36, 36, 51, 44, 23, 0, 
    0, 2, 54, 36, 60, 85, 58, 47, 45, 50, 53, 38, 24, 0, 0, 
    116, 70, 3, 32, 25, 36, 8, 16, 20, 21, 13, 27, 19, 0, 0, 
    19, 31, 0, 0, 12, 18, 45, 25, 24, 16, 24, 38, 27, 0, 0, 
    0, 0, 33, 49, 16, 0, 0, 22, 38, 51, 66, 47, 39, 11, 2, 
    38, 40, 10, 0, 0, 0, 7, 11, 1, 4, 18, 34, 27, 0, 0, 
    
    -- channel=123
    51, 48, 46, 45, 50, 60, 49, 41, 37, 31, 25, 18, 12, 10, 11, 
    50, 47, 41, 39, 47, 48, 59, 51, 34, 34, 34, 34, 36, 37, 34, 
    44, 44, 27, 25, 41, 44, 45, 49, 56, 62, 57, 52, 41, 35, 26, 
    41, 47, 48, 14, 39, 48, 49, 52, 50, 49, 61, 56, 40, 36, 30, 
    80, 96, 87, 39, 36, 60, 77, 64, 56, 54, 54, 61, 54, 46, 43, 
    101, 101, 103, 36, 54, 61, 73, 67, 64, 60, 55, 58, 50, 49, 42, 
    89, 89, 98, 70, 19, 48, 68, 69, 71, 66, 59, 56, 54, 36, 30, 
    91, 97, 93, 93, 93, 49, 67, 62, 78, 80, 65, 54, 54, 43, 36, 
    106, 124, 149, 118, 122, 87, 72, 69, 75, 81, 73, 64, 58, 44, 20, 
    161, 170, 146, 141, 106, 100, 71, 74, 75, 81, 80, 72, 56, 34, 2, 
    173, 158, 101, 62, 55, 60, 49, 51, 70, 74, 69, 66, 51, 41, 13, 
    110, 91, 71, 78, 55, 36, 61, 46, 36, 58, 69, 75, 43, 29, 31, 
    56, 59, 59, 57, 62, 57, 44, 51, 51, 72, 88, 76, 55, 20, 29, 
    48, 49, 44, 30, 21, 31, 37, 37, 37, 39, 53, 65, 48, 19, 12, 
    32, 19, 15, 10, 7, 25, 30, 24, 13, 17, 21, 27, 25, 5, 1, 
    
    -- channel=124
    69, 66, 62, 61, 70, 84, 73, 57, 52, 46, 39, 32, 27, 24, 26, 
    69, 66, 60, 56, 71, 74, 84, 82, 55, 51, 54, 52, 52, 50, 45, 
    62, 62, 41, 41, 71, 78, 85, 84, 77, 78, 73, 66, 52, 43, 33, 
    61, 69, 65, 47, 80, 89, 86, 84, 87, 77, 82, 75, 47, 45, 39, 
    103, 118, 108, 57, 70, 85, 109, 101, 92, 94, 92, 89, 67, 53, 51, 
    120, 119, 120, 56, 81, 103, 113, 102, 97, 94, 93, 98, 69, 52, 47, 
    105, 103, 110, 88, 39, 65, 95, 103, 108, 101, 92, 93, 79, 45, 37, 
    113, 116, 111, 95, 115, 80, 93, 93, 115, 116, 102, 95, 88, 67, 45, 
    128, 149, 175, 149, 136, 106, 83, 103, 115, 119, 111, 106, 96, 63, 22, 
    181, 185, 157, 142, 132, 116, 95, 103, 116, 120, 116, 112, 95, 48, 0, 
    190, 172, 131, 96, 88, 90, 85, 69, 103, 108, 101, 103, 81, 48, 18, 
    122, 104, 70, 90, 84, 75, 83, 73, 72, 97, 101, 107, 64, 35, 33, 
    69, 76, 73, 68, 60, 60, 70, 75, 86, 107, 123, 111, 76, 30, 30, 
    63, 61, 56, 37, 25, 39, 53, 54, 55, 64, 79, 97, 75, 20, 16, 
    38, 22, 17, 13, 7, 29, 38, 23, 15, 24, 32, 33, 27, 6, 0, 
    
    -- channel=125
    32, 33, 26, 28, 41, 53, 49, 33, 35, 35, 31, 30, 28, 26, 31, 
    31, 35, 30, 31, 60, 61, 70, 63, 39, 33, 40, 45, 47, 45, 44, 
    30, 30, 34, 37, 64, 79, 80, 84, 69, 57, 52, 50, 41, 34, 32, 
    33, 31, 43, 54, 74, 82, 90, 92, 86, 56, 56, 51, 36, 39, 42, 
    48, 58, 80, 68, 80, 71, 92, 101, 101, 97, 83, 73, 46, 50, 55, 
    40, 37, 49, 63, 73, 70, 84, 94, 94, 101, 106, 81, 54, 49, 50, 
    27, 27, 34, 78, 52, 53, 87, 87, 85, 95, 102, 91, 72, 40, 38, 
    32, 37, 49, 44, 82, 63, 86, 89, 90, 94, 99, 100, 75, 47, 45, 
    38, 34, 56, 95, 74, 88, 63, 98, 85, 87, 100, 104, 81, 65, 38, 
    63, 59, 41, 72, 41, 67, 54, 98, 90, 85, 96, 107, 86, 56, 40, 
    30, 40, 42, 28, 57, 59, 70, 64, 88, 84, 82, 97, 82, 57, 53, 
    7, 0, 43, 50, 73, 71, 66, 70, 61, 73, 84, 90, 74, 45, 64, 
    25, 21, 23, 40, 60, 76, 54, 72, 77, 74, 87, 85, 85, 56, 47, 
    32, 43, 44, 32, 27, 46, 59, 64, 71, 60, 53, 77, 75, 52, 47, 
    37, 27, 34, 46, 41, 46, 61, 50, 56, 57, 52, 50, 53, 48, 47, 
    
    -- channel=126
    11, 12, 23, 16, 25, 23, 14, 16, 15, 17, 16, 13, 16, 23, 18, 
    11, 11, 24, 13, 25, 33, 23, 23, 19, 23, 24, 23, 24, 30, 27, 
    13, 14, 16, 30, 21, 31, 38, 38, 32, 31, 27, 34, 32, 33, 34, 
    15, 20, 14, 20, 24, 33, 37, 46, 52, 36, 32, 32, 39, 32, 39, 
    20, 19, 13, 5, 25, 41, 32, 28, 44, 43, 43, 35, 51, 51, 54, 
    31, 25, 0, 0, 28, 42, 18, 21, 42, 42, 45, 43, 57, 67, 56, 
    25, 24, 14, 4, 35, 47, 24, 34, 37, 28, 34, 43, 48, 57, 38, 
    24, 27, 26, 6, 14, 39, 37, 42, 35, 18, 26, 37, 38, 41, 39, 
    33, 38, 21, 4, 33, 33, 47, 29, 31, 16, 22, 23, 33, 40, 61, 
    26, 36, 19, 0, 32, 16, 44, 22, 29, 21, 24, 18, 34, 44, 63, 
    25, 17, 0, 17, 24, 19, 37, 33, 36, 30, 34, 27, 38, 57, 56, 
    18, 14, 0, 20, 15, 25, 37, 31, 36, 28, 29, 32, 42, 75, 56, 
    11, 25, 24, 29, 18, 38, 51, 19, 26, 31, 23, 17, 41, 73, 66, 
    26, 34, 40, 50, 57, 52, 48, 45, 48, 51, 34, 24, 40, 70, 81, 
    44, 56, 62, 62, 75, 72, 58, 65, 72, 65, 67, 66, 65, 78, 79, 
    
    -- channel=127
    0, 0, 0, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 45, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    32, 48, 90, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 13, 
    47, 49, 53, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    26, 31, 47, 40, 16, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    29, 34, 54, 29, 43, 34, 1, 0, 0, 0, 0, 0, 0, 0, 7, 
    58, 85, 124, 133, 35, 76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    126, 147, 108, 46, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    130, 106, 65, 28, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    38, 22, 16, 8, 14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=128
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=129
    0, 41, 97, 86, 81, 94, 88, 93, 52, 22, 65, 100, 103, 108, 103, 
    0, 10, 108, 94, 78, 89, 105, 111, 115, 15, 100, 128, 126, 124, 117, 
    0, 0, 77, 99, 129, 71, 83, 124, 109, 62, 140, 162, 151, 143, 132, 
    0, 0, 97, 105, 145, 87, 37, 42, 55, 108, 142, 162, 157, 168, 172, 
    81, 105, 135, 75, 133, 133, 109, 60, 66, 98, 141, 187, 184, 149, 177, 
    144, 148, 149, 87, 128, 130, 98, 54, 62, 88, 136, 206, 195, 152, 158, 
    154, 145, 129, 116, 113, 111, 92, 80, 85, 105, 127, 195, 202, 168, 137, 
    156, 143, 67, 139, 121, 120, 96, 89, 107, 116, 126, 203, 201, 205, 177, 
    142, 131, 78, 135, 128, 115, 104, 67, 112, 88, 107, 59, 180, 175, 196, 
    147, 129, 136, 136, 161, 177, 144, 86, 66, 106, 96, 83, 69, 95, 140, 
    169, 143, 149, 139, 143, 117, 149, 152, 113, 106, 73, 90, 103, 83, 89, 
    176, 138, 164, 156, 152, 111, 122, 129, 124, 62, 92, 99, 107, 84, 58, 
    168, 150, 165, 158, 129, 90, 142, 133, 113, 73, 96, 88, 106, 84, 74, 
    159, 141, 161, 163, 100, 71, 114, 108, 90, 58, 84, 77, 60, 77, 84, 
    148, 131, 146, 163, 134, 124, 92, 84, 58, 59, 70, 74, 49, 76, 85, 
    
    -- channel=130
    0, 21, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 18, 26, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 13, 0, 0, 0, 42, 74, 67, 0, 0, 11, 0, 0, 0, 
    0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 
    0, 0, 0, 0, 0, 5, 0, 0, 1, 1, 0, 0, 0, 0, 10, 
    0, 0, 0, 0, 0, 0, 13, 11, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 25, 0, 0, 22, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 84, 20, 2, 0, 
    0, 14, 0, 0, 0, 0, 0, 0, 17, 0, 0, 0, 95, 93, 24, 
    0, 0, 0, 0, 12, 39, 0, 0, 0, 0, 7, 2, 0, 0, 35, 
    0, 0, 0, 0, 0, 0, 16, 16, 0, 0, 18, 0, 0, 8, 2, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 10, 0, 0, 0, 0, 0, 
    0, 2, 0, 0, 16, 73, 3, 12, 23, 11, 0, 8, 28, 23, 0, 
    0, 3, 10, 0, 0, 0, 0, 25, 31, 24, 0, 4, 8, 3, 0, 
    32, 0, 19, 4, 0, 0, 29, 17, 20, 3, 5, 0, 0, 0, 10, 
    
    -- channel=131
    13, 0, 0, 0, 0, 0, 0, 0, 27, 9, 0, 0, 0, 0, 0, 
    12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 
    11, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    131, 127, 23, 0, 0, 0, 21, 4, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=132
    25, 1, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 
    24, 11, 0, 0, 10, 2, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    21, 19, 0, 0, 25, 21, 13, 10, 0, 0, 18, 5, 0, 0, 0, 
    10, 5, 2, 0, 21, 19, 5, 7, 11, 13, 23, 7, 14, 20, 6, 
    0, 0, 9, 0, 24, 28, 20, 10, 15, 13, 19, 5, 16, 11, 5, 
    1, 7, 5, 0, 14, 25, 21, 14, 20, 18, 21, 12, 15, 2, 0, 
    0, 0, 2, 0, 20, 29, 28, 6, 25, 19, 27, 14, 16, 7, 0, 
    3, 0, 0, 0, 17, 20, 24, 28, 11, 19, 20, 15, 0, 20, 5, 
    3, 0, 0, 11, 15, 16, 25, 23, 9, 0, 8, 0, 22, 16, 2, 
    3, 0, 7, 8, 26, 36, 23, 15, 4, 2, 4, 0, 0, 0, 2, 
    7, 11, 11, 13, 10, 18, 24, 24, 12, 8, 0, 0, 0, 0, 0, 
    11, 8, 14, 17, 19, 0, 7, 9, 14, 0, 0, 0, 2, 0, 0, 
    10, 6, 5, 23, 23, 0, 10, 4, 5, 0, 0, 0, 11, 0, 0, 
    7, 0, 0, 21, 6, 0, 4, 0, 0, 0, 0, 0, 2, 0, 0, 
    4, 0, 0, 26, 16, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=133
    0, 12, 42, 31, 23, 38, 36, 30, 15, 0, 10, 24, 39, 39, 40, 
    0, 0, 34, 27, 2, 7, 37, 35, 22, 10, 4, 13, 19, 28, 37, 
    0, 0, 12, 8, 7, 0, 0, 15, 28, 12, 0, 0, 7, 13, 15, 
    0, 0, 0, 20, 17, 0, 0, 0, 0, 7, 8, 8, 16, 13, 10, 
    12, 12, 3, 0, 0, 0, 7, 4, 0, 4, 9, 4, 0, 0, 0, 
    6, 6, 9, 8, 11, 11, 2, 0, 0, 0, 0, 2, 0, 0, 0, 
    4, 8, 17, 14, 0, 0, 0, 16, 0, 0, 0, 7, 1, 3, 0, 
    4, 20, 24, 25, 10, 5, 0, 5, 17, 5, 17, 41, 42, 5, 4, 
    0, 0, 14, 15, 7, 0, 0, 0, 9, 16, 13, 0, 0, 17, 24, 
    0, 2, 11, 9, 0, 3, 14, 0, 0, 7, 19, 21, 16, 16, 13, 
    0, 0, 4, 2, 6, 0, 0, 4, 14, 17, 17, 14, 16, 9, 18, 
    0, 0, 0, 10, 17, 26, 16, 11, 11, 12, 14, 16, 18, 17, 12, 
    0, 1, 3, 0, 0, 11, 19, 19, 16, 16, 16, 14, 17, 20, 7, 
    2, 2, 0, 1, 5, 23, 26, 17, 16, 15, 9, 9, 9, 11, 14, 
    7, 0, 0, 7, 1, 8, 28, 28, 14, 11, 12, 12, 10, 12, 16, 
    
    -- channel=134
    14, 0, 0, 0, 0, 0, 0, 0, 0, 0, 8, 0, 0, 0, 0, 
    14, 0, 0, 5, 28, 10, 0, 0, 0, 4, 15, 0, 0, 0, 0, 
    12, 5, 0, 4, 46, 21, 0, 0, 0, 19, 20, 11, 15, 16, 9, 
    0, 29, 15, 1, 37, 41, 24, 8, 12, 30, 19, 33, 40, 21, 15, 
    20, 20, 7, 0, 33, 36, 29, 14, 19, 27, 25, 20, 26, 1, 0, 
    9, 13, 0, 6, 36, 37, 11, 24, 25, 33, 22, 25, 22, 2, 0, 
    0, 4, 0, 0, 12, 34, 29, 48, 30, 31, 30, 17, 24, 23, 13, 
    1, 3, 0, 16, 41, 27, 47, 22, 12, 30, 4, 10, 3, 14, 18, 
    0, 4, 14, 25, 42, 45, 48, 20, 12, 2, 4, 0, 0, 0, 4, 
    9, 23, 21, 23, 26, 33, 43, 37, 5, 14, 0, 0, 1, 0, 0, 
    15, 14, 26, 24, 33, 13, 19, 31, 22, 0, 0, 3, 3, 0, 0, 
    13, 6, 30, 38, 24, 22, 12, 22, 10, 0, 1, 4, 6, 1, 0, 
    8, 0, 19, 33, 0, 0, 3, 3, 0, 0, 0, 2, 0, 0, 0, 
    3, 0, 10, 36, 22, 18, 0, 0, 0, 0, 0, 0, 0, 0, 2, 
    0, 0, 12, 30, 26, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=135
    0, 0, 43, 53, 52, 44, 56, 48, 64, 58, 7, 53, 69, 68, 71, 
    0, 0, 7, 39, 54, 46, 36, 48, 55, 80, 5, 65, 69, 68, 70, 
    0, 0, 0, 44, 40, 81, 34, 20, 37, 42, 25, 43, 60, 61, 66, 
    62, 16, 0, 48, 23, 72, 73, 48, 27, 14, 46, 36, 67, 62, 44, 
    56, 33, 48, 62, 17, 53, 61, 59, 27, 22, 32, 39, 70, 71, 28, 
    49, 42, 47, 65, 28, 47, 66, 52, 37, 32, 37, 26, 62, 72, 32, 
    48, 45, 51, 53, 55, 48, 57, 29, 48, 32, 40, 33, 56, 66, 55, 
    48, 42, 89, 18, 55, 52, 48, 58, 37, 31, 49, 0, 41, 58, 53, 
    59, 36, 68, 41, 60, 62, 67, 70, 13, 62, 43, 71, 0, 35, 17, 
    52, 41, 52, 60, 44, 45, 58, 73, 80, 41, 49, 44, 52, 43, 29, 
    47, 54, 37, 61, 57, 67, 34, 52, 63, 53, 46, 38, 49, 56, 37, 
    44, 57, 23, 58, 62, 61, 54, 57, 61, 68, 27, 43, 44, 57, 53, 
    46, 41, 21, 58, 73, 61, 47, 53, 57, 53, 28, 42, 33, 43, 46, 
    47, 41, 12, 45, 74, 75, 53, 50, 49, 40, 27, 42, 45, 28, 40, 
    37, 35, 8, 33, 63, 59, 50, 38, 46, 29, 31, 36, 46, 29, 35, 
    
    -- channel=136
    0, 0, 0, 9, 0, 0, 0, 0, 30, 77, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 7, 0, 0, 0, 119, 0, 0, 0, 0, 0, 
    1, 0, 0, 0, 0, 81, 0, 0, 0, 3, 0, 0, 0, 0, 0, 
    60, 0, 0, 36, 0, 34, 45, 20, 0, 0, 0, 0, 0, 2, 0, 
    36, 0, 0, 92, 0, 0, 16, 64, 0, 0, 0, 0, 0, 56, 0, 
    0, 0, 0, 61, 0, 0, 35, 45, 0, 0, 0, 0, 0, 54, 0, 
    0, 0, 34, 0, 0, 0, 19, 0, 0, 0, 0, 0, 0, 10, 38, 
    14, 0, 83, 0, 10, 0, 15, 0, 0, 0, 0, 0, 0, 0, 0, 
    40, 0, 4, 0, 0, 0, 16, 44, 0, 42, 0, 50, 0, 0, 0, 
    20, 3, 0, 0, 0, 0, 0, 33, 42, 0, 9, 0, 0, 0, 0, 
    0, 33, 0, 0, 0, 39, 0, 0, 21, 9, 9, 0, 0, 24, 0, 
    0, 38, 0, 0, 0, 39, 0, 0, 0, 76, 0, 0, 0, 19, 25, 
    0, 17, 0, 0, 30, 30, 0, 0, 20, 39, 0, 4, 0, 1, 0, 
    10, 22, 0, 0, 42, 2, 0, 2, 19, 29, 0, 0, 21, 0, 0, 
    18, 0, 0, 0, 14, 7, 41, 0, 32, 0, 0, 0, 16, 0, 0, 
    
    -- channel=137
    0, 65, 67, 47, 44, 50, 46, 50, 38, 0, 76, 83, 67, 62, 59, 
    0, 22, 84, 63, 73, 50, 62, 68, 68, 0, 104, 79, 72, 69, 67, 
    0, 0, 92, 60, 110, 38, 51, 61, 50, 48, 99, 83, 79, 80, 76, 
    0, 27, 93, 35, 121, 68, 40, 38, 49, 93, 87, 106, 105, 82, 88, 
    27, 68, 66, 16, 110, 95, 68, 31, 50, 81, 94, 114, 94, 37, 66, 
    59, 71, 60, 26, 97, 88, 60, 35, 57, 76, 89, 117, 89, 29, 35, 
    53, 61, 46, 65, 72, 77, 55, 72, 69, 81, 82, 120, 94, 71, 40, 
    42, 64, 31, 126, 70, 81, 67, 59, 75, 69, 64, 94, 103, 83, 63, 
    26, 58, 76, 117, 84, 98, 77, 50, 83, 42, 65, 21, 92, 57, 88, 
    41, 53, 91, 82, 95, 97, 93, 75, 38, 64, 59, 53, 50, 56, 71, 
    63, 41, 95, 87, 83, 61, 97, 91, 69, 55, 42, 68, 72, 48, 45, 
    66, 33, 102, 99, 91, 72, 87, 84, 73, 25, 64, 60, 75, 44, 36, 
    56, 32, 82, 96, 68, 74, 91, 74, 57, 28, 61, 49, 62, 51, 46, 
    47, 18, 60, 96, 63, 68, 73, 55, 36, 29, 54, 43, 29, 56, 53, 
    35, 21, 40, 105, 74, 61, 35, 48, 20, 29, 44, 44, 32, 48, 55, 
    
    -- channel=138
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 7, 36, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 8, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 0, 
    0, 0, 0, 3, 0, 0, 0, 10, 0, 0, 0, 0, 0, 5, 0, 
    0, 0, 8, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 55, 36, 17, 0, 
    10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 44, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 0, 0, 0, 8, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 19, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 0, 0, 0, 
    0, 18, 0, 0, 10, 0, 0, 0, 12, 2, 0, 0, 10, 2, 0, 
    9, 22, 0, 0, 0, 0, 5, 4, 5, 0, 0, 0, 0, 0, 0, 
    28, 16, 0, 0, 0, 0, 26, 12, 12, 0, 0, 0, 0, 0, 0, 
    
    -- channel=139
    0, 1, 75, 84, 79, 77, 86, 90, 102, 48, 52, 110, 105, 105, 101, 
    0, 0, 52, 77, 110, 89, 86, 105, 104, 81, 80, 132, 122, 115, 111, 
    0, 0, 44, 74, 109, 109, 55, 49, 65, 82, 110, 126, 133, 136, 137, 
    73, 55, 97, 91, 100, 127, 106, 75, 58, 72, 124, 139, 158, 144, 137, 
    131, 119, 131, 101, 86, 115, 111, 81, 58, 72, 116, 150, 159, 144, 120, 
    133, 127, 129, 108, 104, 110, 103, 74, 79, 82, 106, 143, 169, 158, 126, 
    134, 125, 103, 104, 103, 96, 97, 83, 107, 97, 106, 146, 168, 177, 157, 
    132, 118, 95, 95, 124, 113, 106, 84, 95, 97, 105, 83, 148, 157, 153, 
    137, 105, 111, 104, 138, 147, 125, 107, 67, 92, 98, 82, 58, 99, 122, 
    152, 126, 125, 120, 120, 116, 129, 138, 104, 86, 91, 78, 87, 91, 81, 
    152, 129, 126, 135, 134, 122, 102, 111, 125, 90, 77, 87, 92, 85, 69, 
    144, 136, 120, 138, 132, 113, 119, 118, 113, 90, 73, 87, 93, 88, 80, 
    141, 132, 123, 136, 114, 60, 98, 104, 95, 72, 71, 77, 70, 76, 76, 
    135, 122, 110, 135, 134, 95, 98, 82, 69, 61, 66, 69, 63, 62, 79, 
    113, 116, 94, 125, 130, 108, 75, 66, 56, 47, 64, 68, 72, 63, 73, 
    
    -- channel=140
    1, 13, 72, 91, 88, 83, 94, 98, 108, 66, 56, 122, 110, 114, 109, 
    0, 3, 51, 79, 119, 103, 86, 110, 113, 83, 100, 149, 137, 125, 117, 
    0, 2, 56, 90, 115, 119, 72, 57, 63, 83, 143, 147, 152, 152, 153, 
    110, 81, 131, 105, 105, 130, 117, 93, 70, 83, 135, 150, 165, 159, 151, 
    141, 144, 152, 117, 105, 125, 116, 90, 67, 84, 128, 176, 181, 171, 149, 
    150, 145, 149, 116, 118, 119, 111, 83, 92, 95, 123, 165, 194, 184, 161, 
    160, 144, 117, 109, 130, 115, 110, 84, 120, 116, 122, 167, 191, 193, 186, 
    156, 131, 91, 101, 134, 127, 111, 93, 97, 111, 114, 92, 150, 180, 171, 
    166, 130, 109, 120, 143, 164, 146, 120, 84, 98, 106, 99, 86, 106, 136, 
    176, 148, 139, 135, 143, 127, 129, 148, 126, 93, 102, 81, 93, 101, 99, 
    173, 153, 139, 151, 147, 140, 121, 122, 126, 104, 78, 97, 102, 94, 76, 
    168, 159, 141, 147, 139, 110, 131, 127, 122, 94, 86, 96, 99, 93, 87, 
    166, 155, 148, 151, 130, 57, 107, 112, 102, 77, 81, 85, 79, 78, 88, 
    159, 147, 140, 150, 145, 96, 110, 89, 74, 68, 79, 78, 71, 72, 85, 
    133, 138, 123, 135, 144, 120, 78, 68, 63, 53, 73, 75, 79, 74, 81, 
    
    -- channel=141
    20, 0, 45, 56, 53, 53, 65, 63, 68, 75, 4, 54, 68, 70, 70, 
    20, 7, 15, 35, 40, 53, 42, 52, 50, 62, 28, 56, 63, 64, 64, 
    21, 16, 0, 50, 18, 54, 20, 18, 22, 29, 44, 36, 50, 57, 63, 
    84, 40, 60, 63, 0, 40, 64, 46, 27, 16, 35, 34, 51, 56, 36, 
    78, 68, 57, 61, 11, 20, 41, 43, 24, 14, 26, 41, 53, 72, 50, 
    60, 52, 55, 65, 31, 27, 31, 31, 36, 24, 26, 31, 55, 85, 72, 
    64, 52, 52, 43, 33, 18, 42, 22, 41, 24, 30, 34, 52, 68, 80, 
    70, 47, 61, 16, 53, 33, 26, 49, 18, 37, 40, 13, 26, 57, 58, 
    77, 39, 38, 37, 38, 45, 47, 41, 19, 45, 45, 60, 7, 26, 32, 
    72, 62, 39, 45, 28, 22, 24, 39, 72, 45, 39, 38, 52, 52, 30, 
    59, 67, 25, 45, 49, 47, 18, 26, 38, 51, 31, 44, 42, 41, 46, 
    57, 69, 26, 36, 43, 34, 45, 41, 44, 49, 40, 39, 35, 52, 44, 
    61, 67, 37, 33, 40, 6, 34, 37, 38, 46, 33, 37, 29, 27, 43, 
    63, 73, 41, 32, 46, 62, 43, 37, 42, 33, 35, 39, 41, 28, 42, 
    51, 67, 50, 16, 42, 50, 43, 34, 44, 39, 34, 40, 43, 44, 30, 
    
    -- channel=142
    23, 88, 94, 63, 63, 70, 70, 67, 43, 20, 75, 75, 77, 77, 77, 
    23, 65, 110, 58, 42, 35, 57, 64, 54, 2, 95, 52, 59, 67, 71, 
    23, 43, 108, 59, 55, 7, 43, 65, 54, 36, 66, 43, 40, 42, 41, 
    9, 28, 76, 29, 71, 10, 19, 31, 42, 64, 48, 51, 32, 30, 42, 
    9, 52, 40, 8, 71, 34, 24, 17, 41, 53, 46, 61, 28, 8, 47, 
    33, 39, 38, 20, 54, 33, 29, 15, 40, 47, 49, 60, 28, 7, 29, 
    34, 41, 39, 66, 41, 29, 18, 30, 27, 40, 38, 65, 32, 20, 11, 
    25, 47, 41, 91, 19, 40, 10, 41, 48, 30, 49, 55, 68, 31, 25, 
    17, 40, 42, 69, 24, 30, 17, 12, 57, 38, 52, 50, 80, 46, 63, 
    14, 24, 48, 38, 38, 36, 30, 14, 31, 52, 46, 60, 56, 52, 76, 
    25, 17, 48, 38, 33, 23, 56, 40, 23, 44, 48, 57, 58, 38, 48, 
    29, 12, 55, 35, 40, 26, 59, 42, 41, 22, 66, 47, 57, 39, 42, 
    26, 17, 47, 37, 35, 52, 70, 48, 41, 35, 65, 44, 53, 49, 48, 
    25, 23, 43, 39, 13, 50, 56, 55, 43, 40, 59, 48, 38, 63, 50, 
    26, 31, 31, 54, 25, 36, 35, 60, 41, 57, 52, 52, 42, 55, 57, 
    
    -- channel=143
    0, 0, 27, 48, 42, 34, 39, 33, 53, 35, 0, 46, 52, 48, 52, 
    0, 0, 10, 30, 63, 49, 50, 42, 66, 77, 0, 67, 67, 63, 65, 
    0, 0, 0, 13, 63, 104, 45, 44, 67, 30, 26, 68, 86, 79, 75, 
    0, 0, 0, 56, 50, 102, 49, 45, 25, 0, 79, 48, 97, 107, 67, 
    63, 4, 59, 69, 23, 85, 97, 79, 28, 13, 58, 53, 100, 94, 32, 
    66, 52, 73, 52, 47, 82, 93, 50, 33, 16, 51, 59, 100, 95, 37, 
    62, 54, 80, 54, 57, 54, 90, 37, 69, 41, 45, 53, 94, 103, 62, 
    68, 55, 92, 39, 87, 70, 86, 51, 54, 40, 65, 62, 69, 111, 64, 
    79, 40, 82, 41, 86, 82, 77, 104, 11, 46, 69, 28, 21, 84, 39, 
    78, 41, 70, 78, 71, 97, 97, 87, 48, 40, 75, 42, 19, 54, 30, 
    75, 72, 60, 76, 79, 93, 56, 78, 103, 80, 33, 35, 52, 63, 44, 
    70, 83, 39, 97, 102, 99, 56, 71, 84, 77, 9, 51, 58, 57, 42, 
    70, 66, 30, 89, 123, 45, 71, 72, 84, 55, 24, 44, 55, 47, 41, 
    71, 55, 13, 82, 106, 37, 73, 58, 58, 25, 24, 32, 42, 9, 39, 
    58, 46, 7, 68, 91, 86, 71, 42, 48, 0, 22, 30, 28, 19, 35, 
    
    -- channel=144
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=145
    157, 158, 156, 127, 116, 99, 100, 118, 164, 178, 180, 177, 131, 154, 121, 
    182, 182, 174, 101, 110, 121, 134, 161, 182, 184, 179, 184, 186, 169, 179, 
    194, 195, 164, 34, 31, 32, 24, 18, 41, 88, 160, 172, 173, 148, 190, 
    193, 192, 158, 49, 85, 88, 79, 79, 63, 53, 104, 198, 144, 125, 135, 
    193, 182, 153, 40, 75, 97, 76, 67, 81, 86, 76, 143, 172, 129, 101, 
    192, 178, 78, 10, 55, 46, 48, 57, 59, 75, 103, 117, 197, 193, 194, 
    161, 133, 113, 13, 8, 42, 25, 11, 31, 50, 34, 98, 177, 201, 193, 
    135, 77, 82, 70, 44, 9, 23, 23, 32, 21, 23, 44, 64, 99, 196, 
    102, 14, 96, 41, 25, 54, 13, 0, 0, 0, 0, 0, 18, 56, 160, 
    119, 30, 77, 0, 40, 9, 47, 88, 73, 102, 92, 90, 111, 37, 134, 
    136, 1, 6, 0, 0, 4, 0, 13, 45, 34, 26, 34, 37, 21, 102, 
    124, 15, 32, 0, 0, 0, 75, 0, 75, 41, 42, 113, 0, 63, 100, 
    103, 0, 15, 56, 0, 0, 0, 0, 0, 70, 61, 22, 0, 0, 86, 
    107, 94, 39, 48, 14, 0, 0, 0, 2, 102, 113, 40, 0, 11, 80, 
    93, 73, 41, 17, 14, 0, 0, 0, 0, 19, 59, 15, 0, 5, 85, 
    
    -- channel=146
    0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 32, 62, 77, 107, 132, 109, 67, 31, 0, 0, 2, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 51, 28, 0, 0, 23, 31, 
    0, 0, 13, 7, 0, 0, 0, 14, 0, 0, 0, 56, 0, 0, 0, 
    0, 0, 49, 58, 0, 35, 49, 6, 9, 7, 0, 0, 0, 0, 0, 
    17, 5, 0, 0, 63, 22, 20, 34, 48, 40, 58, 48, 20, 0, 0, 
    14, 53, 55, 0, 0, 0, 0, 0, 0, 0, 11, 43, 97, 96, 0, 
    0, 83, 16, 0, 37, 40, 53, 47, 72, 74, 65, 75, 88, 73, 36, 
    0, 0, 0, 119, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 17, 54, 12, 32, 42, 73, 73, 55, 101, 106, 99, 73, 77, 31, 
    0, 0, 0, 0, 20, 32, 0, 0, 54, 19, 28, 0, 43, 0, 0, 
    10, 53, 28, 0, 0, 17, 108, 79, 28, 15, 0, 17, 60, 86, 53, 
    10, 0, 0, 0, 0, 0, 1, 2, 6, 0, 0, 0, 9, 0, 0, 
    0, 13, 0, 3, 0, 0, 0, 0, 0, 65, 108, 41, 19, 0, 0, 
    19, 2, 0, 30, 9, 0, 0, 0, 0, 13, 41, 33, 0, 0, 0, 
    
    -- channel=147
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 12, 21, 23, 31, 7, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 47, 125, 101, 94, 136, 75, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 5, 0, 0, 0, 45, 0, 0, 0, 2, 45, 0, 0, 0, 
    0, 0, 0, 38, 9, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 58, 37, 0, 8, 12, 0, 4, 8, 0, 0, 0, 0, 11, 0, 
    0, 0, 0, 0, 0, 0, 26, 16, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 21, 19, 6, 0, 0, 0, 7, 8, 3, 
    
    -- channel=148
    25, 20, 31, 25, 17, 23, 16, 16, 22, 27, 24, 22, 18, 20, 12, 
    33, 32, 38, 36, 48, 56, 57, 61, 53, 31, 21, 26, 26, 22, 11, 
    39, 40, 36, 42, 80, 90, 82, 84, 89, 83, 25, 26, 28, 16, 11, 
    38, 41, 40, 57, 84, 63, 85, 106, 97, 93, 73, 35, 19, 16, 9, 
    37, 41, 45, 69, 88, 100, 92, 106, 104, 96, 87, 45, 22, 17, 8, 
    35, 43, 34, 82, 87, 88, 104, 103, 101, 106, 106, 75, 51, 38, 39, 
    38, 38, 38, 52, 64, 93, 96, 85, 83, 81, 58, 54, 53, 43, 36, 
    23, 31, 16, 30, 88, 84, 91, 92, 82, 75, 85, 76, 66, 77, 52, 
    19, 21, 28, 44, 66, 56, 45, 35, 30, 23, 20, 21, 47, 68, 47, 
    30, 42, 36, 30, 63, 57, 66, 64, 62, 81, 79, 75, 73, 67, 56, 
    35, 32, 43, 39, 48, 49, 44, 71, 60, 79, 77, 63, 78, 59, 49, 
    50, 49, 32, 45, 40, 41, 69, 43, 50, 32, 45, 65, 32, 69, 46, 
    67, 40, 42, 63, 43, 40, 32, 34, 38, 32, 28, 45, 43, 32, 48, 
    64, 68, 67, 56, 57, 40, 28, 32, 30, 61, 65, 70, 31, 38, 56, 
    75, 71, 66, 57, 56, 41, 31, 36, 42, 52, 64, 63, 33, 39, 57, 
    
    -- channel=149
    0, 0, 0, 0, 7, 17, 20, 15, 10, 3, 0, 3, 0, 0, 0, 
    0, 0, 3, 8, 7, 1, 3, 14, 25, 23, 0, 1, 1, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 2, 3, 3, 
    0, 0, 0, 0, 0, 24, 0, 0, 0, 0, 0, 0, 0, 3, 11, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 0, 0, 
    8, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    5, 1, 0, 0, 0, 0, 0, 0, 0, 11, 2, 0, 8, 21, 10, 
    20, 1, 12, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    8, 13, 6, 0, 0, 12, 20, 0, 0, 0, 0, 0, 0, 0, 19, 
    0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 11, 32, 0, 8, 9, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 22, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=150
    51, 45, 49, 37, 48, 55, 63, 65, 52, 48, 38, 42, 45, 35, 31, 
    64, 61, 57, 64, 63, 72, 71, 65, 59, 33, 29, 37, 39, 14, 32, 
    63, 62, 62, 64, 111, 120, 131, 121, 113, 75, 56, 44, 32, 2, 15, 
    62, 57, 62, 97, 129, 128, 126, 139, 139, 148, 57, 43, 37, 32, 4, 
    58, 58, 73, 106, 114, 115, 130, 137, 130, 135, 116, 77, 57, 49, 59, 
    52, 53, 78, 94, 87, 114, 123, 115, 105, 106, 109, 59, 65, 62, 62, 
    42, 38, 37, 83, 131, 128, 125, 114, 127, 116, 75, 72, 52, 68, 52, 
    30, 23, 46, 57, 107, 65, 86, 73, 59, 55, 60, 50, 58, 79, 64, 
    52, 58, 21, 47, 81, 91, 89, 77, 85, 98, 81, 77, 100, 104, 67, 
    53, 51, 28, 47, 65, 54, 53, 92, 53, 80, 70, 68, 83, 66, 81, 
    60, 66, 30, 48, 41, 58, 80, 56, 52, 65, 60, 64, 78, 78, 86, 
    78, 44, 54, 67, 43, 32, 37, 31, 61, 53, 69, 64, 36, 38, 82, 
    90, 82, 80, 61, 57, 37, 28, 31, 43, 90, 88, 61, 37, 48, 95, 
    98, 87, 74, 60, 66, 35, 30, 40, 54, 39, 69, 45, 33, 57, 96, 
    100, 97, 83, 61, 55, 42, 39, 42, 47, 55, 61, 55, 34, 50, 99, 
    
    -- channel=151
    64, 63, 70, 64, 45, 46, 38, 44, 46, 57, 58, 53, 73, 47, 57, 
    67, 67, 69, 61, 20, 17, 22, 17, 13, 32, 39, 50, 60, 63, 36, 
    70, 69, 73, 105, 22, 43, 47, 54, 37, 26, 12, 51, 67, 59, 15, 
    70, 71, 74, 83, 4, 35, 61, 41, 47, 38, 44, 25, 72, 64, 37, 
    69, 73, 55, 72, 5, 32, 47, 33, 34, 41, 54, 17, 56, 84, 74, 
    56, 70, 89, 75, 0, 33, 36, 27, 28, 33, 19, 32, 36, 71, 69, 
    58, 72, 53, 77, 21, 28, 38, 30, 13, 17, 34, 5, 8, 26, 64, 
    65, 71, 30, 60, 42, 59, 35, 29, 7, 11, 13, 0, 0, 23, 18, 
    73, 81, 23, 44, 25, 11, 39, 54, 46, 39, 62, 44, 28, 35, 4, 
    81, 86, 0, 53, 0, 31, 8, 2, 46, 26, 37, 30, 18, 52, 0, 
    67, 93, 26, 32, 17, 0, 24, 41, 12, 50, 42, 42, 36, 34, 8, 
    63, 94, 0, 38, 42, 0, 0, 37, 0, 32, 27, 6, 71, 0, 0, 
    57, 105, 26, 30, 48, 20, 0, 0, 0, 0, 48, 66, 27, 0, 0, 
    52, 57, 67, 23, 25, 39, 0, 0, 0, 0, 23, 66, 25, 0, 0, 
    50, 53, 59, 29, 18, 24, 9, 8, 7, 11, 13, 37, 26, 0, 0, 
    
    -- channel=152
    0, 0, 0, 46, 0, 0, 0, 0, 0, 0, 0, 0, 27, 0, 36, 
    0, 0, 0, 125, 0, 0, 0, 0, 0, 0, 0, 0, 0, 24, 0, 
    0, 0, 25, 188, 0, 0, 0, 11, 0, 0, 0, 0, 0, 36, 0, 
    0, 0, 26, 168, 0, 0, 43, 0, 0, 0, 0, 0, 13, 18, 0, 
    0, 0, 67, 134, 0, 0, 34, 0, 0, 0, 0, 0, 0, 33, 0, 
    0, 10, 91, 118, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 50, 13, 98, 0, 0, 11, 5, 0, 0, 21, 0, 0, 0, 0, 
    0, 109, 0, 38, 15, 26, 0, 5, 0, 0, 0, 0, 0, 0, 0, 
    19, 138, 0, 139, 0, 0, 16, 56, 0, 0, 33, 0, 0, 0, 0, 
    27, 169, 0, 113, 0, 27, 0, 0, 13, 0, 7, 0, 0, 74, 0, 
    0, 200, 0, 31, 17, 0, 0, 42, 0, 19, 0, 0, 51, 0, 0, 
    0, 205, 0, 0, 81, 0, 0, 100, 0, 23, 0, 0, 170, 0, 0, 
    0, 130, 0, 0, 68, 43, 0, 0, 0, 0, 0, 61, 72, 0, 0, 
    0, 13, 58, 0, 1, 76, 0, 0, 0, 0, 0, 70, 72, 0, 0, 
    1, 6, 30, 47, 0, 36, 5, 0, 0, 0, 0, 27, 62, 0, 0, 
    
    -- channel=153
    96, 98, 99, 62, 74, 88, 86, 90, 112, 101, 90, 102, 73, 78, 50, 
    122, 122, 105, 43, 85, 100, 97, 102, 108, 96, 78, 110, 105, 60, 82, 
    127, 128, 108, 5, 107, 119, 109, 99, 109, 101, 109, 122, 90, 44, 82, 
    127, 121, 106, 30, 139, 140, 109, 124, 123, 125, 114, 121, 95, 57, 61, 
    129, 115, 85, 38, 137, 126, 100, 128, 129, 125, 114, 146, 129, 93, 86, 
    135, 106, 65, 39, 107, 106, 99, 105, 108, 113, 121, 133, 152, 127, 129, 
    131, 88, 88, 43, 93, 113, 99, 87, 98, 105, 62, 91, 128, 125, 134, 
    110, 38, 96, 63, 84, 72, 68, 45, 53, 58, 38, 53, 101, 120, 177, 
    92, 16, 106, 22, 77, 73, 78, 61, 54, 68, 53, 47, 99, 100, 181, 
    98, 0, 83, 0, 81, 39, 70, 86, 98, 99, 90, 93, 103, 52, 157, 
    110, 0, 47, 20, 17, 49, 77, 32, 100, 66, 67, 100, 55, 72, 147, 
    118, 0, 65, 56, 0, 16, 59, 0, 85, 55, 81, 96, 0, 78, 120, 
    127, 27, 71, 85, 15, 0, 0, 11, 31, 115, 96, 37, 1, 37, 140, 
    120, 109, 60, 71, 51, 0, 0, 13, 37, 119, 100, 33, 0, 55, 137, 
    117, 105, 70, 47, 46, 14, 11, 21, 35, 56, 85, 49, 0, 48, 140, 
    
    -- channel=154
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 33, 30, 14, 14, 46, 54, 41, 9, 0, 0, 6, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 0, 
    0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 
    0, 0, 27, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 12, 0, 0, 0, 0, 0, 0, 0, 10, 7, 0, 22, 14, 0, 
    4, 20, 0, 9, 0, 0, 0, 0, 33, 23, 0, 49, 13, 0, 0, 
    0, 0, 0, 34, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 23, 0, 0, 0, 0, 0, 23, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 26, 0, 0, 0, 0, 21, 36, 0, 31, 0, 13, 40, 20, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 5, 0, 0, 
    0, 0, 0, 4, 0, 0, 0, 0, 0, 17, 0, 24, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 0, 0, 0, 
    
    -- channel=155
    157, 157, 149, 117, 110, 120, 143, 155, 164, 163, 155, 156, 165, 150, 151, 
    171, 171, 162, 102, 67, 59, 56, 67, 82, 110, 135, 144, 151, 143, 145, 
    167, 166, 159, 94, 62, 82, 82, 85, 71, 63, 100, 157, 142, 125, 120, 
    167, 163, 144, 103, 57, 114, 108, 86, 91, 100, 106, 110, 153, 137, 112, 
    164, 163, 107, 70, 59, 65, 75, 74, 80, 87, 103, 110, 158, 173, 156, 
    141, 147, 118, 72, 26, 52, 51, 48, 51, 56, 64, 93, 128, 169, 167, 
    119, 112, 78, 79, 68, 57, 62, 46, 47, 61, 49, 43, 73, 105, 161, 
    104, 62, 66, 76, 41, 35, 14, 8, 0, 3, 0, 0, 24, 50, 116, 
    120, 79, 60, 41, 39, 45, 79, 87, 83, 98, 115, 93, 88, 73, 106, 
    131, 64, 32, 26, 14, 25, 10, 16, 76, 42, 52, 49, 49, 46, 64, 
    123, 85, 40, 24, 0, 8, 53, 22, 34, 45, 38, 64, 34, 56, 71, 
    113, 53, 23, 65, 31, 0, 0, 15, 0, 64, 73, 48, 37, 10, 37, 
    105, 108, 58, 61, 43, 9, 0, 0, 8, 73, 130, 97, 14, 14, 47, 
    93, 98, 74, 50, 37, 25, 2, 5, 15, 39, 57, 68, 3, 8, 52, 
    93, 89, 78, 40, 28, 23, 14, 14, 15, 20, 26, 48, 12, 11, 59, 
    
    -- channel=156
    177, 181, 168, 134, 118, 119, 145, 165, 183, 182, 175, 170, 176, 175, 167, 
    184, 185, 173, 100, 65, 57, 58, 64, 76, 118, 155, 159, 170, 168, 165, 
    183, 181, 170, 107, 62, 91, 89, 95, 83, 73, 113, 175, 159, 139, 145, 
    183, 180, 156, 102, 58, 109, 117, 83, 91, 97, 120, 122, 163, 153, 133, 
    178, 176, 121, 56, 63, 68, 65, 73, 78, 86, 104, 117, 169, 188, 173, 
    146, 155, 114, 76, 36, 57, 54, 44, 50, 57, 62, 97, 140, 184, 183, 
    127, 116, 79, 70, 62, 51, 43, 39, 31, 46, 50, 56, 88, 106, 166, 
    111, 68, 55, 89, 45, 59, 46, 20, 1, 9, 0, 0, 21, 49, 122, 
    121, 75, 68, 41, 35, 40, 62, 90, 91, 101, 124, 110, 103, 77, 111, 
    136, 71, 34, 20, 25, 23, 27, 12, 76, 51, 54, 54, 53, 47, 70, 
    128, 82, 45, 28, 14, 16, 57, 46, 44, 70, 54, 85, 61, 44, 85, 
    112, 57, 23, 63, 39, 6, 0, 1, 1, 44, 72, 53, 21, 28, 39, 
    102, 99, 76, 66, 42, 20, 0, 3, 15, 68, 135, 99, 20, 16, 61, 
    101, 100, 72, 57, 37, 26, 12, 11, 16, 54, 52, 65, 5, 15, 60, 
    94, 89, 81, 46, 32, 24, 23, 23, 25, 29, 35, 42, 21, 21, 68, 
    
    -- channel=157
    45, 46, 42, 42, 31, 33, 44, 62, 48, 43, 49, 34, 59, 62, 60, 
    35, 35, 42, 35, 0, 0, 0, 0, 0, 1, 28, 31, 35, 58, 46, 
    27, 27, 27, 51, 0, 0, 0, 0, 0, 0, 0, 29, 47, 52, 32, 
    27, 29, 20, 31, 0, 0, 0, 0, 0, 0, 0, 0, 31, 71, 46, 
    24, 32, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 26, 46, 63, 
    9, 31, 31, 17, 0, 0, 0, 0, 0, 0, 0, 0, 0, 27, 26, 
    9, 12, 1, 13, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 13, 
    17, 15, 0, 39, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    39, 49, 5, 0, 0, 1, 0, 4, 50, 49, 55, 55, 34, 3, 0, 
    26, 50, 0, 31, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    16, 51, 13, 9, 3, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 
    0, 38, 0, 21, 31, 5, 0, 0, 0, 0, 2, 2, 13, 0, 0, 
    0, 41, 28, 0, 13, 29, 9, 2, 0, 7, 41, 51, 15, 0, 0, 
    0, 0, 6, 0, 0, 22, 16, 12, 9, 0, 0, 12, 16, 0, 0, 
    0, 0, 4, 0, 0, 7, 14, 8, 0, 0, 0, 0, 23, 0, 0, 
    
    -- channel=158
    18, 26, 24, 6, 24, 26, 21, 28, 38, 21, 23, 29, 10, 24, 11, 
    21, 23, 15, 0, 27, 32, 24, 26, 36, 35, 24, 45, 30, 13, 34, 
    22, 24, 6, 0, 14, 0, 0, 0, 0, 28, 36, 41, 28, 23, 46, 
    22, 23, 10, 0, 29, 3, 0, 0, 0, 0, 37, 50, 21, 11, 44, 
    27, 17, 0, 0, 26, 11, 0, 0, 0, 0, 0, 36, 39, 9, 16, 
    46, 17, 0, 0, 20, 0, 0, 0, 0, 8, 0, 35, 48, 22, 24, 
    55, 16, 31, 0, 5, 0, 0, 0, 0, 5, 2, 34, 53, 31, 42, 
    48, 8, 48, 10, 5, 1, 0, 0, 11, 13, 5, 25, 45, 38, 65, 
    21, 0, 79, 0, 30, 5, 6, 0, 6, 7, 0, 3, 28, 3, 70, 
    18, 0, 49, 0, 35, 9, 30, 22, 30, 19, 12, 20, 19, 0, 70, 
    26, 0, 35, 11, 9, 15, 19, 0, 45, 0, 13, 32, 0, 25, 50, 
    19, 0, 28, 22, 0, 26, 44, 0, 58, 17, 23, 38, 0, 39, 57, 
    14, 0, 18, 26, 0, 0, 19, 24, 23, 56, 10, 0, 0, 26, 65, 
    14, 4, 0, 11, 10, 0, 18, 22, 30, 70, 27, 0, 0, 39, 49, 
    4, 2, 0, 0, 15, 0, 15, 20, 22, 26, 34, 0, 0, 36, 60, 
    
    -- channel=159
    98, 84, 110, 97, 78, 68, 65, 56, 75, 103, 93, 94, 96, 65, 66, 
    120, 117, 137, 130, 98, 102, 99, 118, 119, 95, 83, 87, 106, 98, 57, 
    126, 125, 146, 130, 56, 75, 74, 83, 87, 72, 52, 94, 110, 95, 39, 
    126, 134, 116, 172, 49, 98, 122, 117, 108, 95, 74, 84, 107, 97, 47, 
    123, 138, 143, 143, 65, 89, 129, 100, 102, 96, 129, 69, 97, 128, 71, 
    109, 150, 105, 116, 34, 79, 92, 86, 87, 77, 94, 63, 80, 126, 125, 
    96, 142, 87, 92, 46, 79, 109, 72, 66, 95, 65, 46, 84, 112, 114, 
    117, 104, 31, 109, 79, 58, 50, 53, 35, 31, 34, 23, 26, 65, 81, 
    107, 88, 25, 93, 27, 47, 46, 55, 3, 0, 53, 3, 0, 72, 39, 
    121, 110, 50, 26, 26, 44, 28, 33, 98, 83, 104, 90, 109, 79, 0, 
    114, 126, 12, 32, 0, 0, 3, 50, 8, 59, 45, 24, 67, 34, 0, 
    129, 130, 20, 31, 32, 0, 0, 56, 0, 56, 56, 71, 63, 35, 0, 
    113, 108, 18, 83, 53, 9, 0, 0, 0, 0, 76, 121, 19, 0, 0, 
    102, 123, 100, 87, 44, 37, 0, 0, 0, 26, 81, 146, 7, 0, 0, 
    113, 106, 108, 65, 32, 27, 0, 0, 0, 12, 33, 97, 3, 0, 0, 
    
    
    others => 0);
end gold_package;
