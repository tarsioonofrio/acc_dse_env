library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
package gold_package is
  type mem is array(0 to 4000000) of integer;

  constant gold : mem := (

    -- gold
    -- channel=0
    339, 337, 348, 352, 355, 322, 362, 390, 368, 304, 254, 262, 281, 302, 312, 
    353, 356, 360, 363, 357, 294, 317, 310, 241, 141, 76, 96, 152, 248, 302, 
    244, 288, 365, 373, 377, 295, 209, 136, 86, 49, 20, 27, 49, 126, 241, 
    79, 153, 340, 365, 315, 226, 127, 60, 46, 64, 64, 60, 40, 50, 177, 
    1, 64, 285, 279, 133, 99, 62, 46, 37, 57, 61, 53, 48, 39, 101, 
    0, 23, 257, 258, 61, 65, 66, 61, 41, 55, 49, 39, 44, 35, 31, 
    0, 1, 183, 288, 126, 99, 70, 64, 38, 44, 30, 31, 33, 34, 54, 
    0, 0, 50, 193, 149, 75, 46, 52, 63, 102, 53, 34, 27, 61, 153, 
    0, 0, 0, 39, 121, 64, 75, 66, 61, 145, 87, 51, 50, 126, 251, 
    4, 0, 0, 0, 16, 58, 55, 36, 37, 88, 48, 17, 43, 219, 280, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 26, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=1
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    12, 10, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 
    37, 31, 24, 24, 25, 26, 24, 24, 37, 35, 29, 19, 25, 24, 12, 
    43, 34, 32, 25, 32, 33, 59, 97, 93, 61, 60, 59, 47, 30, 10, 
    55, 63, 54, 44, 43, 38, 50, 62, 70, 89, 77, 58, 46, 30, 9, 
    
    -- channel=2
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 11, 0, 0, 0, 0, 0, 0, 0, 0, 14, 1, 
    0, 0, 5, 21, 46, 29, 25, 4, 0, 0, 0, 0, 0, 33, 47, 
    0, 0, 0, 0, 11, 11, 0, 0, 0, 0, 0, 0, 8, 28, 24, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 46, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 11, 14, 37, 1, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 17, 6, 0, 6, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 18, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    -- channel=3
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 9, 7, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 16, 16, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 15, 24, 27, 28, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    28, 4, 4, 21, 42, 30, 23, 31, 40, 45, 44, 43, 41, 40, 41, 
    50, 32, 30, 42, 47, 36, 36, 52, 51, 50, 52, 62, 46, 37, 53, 
    
    -- channel=4
    79, 78, 94, 75, 58, 91, 107, 96, 141, 139, 112, 111, 137, 109, 93, 
    79, 97, 103, 72, 61, 96, 88, 100, 115, 113, 117, 111, 134, 95, 96, 
    89, 108, 86, 59, 63, 102, 122, 115, 99, 91, 122, 119, 125, 111, 107, 
    83, 106, 85, 70, 80, 161, 187, 120, 108, 79, 138, 173, 122, 102, 77, 
    82, 103, 81, 84, 120, 156, 137, 113, 156, 158, 177, 199, 151, 85, 57, 
    79, 98, 93, 82, 152, 140, 103, 123, 162, 172, 165, 173, 167, 79, 76, 
    76, 93, 97, 103, 140, 153, 136, 132, 120, 119, 103, 136, 149, 116, 84, 
    90, 95, 90, 99, 104, 113, 130, 134, 134, 129, 114, 89, 102, 117, 75, 
    89, 108, 89, 100, 101, 77, 103, 105, 118, 120, 127, 114, 85, 103, 90, 
    84, 96, 95, 103, 104, 80, 92, 83, 98, 101, 104, 118, 91, 75, 102, 
    82, 114, 114, 94, 112, 97, 96, 93, 76, 89, 101, 115, 115, 82, 97, 
    90, 147, 189, 137, 96, 102, 109, 116, 84, 80, 102, 119, 158, 130, 123, 
    118, 159, 207, 229, 170, 106, 113, 116, 91, 87, 95, 104, 127, 131, 147, 
    101, 152, 202, 211, 240, 214, 184, 127, 103, 100, 101, 113, 103, 121, 145, 
    115, 130, 168, 225, 201, 228, 235, 211, 151, 106, 100, 109, 106, 116, 186, 
    
    -- channel=5
    194, 201, 207, 204, 221, 223, 211, 189, 146, 112, 102, 107, 104, 105, 93, 
    200, 226, 223, 218, 232, 237, 238, 224, 199, 121, 102, 108, 115, 120, 110, 
    187, 209, 226, 237, 236, 250, 246, 242, 235, 166, 143, 129, 120, 124, 120, 
    168, 201, 225, 232, 239, 255, 235, 232, 221, 217, 202, 166, 122, 122, 120, 
    158, 189, 223, 239, 247, 237, 177, 175, 175, 194, 194, 165, 125, 124, 120, 
    136, 184, 206, 226, 235, 209, 124, 120, 149, 148, 138, 114, 107, 124, 120, 
    122, 175, 182, 185, 184, 181, 155, 116, 113, 121, 107, 74, 85, 124, 114, 
    125, 146, 163, 167, 166, 167, 193, 149, 123, 123, 106, 75, 83, 122, 104, 
    139, 136, 144, 151, 157, 154, 155, 168, 145, 130, 101, 75, 86, 124, 86, 
    138, 139, 113, 115, 111, 145, 133, 149, 143, 92, 65, 76, 91, 132, 76, 
    137, 137, 117, 102, 81, 85, 90, 120, 109, 84, 66, 76, 96, 127, 93, 
    136, 130, 129, 134, 135, 103, 118, 109, 74, 58, 46, 61, 85, 115, 120, 
    148, 138, 139, 148, 163, 137, 118, 119, 87, 69, 54, 64, 87, 90, 111, 
    128, 125, 136, 140, 128, 134, 132, 135, 120, 106, 115, 122, 124, 128, 110, 
    130, 131, 132, 138, 134, 141, 157, 140, 143, 125, 145, 152, 145, 145, 130, 
    
    -- channel=6
    422, 440, 462, 476, 453, 405, 389, 364, 315, 244, 247, 198, 89, 84, 165, 
    417, 388, 368, 342, 310, 282, 278, 271, 247, 228, 207, 148, 59, 93, 175, 
    281, 257, 248, 238, 235, 220, 223, 237, 229, 222, 126, 42, 99, 151, 190, 
    199, 201, 205, 206, 217, 215, 212, 230, 232, 209, 70, 44, 149, 201, 196, 
    182, 197, 200, 201, 203, 208, 202, 187, 172, 114, 12, 52, 144, 182, 188, 
    195, 194, 199, 200, 182, 135, 82, 61, 53, 0, 0, 7, 57, 105, 162, 
    201, 193, 191, 177, 126, 55, 0, 0, 9, 0, 0, 0, 14, 30, 91, 
    193, 190, 151, 90, 37, 31, 10, 0, 4, 0, 0, 0, 0, 23, 23, 
    184, 156, 68, 0, 0, 20, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    162, 71, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    126, 0, 0, 0, 6, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    107, 0, 0, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 22, 
    76, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 41, 
    71, 3, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 15, 8, 29, 
    63, 12, 0, 0, 0, 0, 0, 0, 10, 8, 0, 13, 29, 32, 34, 
    
    -- channel=7
    41, 44, 43, 38, 101, 141, 96, 57, 51, 58, 51, 45, 45, 42, 41, 
    42, 44, 53, 70, 154, 209, 205, 175, 87, 66, 76, 71, 69, 58, 55, 
    48, 48, 59, 104, 200, 261, 292, 299, 194, 94, 93, 93, 78, 62, 67, 
    59, 57, 50, 131, 250, 277, 296, 321, 301, 202, 155, 138, 74, 68, 91, 
    54, 54, 70, 141, 246, 243, 258, 299, 340, 330, 298, 236, 127, 112, 125, 
    49, 47, 53, 110, 204, 230, 252, 286, 307, 336, 351, 304, 193, 136, 118, 
    38, 38, 43, 67, 143, 214, 265, 300, 274, 277, 323, 323, 234, 131, 85, 
    52, 50, 62, 79, 102, 144, 227, 292, 276, 264, 313, 328, 259, 159, 97, 
    65, 54, 47, 93, 125, 124, 168, 269, 277, 262, 298, 324, 281, 193, 130, 
    29, 26, 26, 74, 147, 149, 181, 269, 283, 266, 288, 322, 291, 182, 118, 
    0, 3, 54, 134, 201, 230, 245, 244, 284, 276, 276, 308, 272, 169, 126, 
    18, 16, 39, 102, 175, 265, 224, 160, 234, 264, 242, 266, 240, 174, 143, 
    47, 54, 53, 73, 104, 158, 203, 194, 227, 251, 218, 251, 243, 186, 157, 
    71, 85, 113, 123, 126, 131, 163, 201, 233, 231, 216, 252, 253, 191, 169, 
    99, 116, 138, 144, 143, 147, 165, 175, 180, 182, 195, 203, 199, 177, 154, 
    
    -- channel=8
    10, 67, 160, 139, 120, 164, 170, 162, 116, 70, 69, 133, 168, 181, 181, 
    13, 43, 148, 106, 24, 78, 104, 123, 105, 61, 81, 116, 137, 154, 159, 
    17, 24, 124, 110, 0, 10, 53, 83, 83, 58, 74, 97, 96, 100, 110, 
    61, 50, 105, 114, 11, 0, 30, 47, 46, 42, 52, 74, 43, 67, 96, 
    114, 110, 107, 107, 28, 6, 22, 33, 32, 30, 58, 99, 75, 124, 147, 
    119, 106, 120, 105, 43, 12, 24, 25, 21, 20, 46, 101, 95, 144, 181, 
    146, 125, 129, 104, 47, 13, 14, 13, 21, 23, 36, 98, 100, 108, 147, 
    147, 118, 90, 79, 40, 23, 1, 13, 48, 62, 63, 114, 117, 105, 121, 
    145, 113, 53, 52, 26, 17, 2, 12, 79, 80, 79, 113, 119, 120, 143, 
    140, 114, 60, 53, 52, 25, 6, 10, 58, 77, 86, 107, 94, 102, 122, 
    123, 107, 63, 59, 62, 55, 51, 31, 42, 84, 90, 89, 74, 79, 91, 
    123, 121, 72, 33, 44, 53, 71, 56, 59, 84, 100, 80, 69, 80, 85, 
    129, 155, 111, 33, 41, 44, 76, 82, 81, 87, 96, 81, 73, 80, 85, 
    135, 173, 147, 46, 50, 49, 85, 99, 95, 93, 94, 84, 78, 88, 84, 
    138, 167, 150, 37, 47, 70, 91, 100, 92, 96, 90, 87, 85, 89, 87, 
    
    -- channel=9
    25, 36, 7, 26, 16, 0, 15, 28, 37, 39, 54, 43, 39, 83, 76, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 20, 71, 42, 42, 93, 100, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 14, 24, 41, 94, 130, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 21, 23, 66, 100, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 6, 23, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 
    
    
    others => 0);
end gold_package;
