-- https://docs.xilinx.com/r/en-US/ug953-vivado-7series-libraries/BRAM_SINGLE_MACRO

library UNISIM;
use UNISIM.vcomponents.all;
library UNIMACRO;
use unimacro.Vcomponents.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_signed.all;
use IEEE.std_logic_arith.all;

-- BRAM_SINGLE_MACRO: Single Port RAM
--                    7 Series
-- Xilinx HDL Language Template, version 2021.2

-- Note -  This Unimacro model assumes the port directions to be "downto".
--         Simulation of this model with "to" in the port directions could lead to erroneous results.

---------------------------------------------------------------------
--  READ_WIDTH | BRAM_SIZE | READ Depth  | ADDR Width |            --
-- WRITE_WIDTH |           | WRITE Depth |            |  WE Width  --
-- ============|===========|=============|============|============--
--    37-72    |  "36Kb"   |      512    |    9-bit   |    8-bit   --
--    19-36    |  "36Kb"   |     1024    |   10-bit   |    4-bit   --
--    19-36    |  "18Kb"   |      512    |    9-bit   |    4-bit   --
--    10-18    |  "36Kb"   |     2048    |   11-bit   |    2-bit   --
--    10-18    |  "18Kb"   |     1024    |   10-bit   |    2-bit   --
--     5-9     |  "36Kb"   |     4096    |   12-bit   |    1-bit   --
--     5-9     |  "18Kb"   |     2048    |   11-bit   |    1-bit   --
--     3-4     |  "36Kb"   |     8192    |   13-bit   |    1-bit   --
--     3-4     |  "18Kb"   |     4096    |   12-bit   |    1-bit   --
--       2     |  "36Kb"   |    16384    |   14-bit   |    1-bit   --
--       2     |  "18Kb"   |     8192    |   13-bit   |    1-bit   --
--       1     |  "36Kb"   |    32768    |   15-bit   |    1-bit   --
--       1     |  "18Kb"   |    16384    |   14-bit   |    1-bit   --
---------------------------------------------------------------------

entity bram_single is
    generic (
        -- replace ADDR_WIDHT, INPUT_SIZE and ADDRESS_SIZE generics with constants using python
        ADDR_WIDHT      : integer := 10;
        INPUT_SIZE      : integer := 8;
        ADDRESS_SIZE    : integer := 12;

        DEVICE     : string := "7SERIES";
        BRAM_NAME  : string := "default"
        );

    port (
        RST  : in std_logic;
        CLK  : in std_logic;
        EN   : in std_logic;
        WE   : in std_logic;
        DI   : in std_logic_vector(INPUT_SIZE-1 downto 0);
        ADDR : in std_logic_vector(ADDR_WIDHT-1 downto 0);
        DO   : out std_logic_vector(INPUT_SIZE-1 downto 0)
    );
 end bram_single;

  architecture a1 of bram_single is
    signal bram_wr_en    : std_logic_vector(4-1 downto 0);
    signal bram_addr     : std_logic_vector(10-1 downto 0);

    begin
    bram_wr_en <= (others => '1') when WE = '1' else (others => '0');
    bram_addr <= ADDR(10-1 downto 0);
          

    MEM_IWGHT_LAYER0_ENTITY0 : if BRAM_NAME = "iwght_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000018690000112a000008a40000001d00000894fffffa57000004fefffff05b",
            INIT_01 => X"00001da3ffffcfa000000a4b0000188d000013d2fffffebaffffdeecfffffcf0",
            INIT_02 => X"0000000400000000ffffffe5ffffffcafffffff70000000a000000220000001f",
            INIT_03 => X"00000018ffffffddffffffff00000038ffffffd30000002e0000002c00000003",
            INIT_04 => X"ffffffedffffffc3ffffffccffffffc900000018000000200000002100000035",
            INIT_05 => X"ffffffc0ffffffd30000001f0000001bffffffe60000000bffffffdaffffffc6",
            INIT_06 => X"0000000f000000250000001800000017fffffff500000010ffffffe2ffffffc6",
            INIT_07 => X"fffffff3000000320000000700000007ffffffd3fffffff6ffffffd8ffffffd8",
            INIT_08 => X"00000013ffffffcf0000000c00000006ffffffd8000000330000001d00000026",
            INIT_09 => X"ffffffeb0000000bfffffffbffffffff000000240000000500000020fffffff3",
            INIT_0A => X"ffffffdb0000000effffffecfffffff4ffffffdcffffffc1fffffffaffffffdf",
            INIT_0B => X"000000180000002d0000003700000006ffffffe1000000270000000900000032",
            INIT_0C => X"00000016ffffffee0000002d00000021ffffffe6000000020000001200000024",
            INIT_0D => X"ffffffd2fffffffc00000037ffffffc2fffffffbfffffff8ffffffc6ffffffe7",
            INIT_0E => X"0000001000000034000000000000001f00000040ffffffc20000001effffffe6",
            INIT_0F => X"fffffff6ffffffe6ffffffc6ffffffe5ffffffcc0000001e00000052fffffff5",
            INIT_10 => X"fffffffcffffffafffffffbefffffffa0000002b0000004dffffffeb0000002b",
            INIT_11 => X"ffffffc2ffffffe10000003900000044000000220000002bfffffffdffffffcd",
            INIT_12 => X"0000002cfffffff9fffffffa000000330000000b0000003900000001ffffffe1",
            INIT_13 => X"fffffffa0000002f000000450000003b0000002f0000001f0000002600000028",
            INIT_14 => X"fffffff800000021ffffffe400000018ffffffe6fffffff0ffffffef0000001b",
            INIT_15 => X"fffffff4ffffffc6ffffffcaffffffe500000004ffffffd2ffffffd6ffffffd5",
            INIT_16 => X"0000003300000030000000040000001c0000000000000019ffffffd6ffffffe9",
            INIT_17 => X"ffffffc1ffffffb300000005fffffffcffffffbe000000440000000dffffffd6",
            INIT_18 => X"ffffffbc0000001cffffffe400000009fffffff5ffffffd0fffffff000000022",
            INIT_19 => X"0000001100000040000000260000000e000000000000000f0000002500000010",
            INIT_1A => X"ffffffcdfffffff000000000000000340000001fffffffea0000002d00000033",
            INIT_1B => X"00000021ffffffd3ffffffbbffffffc4ffffffc900000009fffffff5fffffff6",
            INIT_1C => X"00000028ffffffc6fffffff200000000ffffffbaffffffc70000000a0000001c",
            INIT_1D => X"ffffffcbfffffff7000000330000003c00000034ffffffff0000002d00000015",
            INIT_1E => X"ffffffd100000017fffffff7fffffff8ffffffde000000030000002fffffffc7",
            INIT_1F => X"0000001c000000390000000bfffffffc0000000afffffff8ffffffc5ffffffc9",
            INIT_20 => X"fffffff8fffffffafffffffb0000000200000003fffffff9ffffffd5fffffff7",
            INIT_21 => X"0000001dffffffdf0000001e0000002bfffffff0ffffffc5ffffffc100000016",
            INIT_22 => X"000000280000003b00000020fffffff30000002d00000031000000170000001b",
            INIT_23 => X"0000003d00000014000000270000002cfffffff70000000600000029ffffffe9",
            INIT_24 => X"0000001dffffffc8ffffffd8fffffff1ffffffd2fffffff50000002500000025",
            INIT_25 => X"ffffffaeffffffbf0000002100000012ffffffe40000001e0000003100000010",
            INIT_26 => X"0000001000000035ffffffdaffffffdcfffffff3000000450000001dffffffe6",
            INIT_27 => X"ffffffd5ffffffe6fffffff7ffffffd00000001cffffffddffffffedffffffcb",
            INIT_28 => X"fffffff9ffffffe2ffffffe300000026fffffffdffffffd9ffffffe0ffffffec",
            INIT_29 => X"0000002cffffffea00000033000000160000002f0000001f0000000100000015",
            INIT_2A => X"ffffffe00000003effffffdbffffffc500000033fffffffbffffffe500000033",
            INIT_2B => X"0000002600000005ffffffd7fffffff800000028ffffffd70000001bfffffff9",
            INIT_2C => X"fffffffeffffffd8000000300000003afffffff30000004b0000000a00000003",
            INIT_2D => X"ffffffddfffffffaffffffebffffffd7ffffffff00000029ffffffc7fffffff9",
            INIT_2E => X"fffffffe0000004dfffffff900000034ffffffe4ffffffdfffffffd9ffffffc9",
            INIT_2F => X"000000030000003d0000001300000019ffffffecffffffbfffffffffffffffd6",
            INIT_30 => X"00000036ffffffff00000007ffffffe9ffffffbcfffffff2ffffffdb0000001b",
            INIT_31 => X"0000000a00000012000000240000000f00000038fffffffb0000003effffffe8",
            INIT_32 => X"0000002900000015fffffffa00000010ffffffe40000000a0000002d00000023",
            INIT_33 => X"0000001900000009ffffffe0ffffffdfffffffd1fffffffdfffffff7ffffffd1",
            INIT_34 => X"ffffffdd0000000dfffffff5ffffffeb0000001afffffff700000010ffffffda",
            INIT_35 => X"0000003100000002ffffffd2ffffffe400000013ffffffefffffffe100000018",
            INIT_36 => X"ffffffdbfffffff50000002b00000042fffffff0000000260000004600000014",
            INIT_37 => X"ffffffccfffffff200000023ffffffdaffffffe4fffffff7fffffff8ffffffcf",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IWGHT_LAYER0_ENTITY0;


    MEM_IFMAP_LAYER0_ENTITY0 : if BRAM_NAME = "ifmap_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000009f000000a20000009c000000a0000000a6000000a50000009f0000009e",
            INIT_01 => X"000000aa000000a9000000a6000000a1000000a0000000a10000009f0000009e",
            INIT_02 => X"0000009400000096000000950000009c000000a0000000a0000000a2000000a7",
            INIT_03 => X"000000740000007e000000890000008f0000008d0000008c0000008f00000095",
            INIT_04 => X"000000a2000000a4000000a0000000a2000000a60000009f0000009700000098",
            INIT_05 => X"000000ab000000ab000000aa000000a30000009f0000009b0000009c000000a3",
            INIT_06 => X"0000008d0000008c0000008b00000091000000970000009a000000a0000000a9",
            INIT_07 => X"000000770000007d000000880000008f0000008e000000910000009300000095",
            INIT_08 => X"000000a5000000a5000000a3000000a0000000a70000009e0000009700000097",
            INIT_09 => X"000000a9000000a7000000a6000000a10000009d0000009e000000a2000000a3",
            INIT_0A => X"0000007200000065000000620000006e00000079000000910000009f000000aa",
            INIT_0B => X"00000078000000820000008b0000008e0000008c0000008f0000008600000078",
            INIT_0C => X"000000a9000000a9000000a7000000a7000000ae000000a00000009b0000009b",
            INIT_0D => X"000000a4000000a20000009d000000b1000000bf000000a7000000a5000000a5",
            INIT_0E => X"0000004a000000500000005c000000620000006700000068000000950000009e",
            INIT_0F => X"0000007f000000880000008c0000008c00000084000000710000005300000056",
            INIT_10 => X"000000a6000000a9000000a3000000a9000000aa000000a10000009c0000009b",
            INIT_11 => X"0000008e0000009200000097000000c3000000f6000000ad000000a4000000a4",
            INIT_12 => X"0000005d000000610000006a0000007000000071000000550000004e0000006f",
            INIT_13 => X"00000081000000850000008a000000800000006900000055000000540000004a",
            INIT_14 => X"000000a7000000a7000000a5000000a100000093000000820000008500000094",
            INIT_15 => X"0000004200000061000000800000009d000000b4000000a3000000a5000000a3",
            INIT_16 => X"0000005e00000072000000770000007a00000076000000590000004200000045",
            INIT_17 => X"000000860000008a0000008c0000006c000000430000003a0000005b00000063",
            INIT_18 => X"000000aa000000a8000000aa00000099000000580000002f0000006d0000007f",
            INIT_19 => X"00000044000000640000007f0000008100000093000000a4000000a6000000a9",
            INIT_1A => X"0000006b000000690000007c000000920000008400000053000000480000004e",
            INIT_1B => X"000000860000008d000000840000004f0000002e0000003f0000005500000073",
            INIT_1C => X"000000a8000000a5000000a70000008f000000460000002a0000006300000083",
            INIT_1D => X"00000058000000740000009000000082000000780000008c000000a1000000ab",
            INIT_1E => X"0000006a0000006600000088000000a30000007c0000004d000000550000005b",
            INIT_1F => X"000000880000008a0000006b0000003900000031000000360000005500000064",
            INIT_20 => X"000000a6000000a3000000a1000000990000007c0000003600000067000000aa",
            INIT_21 => X"00000056000000790000009c0000009d0000007d00000071000000ae000000a5",
            INIT_22 => X"0000005700000071000000920000008a00000051000000500000005400000052",
            INIT_23 => X"00000089000000850000004a0000002800000038000000470000005600000053",
            INIT_24 => X"000000990000009c0000009e000000ae0000009a0000005e00000086000000b4",
            INIT_25 => X"0000005d0000007d00000094000000ae0000009c000000cf000000ed000000cf",
            INIT_26 => X"0000006a000000850000008f000000890000004c0000003b0000004a00000056",
            INIT_27 => X"000000840000005f00000028000000320000004b000000540000005700000056",
            INIT_28 => X"0000007a0000009f0000009b000000b1000000a50000008e0000006c000000b7",
            INIT_29 => X"000000780000007d0000009c000000b7000000a4000000dc000000ed000000d5",
            INIT_2A => X"0000006b0000009b0000009d000000af0000005b0000002d000000500000004e",
            INIT_2B => X"000000680000003b000000290000003b0000004e000000580000006700000057",
            INIT_2C => X"00000086000000ad000000a6000000bb000000aa0000008700000064000000bc",
            INIT_2D => X"0000007500000086000000bd000000b9000000aa000000c7000000c200000075",
            INIT_2E => X"0000005d00000092000000a0000000d20000007d000000260000005400000066",
            INIT_2F => X"0000004c0000003e000000370000004900000055000000680000005e00000053",
            INIT_30 => X"0000009f000000b2000000a6000000ae000000af0000007f0000005a000000bd",
            INIT_31 => X"0000007b000000a0000000d8000000ba00000089000000a8000000a800000061",
            INIT_32 => X"0000005b0000007b0000009b000000c200000096000000320000007300000078",
            INIT_33 => X"000000490000004f0000004900000054000000560000005f0000005400000054",
            INIT_34 => X"000000a7000000ad0000008800000077000000b9000000980000005d000000bd",
            INIT_35 => X"0000008d000000b4000000e2000000bd000000a7000000910000009300000067",
            INIT_36 => X"000000570000007200000095000000ba0000009a00000047000000750000007e",
            INIT_37 => X"0000005e000000610000005a0000006400000063000000500000004800000050",
            INIT_38 => X"000000a70000009c0000006300000069000000ba000000a80000006c000000c2",
            INIT_39 => X"0000009a00000091000000ac000000be000000c60000008a0000007300000064",
            INIT_3A => X"0000006e0000008200000089000000b300000098000000470000006700000092",
            INIT_3B => X"000000750000006100000064000000730000006d0000005f0000005b00000055",
            INIT_3C => X"0000009b0000008c0000004e00000082000000b8000000ac00000084000000c5",
            INIT_3D => X"000000830000008700000091000000f2000000e60000008f0000008200000073",
            INIT_3E => X"000000570000007000000098000000a8000000900000005f0000006c00000079",
            INIT_3F => X"0000008800000079000000670000007800000070000000690000005700000047",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000008a0000007e0000004e000000a8000000bf000000a800000092000000cb",
            INIT_41 => X"00000071000000710000008c000000a2000000ad0000009a000000600000008a",
            INIT_42 => X"0000006d00000087000000940000009c000000ab000000700000006900000065",
            INIT_43 => X"00000090000000970000007d0000006b000000650000005e0000004f0000004e",
            INIT_44 => X"0000009c000000600000005e000000b0000000b7000000a4000000a3000000d6",
            INIT_45 => X"0000007300000066000000740000007200000076000000810000006a00000094",
            INIT_46 => X"0000004b00000085000000800000004400000076000000900000006500000056",
            INIT_47 => X"0000008c000000960000008f0000007400000066000000470000003a0000003c",
            INIT_48 => X"0000008d000000560000007c000000b0000000ad000000a7000000b2000000d4",
            INIT_49 => X"00000093000000810000007c000000860000004d000000680000008700000099",
            INIT_4A => X"000000400000004b0000006b0000007500000084000000960000005c00000055",
            INIT_4B => X"000000970000009a000000a00000009b0000008500000056000000410000002c",
            INIT_4C => X"000000770000005600000090000000b1000000ae000000ab000000bb000000c7",
            INIT_4D => X"000000b8000000910000006c000000810000004600000090000000890000007a",
            INIT_4E => X"0000003400000033000000590000008600000089000000830000004900000074",
            INIT_4F => X"000000950000009e000000a4000000ab000000a3000000790000005a0000002f",
            INIT_50 => X"000000830000006300000098000000b5000000b1000000b3000000c3000000a5",
            INIT_51 => X"000000bf000000b20000007a0000005d000000500000005d00000067000000ab",
            INIT_52 => X"00000018000000260000002e0000003c00000057000000590000006400000096",
            INIT_53 => X"000000780000007f0000008000000090000000900000006c0000003c0000002e",
            INIT_54 => X"00000096000000530000008a000000b5000000b2000000b1000000c300000075",
            INIT_55 => X"000000c2000000be000000b0000000950000008600000085000000db000000f5",
            INIT_56 => X"0000003a0000003100000022000000230000003d0000006e0000007d000000a8",
            INIT_57 => X"000000370000003b000000450000004e00000048000000450000003a0000003d",
            INIT_58 => X"000000d30000006d0000008c000000b1000000b0000000ae000000af0000004f",
            INIT_59 => X"0000007a000000740000007c000000720000007c000000d0000000fc000000fd",
            INIT_5A => X"000000380000003300000032000000340000003c000000440000004400000068",
            INIT_5B => X"0000002a0000002b000000300000003b000000330000002b0000003300000038",
            INIT_5C => X"000000f6000000a5000000a5000000b2000000a8000000900000006000000029",
            INIT_5D => X"000000300000003100000031000000350000003c0000006e000000e3000000fd",
            INIT_5E => X"0000002b0000002e0000002e000000260000002a0000002e0000002a0000002d",
            INIT_5F => X"0000002d000000330000003500000037000000320000002e0000002e0000002a",
            INIT_60 => X"000000fe000000c200000084000000a6000000830000003b0000001d0000001d",
            INIT_61 => X"00000032000000310000003300000032000000320000003d0000008d000000f1",
            INIT_62 => X"0000002a00000026000000270000002300000022000000270000002a0000002f",
            INIT_63 => X"000000330000002e00000032000000380000003b0000003e000000380000002d",
            INIT_64 => X"00000100000000d7000000800000008000000049000000220000001e00000030",
            INIT_65 => X"0000002d0000002e0000003400000034000000320000003600000042000000bb",
            INIT_66 => X"0000002e0000002b00000028000000280000002700000024000000290000002b",
            INIT_67 => X"000000530000004600000032000000360000003b000000400000003e0000003b",
            INIT_68 => X"000000f0000000e00000008000000042000000290000001f0000002300000034",
            INIT_69 => X"0000002f0000002c0000002c0000003600000038000000310000003a0000007c",
            INIT_6A => X"0000003a000000360000002d0000002c0000002c0000002b0000002b0000002e",
            INIT_6B => X"0000004c000000550000004900000033000000240000002b0000002e00000036",
            INIT_6C => X"000000d3000000ca0000004e0000002c000000230000001d0000002300000032",
            INIT_6D => X"0000002d00000028000000300000003a00000030000000360000004100000061",
            INIT_6E => X"000000300000002700000027000000330000002e0000002f000000300000002f",
            INIT_6F => X"000000330000002e0000004300000043000000280000001c000000270000002f",
            INIT_70 => X"000000aa000000680000002e0000002900000021000000200000002300000032",
            INIT_71 => X"0000002d000000360000003a0000003d00000035000000340000003600000040",
            INIT_72 => X"00000027000000280000002a0000002e000000310000002e000000290000002a",
            INIT_73 => X"000000330000000f0000001f0000002f0000003f0000002c0000002800000025",
            INIT_74 => X"000000470000002a0000002b00000025000000260000001f0000002a00000044",
            INIT_75 => X"000000350000003a0000003800000031000000260000001b0000001f00000031",
            INIT_76 => X"00000021000000270000002d0000003200000035000000390000003c00000038",
            INIT_77 => X"000000280000000d0000002600000038000000490000004f0000003e0000002a",
            INIT_78 => X"000000280000002c0000002a000000270000002b00000023000000310000003d",
            INIT_79 => X"0000002f000000240000001d0000001b0000001e000000170000001b0000002a",
            INIT_7A => X"0000002b0000002b00000031000000450000004b000000420000003e00000038",
            INIT_7B => X"000000140000001d0000001a0000003c0000005d0000006d000000550000003c",
            INIT_7C => X"000000260000002800000028000000280000002b0000002d0000003800000036",
            INIT_7D => X"00000012000000130000001d000000190000001d000000160000001a00000024",
            INIT_7E => X"0000002d0000003400000035000000420000004a0000003d0000002f00000020",
            INIT_7F => X"0000001500000022000000180000003000000059000000690000005900000043",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY0;


    MEM_IFMAP_LAYER0_ENTITY1 : if BRAM_NAME = "ifmap_layer0_entity1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"00000071000000730000006d0000007000000076000000740000006f00000070",
            INIT_01 => X"0000007700000075000000750000006f0000006f00000074000000710000006f",
            INIT_02 => X"0000006a0000006b0000006b0000006d000000700000006f0000007100000075",
            INIT_03 => X"000000550000005b0000005f000000610000006100000062000000650000006b",
            INIT_04 => X"0000007200000075000000710000007000000074000000720000006e00000070",
            INIT_05 => X"000000730000007500000077000000710000006e0000006f0000006e00000074",
            INIT_06 => X"0000006400000066000000680000006e00000073000000700000006f00000073",
            INIT_07 => X"000000580000005b0000005f0000006200000061000000660000006600000069",
            INIT_08 => X"0000007500000075000000730000006a0000006f0000006f0000006d0000006e",
            INIT_09 => X"0000007100000072000000730000006f0000006d000000720000007300000073",
            INIT_0A => X"000000550000004d0000004e0000005a000000600000006f0000007200000074",
            INIT_0B => X"000000590000005f000000620000006300000063000000670000006000000056",
            INIT_0C => X"0000007700000078000000750000006e000000700000006d0000006e0000006b",
            INIT_0D => X"00000072000000730000006f00000082000000920000007b0000007500000073",
            INIT_0E => X"0000003f0000004b0000005a0000005a00000057000000500000006f00000070",
            INIT_0F => X"0000005e00000063000000650000006600000062000000550000003e00000046",
            INIT_10 => X"000000740000007800000071000000720000007200000073000000720000006b",
            INIT_11 => X"0000006c0000006f000000720000009c000000d6000000800000007400000071",
            INIT_12 => X"0000005e00000066000000720000006e00000067000000450000003500000050",
            INIT_13 => X"0000005d0000005e000000650000006000000053000000490000004e00000048",
            INIT_14 => X"000000730000007400000071000000730000007000000064000000680000006d",
            INIT_15 => X"000000320000004b000000660000007a0000008a00000076000000740000006f",
            INIT_16 => X"00000060000000740000007a000000790000007100000053000000380000003a",
            INIT_17 => X"0000005f0000006200000069000000540000003a0000003a0000005b00000064",
            INIT_18 => X"000000760000007300000076000000750000004a000000250000005f00000064",
            INIT_19 => X"00000043000000570000006c000000620000006b000000780000007400000075",
            INIT_1A => X"0000006600000063000000760000008e00000082000000540000004b00000053",
            INIT_1B => X"0000005d00000063000000620000003d0000002f00000047000000530000006f",
            INIT_1C => X"0000007400000072000000750000006f000000400000002b0000006000000073",
            INIT_1D => X"000000570000006a000000830000006e0000005e0000006d0000007100000077",
            INIT_1E => X"000000620000005d0000007c00000099000000760000004d000000580000005f",
            INIT_1F => X"0000006100000067000000530000002f000000350000003c000000510000005d",
            INIT_20 => X"0000007a00000075000000710000007c000000790000003a00000069000000a1",
            INIT_21 => X"000000500000006f0000008f0000008d00000069000000590000008700000079",
            INIT_22 => X"0000004f00000067000000870000007d000000470000004e0000005500000051",
            INIT_23 => X"000000670000006a0000003b000000230000003900000049000000520000004d",
            INIT_24 => X"000000760000007400000074000000950000009a000000640000008b000000b0",
            INIT_25 => X"000000550000006e000000830000009900000083000000b4000000d6000000b4",
            INIT_26 => X"000000620000007c000000850000007d00000044000000390000004a00000054",
            INIT_27 => X"000000670000004b0000001e000000310000004c000000550000005500000051",
            INIT_28 => X"0000005900000076000000700000009c000000a90000009700000074000000b7",
            INIT_29 => X"0000006f0000006c000000890000009f00000087000000bf000000e0000000c5",
            INIT_2A => X"000000640000009300000093000000a5000000550000002c000000500000004c",
            INIT_2B => X"000000510000002e000000240000003b0000004f000000580000006600000053",
            INIT_2C => X"0000005d0000007b00000078000000a7000000af000000900000006c000000bf",
            INIT_2D => X"0000006b00000077000000ab000000a10000008e000000ab000000b60000005f",
            INIT_2E => X"000000590000008b00000098000000c900000079000000260000005400000062",
            INIT_2F => X"0000003800000037000000350000004b00000057000000680000005d00000050",
            INIT_30 => X"0000006d0000007b0000007b0000009c000000b40000008600000060000000c2",
            INIT_31 => X"0000007100000095000000ca000000a600000072000000900000009a00000044",
            INIT_32 => X"000000580000007600000095000000bb00000093000000320000007200000072",
            INIT_33 => X"000000370000004a0000004900000057000000570000005f0000005400000053",
            INIT_34 => X"000000740000007c0000006a0000006e000000bc0000009a0000005f000000c0",
            INIT_35 => X"00000083000000ac000000d8000000ae000000950000007d0000008400000048",
            INIT_36 => X"000000550000006e00000090000000b500000098000000470000007200000075",
            INIT_37 => X"0000004900000059000000580000006500000064000000500000004900000050",
            INIT_38 => X"0000007a00000077000000590000006d000000ba000000a70000006b000000c4",
            INIT_39 => X"0000008f0000008c000000a5000000b4000000b90000007b0000006a0000004a",
            INIT_3A => X"0000006d0000008000000085000000af00000098000000470000006400000088",
            INIT_3B => X"0000005f0000005500000060000000740000006e000000600000005d00000056",
            INIT_3C => X"0000007d000000780000005300000089000000b2000000a700000081000000c5",
            INIT_3D => X"00000079000000820000008a000000ec000000dd00000083000000780000005e",
            INIT_3E => X"000000550000006c000000930000009f00000086000000580000006800000070",
            INIT_3F => X"0000006800000060000000560000006e0000006d000000680000005800000048",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000007e0000007d00000056000000aa000000b6000000a400000092000000cb",
            INIT_41 => X"0000006a0000006a0000008400000098000000a30000008f0000005000000079",
            INIT_42 => X"00000069000000820000008d0000008a0000008f0000005a0000006500000065",
            INIT_43 => X"000000680000006c00000058000000530000005b0000005d0000004f0000004c",
            INIT_44 => X"000000950000006000000066000000b6000000b8000000a7000000a6000000d7",
            INIT_45 => X"0000006e0000005b000000690000006600000069000000740000005d00000089",
            INIT_46 => X"000000450000007e00000078000000380000006000000080000000670000005b",
            INIT_47 => X"0000006e00000074000000700000005e0000005d000000460000003800000038",
            INIT_48 => X"0000008b0000005800000083000000b8000000b5000000af000000b8000000d3",
            INIT_49 => X"0000008f000000750000006f00000079000000400000005a0000008000000094",
            INIT_4A => X"0000003b00000044000000630000006d000000750000008b000000600000005c",
            INIT_4B => X"0000006f00000073000000780000007700000069000000450000003e00000029",
            INIT_4C => X"000000790000005a00000095000000b6000000b3000000b0000000bd000000c0",
            INIT_4D => X"000000b00000008600000061000000760000003b00000086000000880000007c",
            INIT_4E => X"000000330000003100000056000000810000007c000000770000004b00000076",
            INIT_4F => X"0000006b0000006f0000007100000079000000760000005b0000005a00000031",
            INIT_50 => X"00000087000000670000009d000000b5000000ad000000b2000000c10000009c",
            INIT_51 => X"000000b6000000ad000000760000005a0000004d0000005a00000069000000af",
            INIT_52 => X"000000210000002e000000340000003d0000004d0000004e0000006400000094",
            INIT_53 => X"00000069000000710000006d0000007b0000007d000000640000004700000039",
            INIT_54 => X"000000990000005700000090000000b3000000a9000000b2000000c800000078",
            INIT_55 => X"000000c0000000c4000000b60000009c0000008d0000008c000000de000000f7",
            INIT_56 => X"000000510000004600000036000000310000003e0000006d00000085000000ac",
            INIT_57 => X"0000005a0000005c000000600000006800000065000000630000005400000055",
            INIT_58 => X"000000d30000007000000092000000b1000000ac000000b7000000c500000069",
            INIT_59 => X"00000085000000850000008d000000840000008f000000e0000000fd000000fc",
            INIT_5A => X"0000005d00000055000000540000005400000052000000570000005d0000007c",
            INIT_5B => X"0000005f00000061000000610000006c00000068000000600000005b0000005e",
            INIT_5C => X"000000f5000000a6000000aa000000b6000000ae000000a80000008900000059",
            INIT_5D => X"000000480000004b0000004c000000500000005800000088000000e7000000fb",
            INIT_5E => X"00000057000000590000005a000000560000005200000051000000510000004f",
            INIT_5F => X"0000005a0000005f0000005e00000060000000600000005e0000005d00000059",
            INIT_60 => X"000000fa000000bd00000088000000b30000009900000066000000570000005b",
            INIT_61 => X"00000054000000530000005500000054000000540000005e0000009f000000f5",
            INIT_62 => X"000000590000005500000056000000530000004f000000520000005400000056",
            INIT_63 => X"000000670000005e00000063000000660000006500000067000000670000005c",
            INIT_64 => X"000000fd000000d500000088000000940000006a000000550000005e0000006f",
            INIT_65 => X"00000052000000530000005a0000005a000000580000005b0000005d000000c6",
            INIT_66 => X"0000005f0000005c000000590000005600000053000000500000005100000052",
            INIT_67 => X"000000890000007b000000690000006c0000006c0000006d0000006e0000006c",
            INIT_68 => X"000000f5000000e5000000910000005f00000053000000560000006300000072",
            INIT_69 => X"0000005300000052000000520000005c0000005e000000570000005c0000008f",
            INIT_6A => X"0000006e0000006a000000610000005a00000058000000560000005300000054",
            INIT_6B => X"0000007d0000008a000000820000006c0000005b0000005f0000006100000069",
            INIT_6C => X"000000e4000000db0000006a000000530000005600000059000000620000006e",
            INIT_6D => X"00000052000000500000005700000061000000570000005e000000680000007e",
            INIT_6E => X"000000660000005d0000005c0000006100000059000000590000005700000054",
            INIT_6F => X"00000060000000620000007e0000008100000065000000550000005d00000065",
            INIT_70 => X"000000c5000000850000005400000058000000580000005c000000610000006c",
            INIT_71 => X"000000530000006000000064000000670000005f0000005e0000006100000064",
            INIT_72 => X"0000005c0000005d0000005f0000005c0000005c00000058000000500000004f",
            INIT_73 => X"0000005d0000003c0000005a0000006e0000007d000000660000005d0000005a",
            INIT_74 => X"0000006b0000004f00000059000000570000005b00000058000000640000007c",
            INIT_75 => X"0000005c00000066000000640000005d00000052000000470000004d00000059",
            INIT_76 => X"00000053000000580000005e0000005f0000006100000063000000630000005e",
            INIT_77 => X"000000550000004000000061000000740000008300000084000000700000005b",
            INIT_78 => X"00000051000000580000005c0000005a0000005b000000550000006600000074",
            INIT_79 => X"000000560000005000000049000000470000004a000000430000004800000055",
            INIT_7A => X"00000058000000580000005f00000071000000770000006d000000650000005f",
            INIT_7B => X"00000040000000520000005200000073000000910000009c0000008200000069",
            INIT_7C => X"00000051000000570000005c000000590000005600000059000000690000006b",
            INIT_7D => X"0000003a0000003f00000049000000450000004900000042000000450000004f",
            INIT_7E => X"000000570000005f000000600000006f00000077000000680000005700000046",
            INIT_7F => X"00000043000000540000004d000000630000008700000092000000830000006d",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY1;


    MEM_IFMAP_LAYER0_ENTITY2 : if BRAM_NAME = "ifmap_layer0_entity2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000002d0000002f000000290000002e00000035000000330000002f00000031",
            INIT_01 => X"0000002c0000002d00000029000000310000003400000029000000290000002c",
            INIT_02 => X"0000002b0000002d0000002d0000002c0000002b000000270000002600000028",
            INIT_03 => X"00000021000000240000002400000026000000290000002b000000270000002c",
            INIT_04 => X"0000002d0000002f0000002b00000031000000380000002d0000002800000033",
            INIT_05 => X"000000210000002800000029000000340000003600000029000000260000002e",
            INIT_06 => X"000000300000003400000037000000350000003200000029000000210000001e",
            INIT_07 => X"00000022000000200000001f00000022000000260000002d0000002e00000032",
            INIT_08 => X"0000002d0000002d0000002c0000002a0000003000000024000000210000002f",
            INIT_09 => X"0000002300000025000000260000003300000039000000300000002b0000002b",
            INIT_0A => X"000000320000002f000000320000003400000031000000360000002f00000027",
            INIT_0B => X"0000002100000022000000220000002300000027000000330000003700000030",
            INIT_0C => X"00000030000000300000002e0000002b0000002c0000001f0000002000000028",
            INIT_0D => X"000000360000002f000000290000004b0000005f000000390000002d0000002c",
            INIT_0E => X"0000003200000042000000540000004c000000410000002f000000430000003a",
            INIT_0F => X"0000002400000027000000270000002b0000002e0000002d0000002700000034",
            INIT_10 => X"0000002c0000002f000000280000002b0000002f000000310000003000000029",
            INIT_11 => X"000000470000003c000000380000006b000000a40000003b0000002a00000029",
            INIT_12 => X"0000005d00000069000000760000006f00000062000000380000001f00000032",
            INIT_13 => X"00000024000000240000002e000000300000002d0000002f0000004600000043",
            INIT_14 => X"0000002900000029000000270000002c00000035000000390000004000000036",
            INIT_15 => X"0000001f0000002b0000003a0000004e000000550000002a0000002700000025",
            INIT_16 => X"00000060000000740000007a000000780000006e0000004c0000002d0000002b",
            INIT_17 => X"000000280000002c0000003a00000031000000250000002f0000005600000061",
            INIT_18 => X"0000002b000000280000002b000000300000001c000000110000005000000039",
            INIT_19 => X"00000039000000460000004b0000003b0000003400000027000000250000002a",
            INIT_1A => X"0000005e0000005a0000006c00000084000000790000004a0000004000000048",
            INIT_1B => X"00000027000000300000003a0000002400000027000000450000004d00000067",
            INIT_1C => X"00000027000000240000002a0000003800000029000000260000005c0000005a",
            INIT_1D => X"0000004f0000005d0000006b0000004d00000031000000330000003300000031",
            INIT_1E => X"0000005800000051000000700000008c0000006b000000450000005200000058",
            INIT_1F => X"00000027000000330000003200000020000000310000003a0000004a00000054",
            INIT_20 => X"00000032000000290000002b00000052000000710000003b0000006900000090",
            INIT_21 => X"0000004a0000006500000080000000790000004e0000003b0000005f00000042",
            INIT_22 => X"000000460000005d0000007b000000700000003d00000049000000520000004d",
            INIT_23 => X"0000002d0000003b000000230000001b00000035000000430000004c00000045",
            INIT_24 => X"0000003c0000002f000000330000007000000095000000690000008f000000a3",
            INIT_25 => X"0000004f0000006b0000007d0000009100000077000000a6000000c600000092",
            INIT_26 => X"00000059000000720000007a000000700000003a00000035000000470000004f",
            INIT_27 => X"000000390000002c0000000f0000002b000000470000004e0000004e0000004a",
            INIT_28 => X"0000002f00000033000000320000007a000000a80000009e0000007a000000af",
            INIT_29 => X"0000006800000068000000840000009b00000083000000bc000000e2000000b3",
            INIT_2A => X"0000005c0000008a000000890000009a0000004d000000280000004d00000045",
            INIT_2B => X"0000002e0000001f000000210000003b000000490000004f000000600000004d",
            INIT_2C => X"0000002c000000370000003b00000088000000b20000009900000074000000bd",
            INIT_2D => X"0000005f0000006a0000009f0000009700000085000000a4000000bc00000050",
            INIT_2E => X"00000052000000820000008e000000c000000071000000220000004f00000059",
            INIT_2F => X"0000001a00000030000000370000004e000000510000005e000000580000004b",
            INIT_30 => X"0000002f000000350000004400000085000000b90000009000000069000000c2",
            INIT_31 => X"0000006200000081000000b7000000940000005e0000007e000000980000002c",
            INIT_32 => X"000000530000006f0000008c000000b20000008c0000002f0000006d00000069",
            INIT_33 => X"000000180000004000000049000000590000005100000055000000500000004f",
            INIT_34 => X"000000320000003a0000004200000062000000c0000000a300000067000000c1",
            INIT_35 => X"000000750000009d000000c80000009b0000007f000000670000007800000027",
            INIT_36 => X"000000500000006800000088000000ae00000093000000440000006d0000006b",
            INIT_37 => X"000000220000004500000051000000630000005e00000048000000460000004c",
            INIT_38 => X"000000370000003e000000430000006d000000bc000000ac00000070000000c4",
            INIT_39 => X"000000860000008c0000009f000000a9000000a9000000670000005800000022",
            INIT_3A => X"000000690000007a0000007f000000aa00000095000000460000005f0000007d",
            INIT_3B => X"0000002f00000035000000500000006f000000680000005a0000005b00000053",
            INIT_3C => X"0000004d000000580000004d0000008e000000b5000000ae00000088000000c5",
            INIT_3D => X"000000700000008200000089000000e6000000d3000000740000005d00000034",
            INIT_3E => X"00000050000000650000008a00000092000000760000004b0000005f00000065",
            INIT_3F => X"0000003000000030000000360000005d00000063000000630000005700000044",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"000000710000007e0000005a000000ac000000bc000000b2000000a0000000cc",
            INIT_41 => X"0000005a00000058000000750000008d0000009b000000850000002500000052",
            INIT_42 => X"00000061000000760000007e0000006d000000680000003a000000570000005c",
            INIT_43 => X"0000002e000000370000002d00000037000000520000005e0000004d00000048",
            INIT_44 => X"000000910000006600000069000000ba000000c2000000b8000000b4000000d7",
            INIT_45 => X"000000620000004900000059000000590000005f000000690000003d0000006f",
            INIT_46 => X"0000003d00000073000000690000002000000040000000660000005f00000058",
            INIT_47 => X"000000360000004000000044000000400000004e000000410000003500000033",
            INIT_48 => X"0000008f0000006000000085000000bc000000c1000000bd000000c0000000cd",
            INIT_49 => X"0000008500000064000000600000006c00000037000000500000006f0000008d",
            INIT_4A => X"000000340000003a000000560000005c0000005d000000780000005d0000005d",
            INIT_4B => X"0000002e0000002d000000360000003e0000003b000000280000003c00000027",
            INIT_4C => X"000000840000006300000098000000b8000000b9000000b5000000bb000000b4",
            INIT_4D => X"000000a80000007b000000560000006c000000330000007e0000008700000082",
            INIT_4E => X"000000320000002c0000004e0000007600000069000000670000004900000076",
            INIT_4F => X"0000002e000000320000003400000040000000440000003c0000005d00000034",
            INIT_50 => X"000000920000006f000000a0000000b4000000ac000000af000000bb00000092",
            INIT_51 => X"000000b1000000ad000000740000005600000049000000570000006f000000b9",
            INIT_52 => X"000000290000003300000036000000390000003f000000420000006500000094",
            INIT_53 => X"0000003f000000450000003d0000004c000000520000004b0000005300000045",
            INIT_54 => X"0000009f0000005b00000093000000b3000000a8000000b0000000c80000007c",
            INIT_55 => X"000000c5000000d0000000c0000000a40000009300000090000000e1000000fa",
            INIT_56 => X"0000006600000057000000440000003a0000003e0000006d0000008f000000b5",
            INIT_57 => X"00000073000000700000007000000078000000770000007a0000006f0000006e",
            INIT_58 => X"000000d10000007100000096000000b6000000b1000000c0000000d500000085",
            INIT_59 => X"000000980000009c000000a2000000950000009d000000e8000000fc000000f7",
            INIT_5A => X"0000007d000000730000006e0000006f00000065000000680000007700000094",
            INIT_5B => X"0000008400000089000000840000008e0000008d000000870000008200000083",
            INIT_5C => X"000000ed000000a4000000ae000000c0000000bc000000bc000000a800000087",
            INIT_5D => X"000000650000006b00000069000000690000006f00000099000000e4000000f1",
            INIT_5E => X"000000800000007e0000007d0000007d00000074000000710000007800000073",
            INIT_5F => X"000000850000008b000000860000008700000089000000890000008b00000084",
            INIT_60 => X"000000f2000000b500000089000000bf000000b000000086000000820000008d",
            INIT_61 => X"00000074000000780000007900000077000000760000007f000000af000000f5",
            INIT_62 => X"000000820000007d0000007d0000007800000071000000730000007500000075",
            INIT_63 => X"000000950000008c00000090000000920000008e0000008e0000009100000086",
            INIT_64 => X"000000f9000000d10000008f000000a7000000880000007c0000008c000000a2",
            INIT_65 => X"00000073000000790000007f0000007f0000007d0000008000000076000000cd",
            INIT_66 => X"0000008a00000086000000830000007b00000075000000710000007000000071",
            INIT_67 => X"000000b6000000a7000000980000009a00000095000000930000009800000096",
            INIT_68 => X"000000f7000000ea000000a40000007e0000007a0000008200000093000000a5",
            INIT_69 => X"00000077000000770000007700000081000000830000007b0000007200000099",
            INIT_6A => X"0000009a000000960000008d000000830000007f0000007b0000007700000077",
            INIT_6B => X"000000a9000000b6000000b20000009e0000008a0000008c0000008d00000096",
            INIT_6C => X"000000ea000000e90000008a0000007e000000850000008a00000095000000a2",
            INIT_6D => X"00000077000000740000007b000000850000007c000000810000007e0000008c",
            INIT_6E => X"000000940000008b0000008a0000008c00000084000000820000007e0000007a",
            INIT_6F => X"0000008b0000008e000000b0000000b600000099000000850000008b00000093",
            INIT_70 => X"000000d30000009f0000007d0000008a0000008d0000008f00000093000000a1",
            INIT_71 => X"0000007800000083000000870000008b00000082000000800000007900000077",
            INIT_72 => X"000000880000008a0000008b0000008800000087000000820000007800000076",
            INIT_73 => X"00000088000000670000008c000000a4000000b2000000970000008a00000087",
            INIT_74 => X"0000008500000071000000840000008b000000920000008900000094000000b1",
            INIT_75 => X"0000008000000089000000870000008000000075000000690000006900000072",
            INIT_76 => X"0000007d0000008300000088000000890000008a0000008b0000008900000083",
            INIT_77 => X"0000007f0000006c00000092000000a8000000b5000000b30000009a00000085",
            INIT_78 => X"000000700000007d000000860000008b0000008f0000008400000094000000a8",
            INIT_79 => X"00000078000000730000006c0000006a0000006d000000660000006800000073",
            INIT_7A => X"0000007f0000007f00000086000000980000009c000000900000008700000080",
            INIT_7B => X"0000006b0000007e00000082000000a4000000be000000c5000000aa00000090",
            INIT_7C => X"000000730000007b0000008400000086000000860000008400000095000000a0",
            INIT_7D => X"00000059000000620000006c000000680000006c000000650000006900000072",
            INIT_7E => X"0000007b00000082000000830000009100000098000000890000007600000064",
            INIT_7F => X"0000006e000000810000007c00000091000000af000000b6000000a700000091",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_IFMAP_LAYER0_ENTITY2;


    MEM_GOLD_LAYER0_ENTITY0 : if BRAM_NAME = "gold_layer0_entity0" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"0000001d0000000f0000000d00000017000000140000000f0000001200000012",
            INIT_01 => X"00000016000000150000000c0000000600000001000000000000000a0000001d",
            INIT_02 => X"0000000000000003000000080000000400000013000000130000000f00000012",
            INIT_03 => X"0000000b000000000000000b0000000500000000000000000000000000000004",
            INIT_04 => X"00000000000000000000001e000000200000001b000000120000001b00000013",
            INIT_05 => X"0000000c00000000000000010000000100000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000110000000b00000019",
            INIT_07 => X"0000000300000003000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"0000000000000000000000040000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000001000000000000000000000000000000000000000000000000",
            INIT_0B => X"00000000000000000000001c0000000400000000000000000000000000000000",
            INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_0D => X"0000000000000000000000000000000200000000000000000000000000000000",
            INIT_0E => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_0F => X"000000000000000b000000000000000000000000000000000000000000000000",
            INIT_10 => X"000000000000000000000000000000000000000b000000000000000000000000",
            INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_12 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_15 => X"00000000000000000000000000000000000000000000000b0000000000000000",
            INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000020",
            INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"000000000000000000000000000000000000000000000000000000000000000b",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_2B => X"000000000000000d000000000000000000000000000000000000000000000000",
            INIT_2C => X"0000000000000000000000070000000400000000000000000000000000000000",
            INIT_2D => X"0000000000000000000000000000000000000006000000000000000000000000",
            INIT_2E => X"0000000000000000000000000000000000000000000000010000000000000000",
            INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_30 => X"0000000a0000003f0000000f0000001a0000000f000000000000000000000000",
            INIT_31 => X"0000002000000025000000380000003a00000032000000000000000000000000",
            INIT_32 => X"000000000000003a0000002c0000002000000027000000250000002900000022",
            INIT_33 => X"000000240000001f00000020000000200000001d0000001d0000001e00000000",
            INIT_34 => X"0000000e0000002f0000002f000000300000002100000028000000220000001e",
            INIT_35 => X"000000330000002f00000023000000220000001d00000019000000210000000f",
            INIT_36 => X"0000002a000000410000003100000033000000290000003a0000002800000034",
            INIT_37 => X"0000001a0000002d000000210000001c000000170000001f0000002a00000030",
            INIT_38 => X"000000000000000000000000000000000000000000000000000000290000001c",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3D => X"00000000000000000000000000000000000000060000000e0000001800000003",
            INIT_3E => X"000000000000000100000002000000000000000000000000000000000000000b",
            INIT_3F => X"0000001e0000000000000000000000000000000000000006000000000000001b",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000001d00000000000000030000000500000014000000110000000000000000",
            INIT_41 => X"00000000000000170000000f0000000300000000000000080000000000000010",
            INIT_42 => X"00000003000000440000000000000004000000060000000a0000001a00000000",
            INIT_43 => X"00000000000000000000000b0000001700000002000000000000000b00000000",
            INIT_44 => X"00000004000000000000003700000000000000000000000b0000001e0000000c",
            INIT_45 => X"000000060000000000000006000000140000002000000002000000110000000a",
            INIT_46 => X"000000110000000000000000000000200000000000000000000000000000002d",
            INIT_47 => X"00000000000000080000001100000004000000280000001d0000000000000008",
            INIT_48 => X"00000000000000060000000000000010000000000000000b0000000b00000000",
            INIT_49 => X"00000012000000090000000e0000002700000000000000240000001800000000",
            INIT_4A => X"00000000000000000000000c0000000000000000000000000000001500000012",
            INIT_4B => X"000000110000002d000000280000000d0000005800000000000000230000002b",
            INIT_4C => X"00000036000000000000000b0000001f000000220000001b0000000000000000",
            INIT_4D => X"0000001a000000210000001f0000000700000000000000450000001200000023",
            INIT_4E => X"000000380000002a0000002f0000002f0000002e00000028000000220000001e",
            INIT_4F => X"0000002a00000024000000240000002500000027000000000000002500000033",
            INIT_50 => X"000000520000002e0000002c0000003a0000002e0000002f000000360000002f",
            INIT_51 => X"0000002e0000002f0000002a0000002a000000260000002b0000001300000000",
            INIT_52 => X"000000190000002c000000330000002b00000028000000450000002a0000002f",
            INIT_53 => X"0000002e0000002d000000310000002e00000024000000230000002800000019",
            INIT_54 => X"00000000000000000000000000000000000000000000001f0000003a00000043",
            INIT_55 => X"00000000000000000000000a0000000200000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"00000000000000030000001c0000001f00000000000000170000000800000010",
            INIT_58 => X"0000002b00000000000000000000000000000000000000000000002a00000000",
            INIT_59 => X"00000000000000000000003f0000002d00000042000000000000000000000011",
            INIT_5A => X"0000002c00000028000000000000000e00000000000000000000000000000071",
            INIT_5B => X"0000006c000000000000002a0000003b000000260000005a0000000000000025",
            INIT_5C => X"0000003c000000480000005d0000002400000034000000000000002300000005",
            INIT_5D => X"0000003100000059000000000000003e0000001e000000520000002f00000000",
            INIT_5E => X"00000000000000600000003e000000610000002c000000000000000000000037",
            INIT_5F => X"0000001500000073000000480000002500000031000000120000005c00000073",
            INIT_60 => X"00000075000000000000006a0000004a0000005a000000000000000000000038",
            INIT_61 => X"0000003100000028000000650000004d000000370000000c0000001200000047",
            INIT_62 => X"000000500000004f0000000000000046000000380000008b0000000600000000",
            INIT_63 => X"0000002a0000000b000000840000004200000068000000130000002500000006",
            INIT_64 => X"000000040000005b0000001600000029000000000000002c0000002e00000013",
            INIT_65 => X"0000001800000064000000000000009f0000003a0000004a0000000000000000",
            INIT_66 => X"0000000000000000000000170000005a0000003b000000300000004d00000000",
            INIT_67 => X"000000200000004c0000009300000000000000940000003c0000000f0000000c",
            INIT_68 => X"0000003100000020000000230000001d0000001a000000410000008300000071",
            INIT_69 => X"0000003c0000003a00000073000000d8000000000000004e0000002b0000001d",
            INIT_6A => X"0000005f0000004f000000400000003e0000003c0000003d0000003800000047",
            INIT_6B => X"0000003e0000003f0000004900000042000000af000000820000000000000012",
            INIT_6C => X"000000450000006a0000003d0000004800000050000000400000003800000039",
            INIT_6D => X"000000410000003c000000420000004d000000390000005a000000cb00000000",
            INIT_6E => X"0000003e0000004b000000760000007b000000380000004e0000004d00000048",
            INIT_6F => X"0000005500000044000000380000004400000043000000350000004800000054",
            INIT_70 => X"00000008000000080000000000000000000000800000006f0000001a0000003a",
            INIT_71 => X"0000000000000000000000000000000400000000000000050000000300000006",
            INIT_72 => X"0000000a000000070000000c0000000a00000007000000050000000600000000",
            INIT_73 => X"0000000000000006000000240000000000000000000000000000001a00000049",
            INIT_74 => X"0000000000000007000000040000000400000000000000000000000400000000",
            INIT_75 => X"000000000000001700000007000000150000001a0000000d0000000000000000",
            INIT_76 => X"00000037000000000000000d0000000500000009000000250000002800000000",
            INIT_77 => X"000000000000000100000000000000000000000000000000000000050000001b",
            INIT_78 => X"0000000e0000000600000056000000800000000b000000130000005a00000026",
            INIT_79 => X"0000000000000000000000180000000f00000025000000250000000000000000",
            INIT_7A => X"0000001f0000001a0000002a0000000000000000000000000000000800000000",
            INIT_7B => X"000000070000000600000027000000090000000000000000000000000000003a",
            INIT_7C => X"00000011000000090000000a0000000000000021000000000000000400000000",
            INIT_7D => X"0000001c00000007000000150000001d00000017000000000000000b00000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000160000001900000010",
            INIT_7F => X"000000040000000b000000040000001000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY0;


    MEM_GOLD_LAYER0_ENTITY1 : if BRAM_NAME = "gold_layer0_entity1" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000000000000000000000000000040000001a00000000000000000000001c",
            INIT_01 => X"00000011000000040000000900000000000000000000002f0000000300000000",
            INIT_02 => X"0000001b0000000000000000000000000000000c0000004a0000000000000000",
            INIT_03 => X"000000850000009c00000046000000000000000000000000000000000000001f",
            INIT_04 => X"000000000000001b000000410000002000000000000000000000000000000028",
            INIT_05 => X"000000000000000000000000000000460000000f000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000002",
            INIT_08 => X"0000000000000011000000000000000000000012000000070000000400000000",
            INIT_09 => X"0000000000000000000000080000000000000000000000000000000000000000",
            INIT_0A => X"0000000000000000000000000000001300000000000000000000000000000000",
            INIT_0B => X"0000001300000014000000000000000000000000000000000000000000000000",
            INIT_0C => X"000000a2000000a30000009d0000000000000022000000280000000000000004",
            INIT_0D => X"0000007c00000094000000ad000000b7000000ac0000009d000000a4000000a5",
            INIT_0E => X"000000ac000000a8000000ad000000a20000009200000092000000840000007c",
            INIT_0F => X"0000003e0000002e0000003a0000007a000000a0000000a90000008c000000a0",
            INIT_10 => X"000000af000000b0000000ac0000006a000000890000008b0000006e0000004e",
            INIT_11 => X"000000270000000a0000001e000000070000002d00000048000000730000008e",
            INIT_12 => X"00000059000000a2000000aa000000a40000002b0000004d000000670000003a",
            INIT_13 => X"000000250000001b0000002d000000330000000c00000015000000270000004d",
            INIT_14 => X"00000043000000470000004e00000060000000940000001f000000170000003a",
            INIT_15 => X"0000002f0000001c000000170000003900000031000000000000001f0000002f",
            INIT_16 => X"00000031000000450000003b00000025000000990000008e0000001200000016",
            INIT_17 => X"0000000e0000001700000012000000100000002a0000003e000000000000002d",
            INIT_18 => X"0000002f0000002d0000003e000000320000002f0000009f000000620000002a",
            INIT_19 => X"0000000a0000001c000000260000000e00000010000000280000003200000000",
            INIT_1A => X"0000001e00000029000000270000002e0000002600000037000000620000002c",
            INIT_1B => X"0000002b00000000000000140000004100000022000000090000002d0000002f",
            INIT_1C => X"00000042000000540000000d000000300000003600000022000000550000000e",
            INIT_1D => X"00000000000000240000000500000010000000790000002d0000000f00000026",
            INIT_1E => X"000000060000001d000000340000002d00000028000000080000002000000035",
            INIT_1F => X"00000017000000000000002300000015000000000000008a0000006200000009",
            INIT_20 => X"000000000000000000000000000000000000000600000000000000000000001a",
            INIT_21 => X"000000000000003a000000060000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000003400000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_28 => X"0000002300000022000000000000000000000000000000000000000000000000",
            INIT_29 => X"000000170000001d0000002400000026000000270000001e0000002000000025",
            INIT_2A => X"0000002a0000002c00000023000000180000001e00000024000000260000001a",
            INIT_2B => X"000000000000001d0000000e0000001d0000000f00000020000000280000001f",
            INIT_2C => X"000000210000002800000039000000060000001c0000002b0000002000000009",
            INIT_2D => X"00000000000000000000002e0000002100000006000000000000001a00000027",
            INIT_2E => X"0000000f00000029000000210000004c000000000000002c0000002500000000",
            INIT_2F => X"0000000000000009000000000000004800000000000000000000000400000024",
            INIT_30 => X"0000000b00000009000000560000000200000026000000000000004a00000000",
            INIT_31 => X"0000000000000006000000000000000000000059000000000000000000000000",
            INIT_32 => X"00000000000000130000003e0000001a000000000000000a000000000000002b",
            INIT_33 => X"00000000000000000000001400000000000000000000008e0000000000000000",
            INIT_34 => X"0000000000000000000000360000003f00000000000000200000000000000000",
            INIT_35 => X"0000000000000000000000150000000a00000000000000000000006600000000",
            INIT_36 => X"0000000000000000000000000000004200000038000000000000000000000000",
            INIT_37 => X"0000000200000000000000080000000f0000001d000000000000000000000042",
            INIT_38 => X"0000000000000024000000000000000000000011000000040000002100000000",
            INIT_39 => X"00000000000000000000000000000023000000210000001e0000000000000025",
            INIT_3A => X"00000000000000050000000200000000000000270000000f000000000000002c",
            INIT_3B => X"0000007800000000000000040000002a0000001400000034000000300000000c",
            INIT_3C => X"0000000900000008000000000000000000000000000000220000000000000000",
            INIT_3D => X"0000000000000040000000000000001400000020000000000000000000000001",
            INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3F => X"0000000000000000000000000000004300000021000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_41 => X"000000000000000000000000000000000000005d000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000002b00000000000000000000000400000000000000000000000000000000",
            INIT_45 => X"000000370000003a00000030000000290000002f0000002c0000002d00000030",
            INIT_46 => X"000000350000002c000000310000002a0000002700000026000000250000002a",
            INIT_47 => X"0000000c0000003b000000290000001f000000000000002d0000002e00000030",
            INIT_48 => X"0000002e000000290000001c000000250000001f0000000e0000000000000000",
            INIT_49 => X"000000000000000000000000000000230000002d0000003b0000003200000035",
            INIT_4A => X"000000320000002300000000000000000000001a000000040000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000001900000025",
            INIT_4C => X"0000000000000018000000120000000000000000000000110000000000000006",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000300000003000000380000000b00000000000000000000000500000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000070000003a00000007000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000200000000000000000000000000000000",
            INIT_53 => X"000000000000000d000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000050000001a00000000000000000000000000000000",
            INIT_55 => X"000000000000000000000008000000000000000400000018000000030000000f",
            INIT_56 => X"0000000800000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000001f00000000000000000000000a00000011",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000b0000000c0000000c000000040000000800000008000000110000000a",
            INIT_62 => X"00000000000000060000000800000011000000230000002d000000210000000b",
            INIT_63 => X"00000042000000230000000500000000000000080000000c0000000a0000000a",
            INIT_64 => X"00000033000000350000000a000000170000000a000000000000000000000000",
            INIT_65 => X"0000000000000000000000090000001600000037000000050000000800000005",
            INIT_66 => X"0000000500000000000000000000000c0000000e000000000000000000000000",
            INIT_67 => X"000000040000001a000000000000000200000000000000000000000800000008",
            INIT_68 => X"0000000e0000000200000000000000010000000e000000000000000600000010",
            INIT_69 => X"0000000000000000000000000000000700000000000000090000000000000000",
            INIT_6A => X"0000003e0000000300000006000000000000000f000000000000000000000000",
            INIT_6B => X"0000000700000015000000140000000000000000000000000000000000000028",
            INIT_6C => X"0000000000000012000000180000001c00000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000001100000000000000110000000000000031",
            INIT_6E => X"0000003500000035000000020000000000000000000000000000000000000000",
            INIT_6F => X"000000000000000e000000050000000000000009000000000000000e00000021",
            INIT_70 => X"0000000000000000000000260000000000000000000000000000000100000000",
            INIT_71 => X"0000000c00000000000000000000000000000030000000260000000000000000",
            INIT_72 => X"0000000000000000000000000000000900000023000000000000000400000000",
            INIT_73 => X"000000000000000300000018000000000000000000000011000000360000004e",
            INIT_74 => X"0000000000000037000000510000001e00000000000000000000000000000007",
            INIT_75 => X"0000000c00000021000000350000000a00000005000000000000000000000000",
            INIT_76 => X"0000000000000000000000030000000500000004000000280000005600000000",
            INIT_77 => X"0000001800000000000000160000000000000000000000000000000000000000",
            INIT_78 => X"000000000000000000000000000000000000000000000000000000000000003f",
            INIT_79 => X"0000000b0000004f000000180000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000300000000000000220000000000000000000000000000001400000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000012",
            INIT_7D => X"0000000800000015000000090000000e0000000a000000130000000d00000000",
            INIT_7E => X"0000000200000006000000130000001b000000220000001c0000000c00000006",
            INIT_7F => X"0000001a0000000f000000360000000f0000000d000000090000000b00000008",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY1;


    MEM_GOLD_LAYER0_ENTITY2 : if BRAM_NAME = "gold_layer0_entity2" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000260000000a0000001a000000210000002400000035000000340000001f",
            INIT_01 => X"00000020000000280000003300000051000000080000000a0000000b00000024",
            INIT_02 => X"00000014000000330000001a000000190000002b0000004b0000005e00000053",
            INIT_03 => X"0000005b000000360000002f000000450000002e00000019000000120000000e",
            INIT_04 => X"000000150000005e000000710000001b000000150000003b000000420000005d",
            INIT_05 => X"000000670000003b000000330000003b00000064000000440000007e00000035",
            INIT_06 => X"00000013000000280000009e0000007f00000001000000250000003900000038",
            INIT_07 => X"000000500000007f0000005b0000002e0000004b0000007d0000007e000000bd",
            INIT_08 => X"0000005a0000001700000043000000940000007a000000150000003c00000047",
            INIT_09 => X"0000003b0000004600000081000000780000004e00000065000000a800000075",
            INIT_0A => X"000000a5000000390000003900000040000000a50000008e000000330000004c",
            INIT_0B => X"0000004b000000480000004c000000780000005f000000500000006a00000085",
            INIT_0C => X"0000005900000066000000380000007300000066000000b8000000b000000026",
            INIT_0D => X"0000000e0000002b0000002c000000410000006500000033000000510000004e",
            INIT_0E => X"000000790000005f000000330000006f0000007500000086000000b3000000c0",
            INIT_0F => X"000000c700000027000000270000002f00000025000000400000005a00000042",
            INIT_10 => X"00000079000000b900000091000000650000009e000000a20000008b000000ab",
            INIT_11 => X"000000cb000000c100000068000000710000005a00000047000000400000003c",
            INIT_12 => X"0000006f0000007c000000850000008a000000a5000000e7000000c90000009d",
            INIT_13 => X"000000b1000000a10000008c0000008e0000008a000000880000008000000078",
            INIT_14 => X"00000084000000760000007100000070000000750000007a000000af000000e5",
            INIT_15 => X"000000ef000000a6000000850000009d000000a30000009a000000950000008c",
            INIT_16 => X"0000009b0000008c000000820000007700000073000000790000008000000088",
            INIT_17 => X"00000074000000a70000007f0000008f00000097000000ab000000a300000093",
            INIT_18 => X"0000009a0000008500000086000000880000007c0000007e000000890000007f",
            INIT_19 => X"0000000000000000000000000000000000000000000000000000008d000000af",
            INIT_1A => X"00000000000000000000000b0000001c00000013000000000000000000000000",
            INIT_1B => X"0000000b00000000000000000000000000000000000000000000000000000000",
            INIT_1C => X"00000000000000000000001e0000001400000000000000000000003300000014",
            INIT_1D => X"000000280000001c0000003e000000000000000000000000000000000000003f",
            INIT_1E => X"00000019000000000000001e0000000700000000000000000000000000000000",
            INIT_1F => X"000000000000000000000000000000000000000c000000000000000000000000",
            INIT_20 => X"0000000000000000000000000000000e000000060000001a0000000000000000",
            INIT_21 => X"000000000000001d000000040000000f00000000000000000000000000000009",
            INIT_22 => X"00000002000000000000002f0000002500000000000000000000000800000000",
            INIT_23 => X"000000260000000000000006000000000000000000000000000000030000004f",
            INIT_24 => X"0000000d0000000d00000018000000000000000000000000000000000000001c",
            INIT_25 => X"0000000800000018000000000000000900000000000000050000000000000000",
            INIT_26 => X"0000000000000000000000070000000000000002000000000000000000000000",
            INIT_27 => X"000000000000001c0000000000000000000000000000001e0000003d00000000",
            INIT_28 => X"0000003200000022000000000000002e00000000000000000000000000000010",
            INIT_29 => X"000000000000000d0000003a0000002600000036000000000000000000000003",
            INIT_2A => X"000000000000001500000012000000000000000a000000000000000000000000",
            INIT_2B => X"00000008000000000000000000000001000000310000001f0000002e00000000",
            INIT_2C => X"0000001900000000000000000000000000000000000000220000000000000000",
            INIT_2D => X"0000004100000021000000160000000000000000000000000000000d0000000f",
            INIT_2E => X"0000000c000000370000003f00000052000000a2000000000000000000000000",
            INIT_2F => X"000000360000000d000000000000000000000000000000020000000000000006",
            INIT_30 => X"0000000000000000000000000000000200000000000000560000004100000000",
            INIT_31 => X"0000002500000000000000020000000000000000000000030000000000000000",
            INIT_32 => X"000000070000000000000000000000010000000000000000000000060000003e",
            INIT_33 => X"0000003600000018000000000000000c0000004200000000000000000000000a",
            INIT_34 => X"0000000000000005000000000000000000000000000000090000001300000024",
            INIT_35 => X"0000000000000000000000000000000000000000000000040000000000000000",
            INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_3A => X"00000000000000000000000000000000000000000000001f0000000400000000",
            INIT_3B => X"0000000000000000000000000000000000000000000000000000000b00000000",
            INIT_3C => X"0000000000000001000000020000000000000007000000000000002d00000005",
            INIT_3D => X"0000000200000000000000000000000000000000000000000000000000000002",
            INIT_3E => X"000000060000000100000010000000000000000300000000000000000000003b",
            INIT_3F => X"0000005d000000000000000000000000000000000000002c0000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"00000000000000000000000000000000000000000000000e0000000000000000",
            INIT_41 => X"00000000000000520000000000000000000000000000000f0000001c00000000",
            INIT_42 => X"0000000000000000000000000000000400000000000000130000001200000000",
            INIT_43 => X"00000000000000000000002d000000000000000500000000000000170000000c",
            INIT_44 => X"000000000000001100000000000000160000000000000000000000030000001d",
            INIT_45 => X"0000001b00000000000000110000000000000008000000000000000000000012",
            INIT_46 => X"00000003000000000000003b0000000000000019000000090000000000000000",
            INIT_47 => X"0000000000000012000000120000000000000000000000050000000000000010",
            INIT_48 => X"0000002d000000000000000000000058000000000000000d0000003300000000",
            INIT_49 => X"0000001d0000002c0000003e0000003300000028000000020000000000000004",
            INIT_4A => X"0000004e0000004e0000002e000000000000003b000000000000003600000070",
            INIT_4B => X"0000005a000000530000005a00000058000000560000004f0000004900000044",
            INIT_4C => X"0000004c0000004a00000048000000490000000000000008000000480000006f",
            INIT_4D => X"000000600000005a0000005e0000005d000000570000005b0000005b00000054",
            INIT_4E => X"00000057000000530000004d000000450000005000000031000000000000008a",
            INIT_4F => X"0000006700000067000000500000005e00000074000000610000006400000061",
            INIT_50 => X"00000052000000520000005200000049000000550000005f0000004900000041",
            INIT_51 => X"0000002e000000330000002e0000002f00000045000000530000006b0000005e",
            INIT_52 => X"000000270000001c000000230000002b0000002f000000310000002f0000002f",
            INIT_53 => X"000000340000002d000000350000003200000032000000240000002700000026",
            INIT_54 => X"0000002400000015000000130000002100000004000000250000001300000055",
            INIT_55 => X"0000002c000000380000002e000000340000003b0000001a000000280000002d",
            INIT_56 => X"00000027000000040000000b0000000a0000004f0000001a0000000000000000",
            INIT_57 => X"0000001a0000002300000025000000360000002c000000790000000000000039",
            INIT_58 => X"000000530000000e000000000000001200000000000000530000001800000008",
            INIT_59 => X"00000000000000000000001a0000002c000000490000000a0000006300000000",
            INIT_5A => X"0000000000000039000000000000001e000000000000000b0000005f00000008",
            INIT_5B => X"00000000000000000000000000000000000000490000002e0000000000000038",
            INIT_5C => X"00000015000000000000000d00000004000000230000000000000000000000bf",
            INIT_5D => X"000000a400000000000000000000000a0000005000000061000000000000000c",
            INIT_5E => X"0000000100000000000000000000000d000000270000001e0000000000000000",
            INIT_5F => X"000000000000007c000000000000000800000000000000680000004500000000",
            INIT_60 => X"0000003c00000000000000170000000000000012000000220000002a00000000",
            INIT_61 => X"000000000000002200000006000000310000001c000000000000000300000011",
            INIT_62 => X"000000000000004a00000000000000180000000a000000440000003a00000026",
            INIT_63 => X"0000004800000005000000000000000a000000170000000e0000002a00000019",
            INIT_64 => X"0000000b00000000000000a30000000000000011000000510000001c00000056",
            INIT_65 => X"0000001e0000002d000000280000001400000000000000000000000000000056",
            INIT_66 => X"0000000000000000000000000000009800000000000000280000004000000000",
            INIT_67 => X"00000000000000110000000e0000001000000010000000090000000000000000",
            INIT_68 => X"0000000a0000000500000009000000000000001f000000480000004100000003",
            INIT_69 => X"0000000000000017000000080000001000000017000000140000001000000008",
            INIT_6A => X"0000000d00000009000000000000001100000000000000000000007400000010",
            INIT_6B => X"0000000d00000000000000000000002600000000000000090000000d00000010",
            INIT_6C => X"0000001000000018000000090000000c00000016000000000000000000000019",
            INIT_6D => X"0000000000000000000000000000000000000003000000310000000b00000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000001000000000000000000000000000000000000000400000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000012000000040000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000005",
            INIT_75 => X"0000000000000008000000380000000000000000000000270000000100000000",
            INIT_76 => X"0000000000000004000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"000000000000000f000000000000000000000000000000000000001400000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000012000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY2;


    MEM_GOLD_LAYER0_ENTITY3 : if BRAM_NAME = "gold_layer0_entity3" generate
        BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
        generic map (
            BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
            DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
            DO_REG => 0,                     -- Optional output register (0 or 1)
            INIT => X"000000000000000000",   -- Initial values on output port
            INIT_FILE => "NONE",
            WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
            SRVAL => X"000000000000000000",  -- Set/Reset value for port output
            WRITE_MODE => "WRITE_FIRST",     -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
            -- The following INIT_xx declarations specify the initial contents of the RAM
            INIT_00 => X"000000300000001e000000000000000000000000000000000000000000000011",
            INIT_01 => X"00000001000000240000001c000000000000000000000000000000000000003e",
            INIT_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_05 => X"0000000200000000000000000000000000000000000000000000000000000000",
            INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_09 => X"000000360000002f000000000000000000000013000000000000000000000000",
            INIT_0A => X"0000002b000000360000003b0000003900000030000000350000003500000033",
            INIT_0B => X"0000003600000038000000300000002700000028000000250000002000000020",
            INIT_0C => X"000000020000000200000023000000390000003b000000420000003300000039",
            INIT_0D => X"0000003900000036000000130000003000000027000000110000000600000006",
            INIT_0E => X"00000000000000040000000000000000000000000000001e0000003d00000037",
            INIT_0F => X"0000004000000037000000320000000000000015000000170000000000000001",
            INIT_10 => X"0000000000000000000000170000000000000000000000000000001e00000012",
            INIT_11 => X"0000003300000044000000100000003400000012000000000000000000000000",
            INIT_12 => X"0000000000000000000000090000001000000000000000000000000600000025",
            INIT_13 => X"0000002b0000000d0000000b00000038000000310000000f0000000000000000",
            INIT_14 => X"000000000000000000000000000000000000002a000000000000000b00000008",
            INIT_15 => X"000000170000002e000000110000000e0000003d000000070000002c00000000",
            INIT_16 => X"0000000400000000000000000000000000000000000000130000000300000008",
            INIT_17 => X"000000000000000a0000002e0000002200000000000000250000000000000019",
            INIT_18 => X"0000001100000015000000000000000200000000000000000000000f00000013",
            INIT_19 => X"0000002c000000000000000c00000000000000000000001c0000000000000009",
            INIT_1A => X"000000140000000e000000160000002100000000000000000000000000000000",
            INIT_1B => X"0000000000000005000000060000001f00000000000000000000000300000000",
            INIT_1C => X"00000000000000150000001400000005000000280000001e0000000000000000",
            INIT_1D => X"000000000000000000000000000000000000001700000011000000060000002c",
            INIT_1E => X"0000003c00000032000000000000000000000000000000000000000000000000",
            INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_20 => X"00000000000000000000004f0000000000000000000000000000000000000000",
            INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_22 => X"0000000000000000000000000000002800000000000000000000000000000000",
            INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_25 => X"0000002700000000000000000000000000000000000000000000000000000000",
            INIT_26 => X"0000002f0000002b00000028000000200000002c000000290000002300000022",
            INIT_27 => X"00000024000000280000002e000000290000001e0000001d0000002900000032",
            INIT_28 => X"000000050000002e00000030000000430000000e000000210000002c00000024",
            INIT_29 => X"00000028000000020000003f0000002c00000015000000190000002900000021",
            INIT_2A => X"0000001c00000000000000100000002400000028000000200000002a00000029",
            INIT_2B => X"000000240000002e000000000000005c0000000b0000001a000000320000000c",
            INIT_2C => X"0000001800000023000000000000001900000025000000270000000c00000038",
            INIT_2D => X"000000130000000000000041000000050000002c00000000000000260000001a",
            INIT_2E => X"0000001200000038000000140000000000000025000000240000002a00000027",
            INIT_2F => X"00000000000000000000002f0000003700000000000000240000001a0000002b",
            INIT_30 => X"0000001d000000070000002a0000003400000000000000430000002500000016",
            INIT_31 => X"000000150000000000000000000000460000000e000000240000001100000020",
            INIT_32 => X"00000025000000000000000d000000280000002b00000000000000390000001c",
            INIT_33 => X"0000000b0000003500000000000000020000003400000029000000060000000b",
            INIT_34 => X"0000000d0000000d00000011000000000000002c000000110000000000000018",
            INIT_35 => X"000000000000001b0000000e0000000000000034000000000000003f00000000",
            INIT_36 => X"00000000000000000000001a00000000000000000000002b000000050000003f",
            INIT_37 => X"0000000f0000002c0000001d00000000000000140000002a0000000000000039",
            INIT_38 => X"0000003800000000000000000000002f00000010000000000000000f0000002f",
            INIT_39 => X"0000000f0000002b000000270000000500000000000000320000002900000000",
            INIT_3A => X"0000000000000000000000000000000000000021000000110000000800000008",
            INIT_3B => X"0000000000000003000000070000000000000000000000000000000500000052",
            INIT_3C => X"0000002e00000022000000000000000000000014000000030000000000000000",
            INIT_3D => X"0000000200000000000000000000000100000005000000020000000600000000",
            INIT_3E => X"000000000000000d000000220000000000000000000000090000000000000000",
            INIT_3F => X"0000000000000000000000000000000100000000000000000000000600000009",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INIT_40 => X"0000000000000000000000140000000400000000000000000000001300000015",
            INIT_41 => X"0000001a0000001200000000000000000000000c000000000000000000000000",
            INIT_42 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_43 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_44 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_45 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_46 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_47 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_48 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_49 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_4F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_50 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_51 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_52 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_53 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_54 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_55 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_56 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_57 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_58 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_59 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_5F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_60 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_61 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_62 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_63 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_64 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_65 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_66 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_67 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_68 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_69 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_6F => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_70 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_71 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_72 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_73 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_74 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_75 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_76 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_77 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_78 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_79 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INIT_7F => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INITP_xx are for the parity bits
            INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000",

            -- The next set of INIT_xx are valid when configured as 36Kb
            INITP_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
            INITP_0F => X"0000000000000000000000000000000000000000000000000000000000000000"
        )
        port map (
            DO => DO,      -- Output data, width defined by READ_WIDTH parameter
            ADDR => bram_addr,  -- Input address, width defined by read/write port depth
            CLK => CLK,    -- 1-bit input clock
            DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
            EN => EN,      -- 1-bit input RAM enable
            REGCE => '1', -- 1-bit input output register enable
            RST => RST,    -- 1-bit input reset
            WE => bram_wr_en       -- Input write enable, width defined by write port depth
        );
    -- End of BRAM_SINGLE_MACRO_inst instantiation
    end generate MEM_GOLD_LAYER0_ENTITY3;

MEM_EMPTY_36Kb : if BRAM_NAME = "default" generate
    BRAM_SINGLE_MACRO_inst : BRAM_SINGLE_MACRO
    generic map (
        BRAM_SIZE => "36Kb",             -- Target BRAM, "18Kb" or "36Kb"
        DEVICE => DEVICE,                -- Target Device: "VIRTEX5", "7SERIES", "VIRTEX6, "SPARTAN6"
        DO_REG => 0,                     -- Optional output register (0 or 1)
        INIT => X"000000000000000000",   -- Initial values on output port
        INIT_FILE => "NONE",
        WRITE_WIDTH => INPUT_SIZE, -- 0, -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        READ_WIDTH => INPUT_SIZE, -- 0,  -- Valid values are 1-72 (37-72 only valid when BRAM_SIZE="36Kb")
        SRVAL => X"000000000000000000",  -- Set/Reset value for port output
        WRITE_MODE => "WRITE_FIRST"      -- "WRITE_FIRST", "READ_FIRST" or "NO_CHANGE"
    )
    port map (
        DO => DO,      -- Output data, width defined by READ_WIDTH parameter
        ADDR => bram_addr,  -- Input address, width defined by read/write port depth
        CLK => CLK,    -- 1-bit input clock
        DI => DI,      -- Input data port, width defined by WRITE_WIDTH parameter
        EN => EN,      -- 1-bit input RAM enable
        REGCE => '1', -- 1-bit input output register enable
        RST => RST,    -- 1-bit input reset
        WE => bram_wr_en       -- Input write enable, width defined by write port depth
    );
-- End of BRAM_SINGLE_MACRO_inst instantiation
end generate;


end a1;